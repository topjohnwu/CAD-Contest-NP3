//
// Conformal-LEC Version 15.20-d250 ( 18-Apr-2016) ( 64 bit executable)
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n12345 , n12346 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 ;
output n12345 , n12346 ;

wire n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , 
     n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , 
     n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , 
     n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , 
     n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , 
     n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , 
     n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , 
     n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , 
     n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , 
     n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , 
     n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , 
     n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , 
     n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , 
     n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , 
     n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , 
     n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , 
     n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , 
     n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , 
     n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , 
     n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , 
     n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , 
     n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , 
     n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , 
     n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , 
     n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , 
     n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , 
     n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , 
     n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , 
     n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , 
     n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , 
     n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , 
     n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , 
     n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , 
     n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , 
     n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , 
     n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , 
     n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , 
     n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , 
     n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , 
     n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , 
     n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , 
     n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , 
     n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , 
     n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , 
     n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , 
     n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , 
     n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , 
     n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , 
     n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , 
     n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , 
     n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , 
     n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , 
     n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , 
     n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , 
     n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , 
     n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , 
     n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , 
     n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , 
     n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , 
     n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , 
     n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , 
     n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , 
     n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , 
     n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , 
     n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , 
     n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , 
     n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , 
     n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , 
     n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , 
     n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , 
     n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , 
     n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , 
     n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , 
     n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , 
     n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , 
     n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , 
     n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , 
     n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , 
     n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , 
     n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , 
     n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , 
     n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , 
     n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , 
     n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , 
     n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , 
     n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , 
     n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , 
     n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , 
     n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , 
     n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , 
     n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , 
     n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , 
     n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , 
     n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , 
     n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , 
     n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , 
     n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , 
     n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , 
     n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , 
     n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , 
     n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , 
     n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , 
     n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , 
     n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , 
     n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , 
     n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , 
     n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , 
     n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , 
     n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , 
     n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , 
     n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , 
     n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , 
     n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , 
     n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , 
     n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , 
     n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , 
     n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , 
     n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , 
     n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , 
     n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , 
     n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , 
     n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , 
     n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , 
     n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , 
     n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , 
     n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , 
     n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , 
     n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , 
     n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , 
     n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , 
     n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , 
     n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , 
     n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , 
     n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , 
     n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , 
     n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , 
     n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , 
     n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , 
     n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , 
     n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , 
     n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , 
     n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , 
     n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , 
     n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , 
     n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , 
     n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , 
     n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , 
     n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , 
     n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , 
     n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , 
     n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , 
     n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , 
     n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , 
     n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , 
     n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , 
     n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , 
     n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , 
     n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , 
     n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , 
     n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , 
     n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , 
     n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , 
     n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , 
     n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , 
     n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , 
     n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , 
     n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , 
     n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , 
     n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , 
     n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , 
     n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , 
     n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , 
     n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , 
     n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , 
     n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , 
     n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , 
     n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , 
     n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , 
     n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , 
     n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , 
     n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , 
     n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , 
     n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , 
     n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , 
     n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , 
     n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , 
     n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , 
     n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , 
     n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , 
     n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , 
     n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , 
     n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , 
     n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , 
     n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , 
     n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , 
     n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , 
     n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , 
     n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , 
     n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , 
     n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , 
     n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , 
     n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , 
     n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , 
     n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , 
     n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , 
     n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , 
     n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , 
     n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , 
     n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , 
     n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , 
     n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , 
     n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , 
     n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , 
     n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , 
     n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , 
     n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , 
     n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , 
     n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , 
     n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , 
     n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , 
     n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , 
     n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , 
     n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , 
     n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , 
     n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , 
     n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , 
     n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , 
     n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , 
     n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , 
     n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , 
     n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , 
     n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , 
     n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , 
     n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , 
     n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , 
     n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , 
     n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , 
     n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , 
     n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , 
     n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , 
     n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , 
     n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , 
     n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , 
     n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , 
     n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , 
     n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , 
     n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , 
     n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , 
     n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , 
     n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , 
     n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , 
     n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , 
     n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , 
     n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , 
     n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , 
     n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , 
     n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , 
     n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , 
     n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , 
     n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , 
     n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , 
     n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , 
     n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , 
     n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , 
     n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , 
     n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , 
     n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , 
     n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , 
     n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , 
     n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , 
     n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , 
     n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , 
     n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , 
     n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , 
     n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , 
     n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , 
     n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , 
     n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , 
     n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , 
     n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , 
     n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , 
     n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , 
     n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , 
     n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , 
     n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , 
     n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , 
     n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , 
     n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , 
     n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , 
     n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , 
     n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , 
     n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , 
     n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , 
     n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , 
     n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , 
     n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , 
     n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , 
     n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , 
     n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , 
     n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , 
     n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , 
     n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , 
     n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , 
     n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , 
     n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , 
     n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , 
     n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , 
     n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , 
     n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , 
     n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , 
     n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , 
     n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , 
     n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , 
     n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , 
     n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , 
     n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , 
     n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , 
     n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , 
     n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , 
     n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , 
     n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , 
     n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , 
     n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , 
     n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , 
     n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , 
     n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , 
     n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , 
     n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , 
     n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , 
     n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , 
     n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , 
     n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , 
     n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , 
     n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , 
     n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , 
     n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , 
     n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , 
     n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , 
     n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , 
     n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , 
     n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , 
     n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , 
     n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , 
     n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , 
     n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , 
     n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , 
     n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , 
     n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , 
     n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , 
     n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , 
     n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , 
     n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , 
     n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , 
     n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , 
     n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , 
     n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , 
     n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , 
     n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , 
     n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , 
     n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , 
     n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , 
     n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , 
     n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , 
     n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , 
     n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , 
     n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , 
     n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , 
     n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , 
     n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , 
     n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , 
     n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , 
     n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , 
     n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , 
     n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , 
     n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , 
     n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , 
     n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , 
     n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , 
     n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , 
     n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , 
     n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , 
     n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , 
     n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , 
     n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , 
     n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , 
     n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , 
     n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , 
     n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , 
     n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , 
     n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , 
     n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , 
     n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , 
     n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , 
     n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , 
     n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , 
     n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , 
     n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , 
     n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , 
     n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , 
     n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , 
     n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , 
     n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , 
     n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , 
     n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , 
     n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , 
     n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , 
     n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , 
     n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , 
     n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , 
     n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , 
     n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , 
     n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , 
     n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , 
     n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , 
     n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , 
     n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , 
     n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , 
     n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , 
     n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , 
     n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , 
     n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , 
     n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , 
     n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , 
     n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , 
     n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , 
     n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , 
     n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , 
     n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , 
     n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , 
     n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , 
     n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , 
     n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , 
     n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , 
     n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , 
     n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , 
     n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , 
     n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , 
     n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , 
     n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , 
     n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , 
     n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , 
     n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , 
     n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , 
     n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , 
     n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , 
     n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , 
     n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , 
     n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , 
     n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , 
     n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , 
     n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , 
     n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , 
     n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , 
     n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , 
     n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , 
     n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , 
     n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , 
     n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , 
     n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , 
     n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , 
     n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , 
     n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , 
     n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , 
     n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , 
     n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , 
     n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , 
     n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , 
     n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , 
     n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , 
     n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , 
     n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , 
     n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , 
     n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , 
     n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , 
     n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , 
     n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , 
     n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , 
     n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , 
     n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , 
     n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , 
     n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , 
     n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , 
     n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , 
     n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , 
     n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , 
     n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , 
     n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , 
     n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , 
     n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , 
     n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , 
     n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , 
     n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , 
     n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , 
     n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , 
     n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , 
     n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , 
     n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , 
     n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , 
     n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , 
     n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , 
     n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , 
     n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , 
     n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , 
     n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , 
     n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , 
     n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , 
     n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , 
     n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , 
     n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , 
     n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , 
     n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , 
     n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , 
     n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , 
     n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , 
     n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , 
     n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , 
     n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , 
     n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , 
     n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , 
     n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , 
     n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , 
     n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , 
     n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , 
     n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , 
     n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , 
     n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , 
     n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , 
     n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , 
     n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , 
     n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , 
     n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , 
     n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , 
     n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , 
     n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , 
     n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , 
     n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , 
     n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , 
     n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , 
     n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , 
     n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , 
     n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , 
     n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , 
     n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , 
     n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , 
     n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , 
     n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , 
     n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , 
     n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , 
     n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , 
     n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , 
     n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , 
     n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , 
     n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , 
     n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , 
     n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , 
     n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , 
     n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , 
     n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , 
     n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , 
     n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , 
     n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , 
     n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , 
     n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , 
     n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , 
     n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , 
     n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , 
     n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , 
     n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , 
     n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , 
     n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , 
     n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , 
     n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , 
     n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , 
     n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , 
     n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , 
     n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , 
     n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , 
     n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , 
     n6803 , n6804 , n6805 ;
buf ( n12346 , n3996 );
buf ( n12345 , n6805 );
buf ( n1026 , n172 );
buf ( n1027 , n295 );
buf ( n1028 , n114 );
buf ( n1029 , n4 );
buf ( n1030 , n13 );
buf ( n1031 , n477 );
buf ( n1032 , n151 );
buf ( n1033 , n18 );
buf ( n1034 , n364 );
buf ( n1035 , n408 );
buf ( n1036 , n160 );
buf ( n1037 , n190 );
buf ( n1038 , n339 );
buf ( n1039 , n174 );
buf ( n1040 , n181 );
buf ( n1041 , n204 );
buf ( n1042 , n302 );
buf ( n1043 , n478 );
buf ( n1044 , n435 );
buf ( n1045 , n328 );
buf ( n1046 , n39 );
buf ( n1047 , n182 );
buf ( n1048 , n327 );
buf ( n1049 , n372 );
buf ( n1050 , n467 );
buf ( n1051 , n307 );
buf ( n1052 , n154 );
buf ( n1053 , n145 );
buf ( n1054 , n127 );
buf ( n1055 , n410 );
buf ( n1056 , n143 );
buf ( n1057 , n169 );
buf ( n1058 , n432 );
buf ( n1059 , n280 );
buf ( n1060 , n142 );
buf ( n1061 , n324 );
buf ( n1062 , n36 );
buf ( n1063 , n237 );
buf ( n1064 , n359 );
buf ( n1065 , n87 );
buf ( n1066 , n215 );
buf ( n1067 , n454 );
buf ( n1068 , n336 );
buf ( n1069 , n32 );
buf ( n1070 , n136 );
buf ( n1071 , n281 );
buf ( n1072 , n325 );
buf ( n1073 , n199 );
buf ( n1074 , n140 );
buf ( n1075 , n135 );
buf ( n1076 , n148 );
buf ( n1077 , n138 );
buf ( n1078 , n49 );
buf ( n1079 , n445 );
buf ( n1080 , n278 );
buf ( n1081 , n206 );
buf ( n1082 , n17 );
buf ( n1083 , n299 );
buf ( n1084 , n398 );
buf ( n1085 , n90 );
buf ( n1086 , n92 );
buf ( n1087 , n357 );
buf ( n1088 , n149 );
buf ( n1089 , n387 );
buf ( n1090 , n420 );
buf ( n1091 , n499 );
buf ( n1092 , n98 );
buf ( n1093 , n335 );
buf ( n1094 , n439 );
buf ( n1095 , n475 );
buf ( n1096 , n482 );
buf ( n1097 , n144 );
buf ( n1098 , n202 );
buf ( n1099 , n179 );
buf ( n1100 , n100 );
buf ( n1101 , n453 );
buf ( n1102 , n103 );
buf ( n1103 , n373 );
buf ( n1104 , n483 );
buf ( n1105 , n238 );
buf ( n1106 , n342 );
buf ( n1107 , n470 );
buf ( n1108 , n77 );
buf ( n1109 , n63 );
buf ( n1110 , n170 );
buf ( n1111 , n405 );
buf ( n1112 , n10 );
buf ( n1113 , n7 );
buf ( n1114 , n27 );
buf ( n1115 , n244 );
buf ( n1116 , n388 );
buf ( n1117 , n165 );
buf ( n1118 , n166 );
buf ( n1119 , n493 );
buf ( n1120 , n55 );
buf ( n1121 , n495 );
buf ( n1122 , n487 );
buf ( n1123 , n500 );
buf ( n1124 , n81 );
buf ( n1125 , n257 );
buf ( n1126 , n448 );
buf ( n1127 , n59 );
buf ( n1128 , n226 );
buf ( n1129 , n191 );
buf ( n1130 , n137 );
buf ( n1131 , n129 );
buf ( n1132 , n194 );
buf ( n1133 , n407 );
buf ( n1134 , n109 );
buf ( n1135 , n221 );
buf ( n1136 , n68 );
buf ( n1137 , n218 );
buf ( n1138 , n437 );
buf ( n1139 , n447 );
buf ( n1140 , n455 );
buf ( n1141 , n371 );
buf ( n1142 , n390 );
buf ( n1143 , n65 );
buf ( n1144 , n292 );
buf ( n1145 , n163 );
buf ( n1146 , n61 );
buf ( n1147 , n44 );
buf ( n1148 , n6 );
buf ( n1149 , n217 );
buf ( n1150 , n314 );
buf ( n1151 , n461 );
buf ( n1152 , n250 );
buf ( n1153 , n121 );
buf ( n1154 , n64 );
buf ( n1155 , n449 );
buf ( n1156 , n310 );
buf ( n1157 , n112 );
buf ( n1158 , n26 );
buf ( n1159 , n51 );
buf ( n1160 , n348 );
buf ( n1161 , n392 );
buf ( n1162 , n249 );
buf ( n1163 , n424 );
buf ( n1164 , n115 );
buf ( n1165 , n201 );
buf ( n1166 , n396 );
buf ( n1167 , n85 );
buf ( n1168 , n219 );
buf ( n1169 , n24 );
buf ( n1170 , n356 );
buf ( n1171 , n230 );
buf ( n1172 , n20 );
buf ( n1173 , n394 );
buf ( n1174 , n93 );
buf ( n1175 , n451 );
buf ( n1176 , n267 );
buf ( n1177 , n304 );
buf ( n1178 , n76 );
buf ( n1179 , n171 );
buf ( n1180 , n241 );
buf ( n1181 , n349 );
buf ( n1182 , n350 );
buf ( n1183 , n380 );
buf ( n1184 , n3 );
buf ( n1185 , n258 );
buf ( n1186 , n25 );
buf ( n1187 , n214 );
buf ( n1188 , n481 );
buf ( n1189 , n161 );
buf ( n1190 , n429 );
buf ( n1191 , n271 );
buf ( n1192 , n353 );
buf ( n1193 , n469 );
buf ( n1194 , n38 );
buf ( n1195 , n232 );
buf ( n1196 , n188 );
buf ( n1197 , n293 );
buf ( n1198 , n246 );
buf ( n1199 , n119 );
buf ( n1200 , n463 );
buf ( n1201 , n395 );
buf ( n1202 , n494 );
buf ( n1203 , n247 );
buf ( n1204 , n303 );
buf ( n1205 , n337 );
buf ( n1206 , n287 );
buf ( n1207 , n0 );
buf ( n1208 , n133 );
buf ( n1209 , n321 );
buf ( n1210 , n414 );
buf ( n1211 , n502 );
buf ( n1212 , n284 );
buf ( n1213 , n367 );
buf ( n1214 , n34 );
buf ( n1215 , n9 );
buf ( n1216 , n362 );
buf ( n1217 , n15 );
buf ( n1218 , n393 );
buf ( n1219 , n168 );
buf ( n1220 , n436 );
buf ( n1221 , n122 );
buf ( n1222 , n426 );
buf ( n1223 , n29 );
buf ( n1224 , n110 );
buf ( n1225 , n511 );
buf ( n1226 , n162 );
buf ( n1227 , n460 );
buf ( n1228 , n476 );
buf ( n1229 , n312 );
buf ( n1230 , n320 );
buf ( n1231 , n316 );
buf ( n1232 , n153 );
buf ( n1233 , n260 );
buf ( n1234 , n427 );
buf ( n1235 , n464 );
buf ( n1236 , n415 );
buf ( n1237 , n263 );
buf ( n1238 , n377 );
buf ( n1239 , n366 );
buf ( n1240 , n57 );
buf ( n1241 , n262 );
buf ( n1242 , n497 );
buf ( n1243 , n54 );
buf ( n1244 , n401 );
buf ( n1245 , n50 );
buf ( n1246 , n400 );
buf ( n1247 , n62 );
buf ( n1248 , n265 );
buf ( n1249 , n183 );
buf ( n1250 , n459 );
buf ( n1251 , n78 );
buf ( n1252 , n173 );
buf ( n1253 , n220 );
buf ( n1254 , n277 );
buf ( n1255 , n228 );
buf ( n1256 , n14 );
buf ( n1257 , n466 );
buf ( n1258 , n235 );
buf ( n1259 , n42 );
buf ( n1260 , n37 );
buf ( n1261 , n52 );
buf ( n1262 , n31 );
buf ( n1263 , n99 );
buf ( n1264 , n355 );
buf ( n1265 , n431 );
buf ( n1266 , n286 );
buf ( n1267 , n30 );
buf ( n1268 , n229 );
buf ( n1269 , n126 );
buf ( n1270 , n306 );
buf ( n1271 , n309 );
buf ( n1272 , n2 );
buf ( n1273 , n91 );
buf ( n1274 , n243 );
buf ( n1275 , n167 );
buf ( n1276 , n223 );
buf ( n1277 , n253 );
buf ( n1278 , n368 );
buf ( n1279 , n33 );
buf ( n1280 , n313 );
buf ( n1281 , n86 );
buf ( n1282 , n180 );
buf ( n1283 , n276 );
buf ( n1284 , n240 );
buf ( n1285 , n196 );
buf ( n1286 , n340 );
buf ( n1287 , n403 );
buf ( n1288 , n70 );
buf ( n1289 , n472 );
buf ( n1290 , n130 );
buf ( n1291 , n384 );
buf ( n1292 , n402 );
buf ( n1293 , n16 );
buf ( n1294 , n224 );
buf ( n1295 , n434 );
buf ( n1296 , n389 );
buf ( n1297 , n264 );
buf ( n1298 , n326 );
buf ( n1299 , n421 );
buf ( n1300 , n411 );
buf ( n1301 , n473 );
buf ( n1302 , n334 );
buf ( n1303 , n501 );
buf ( n1304 , n212 );
buf ( n1305 , n40 );
buf ( n1306 , n118 );
buf ( n1307 , n291 );
buf ( n1308 , n471 );
buf ( n1309 , n8 );
buf ( n1310 , n124 );
buf ( n1311 , n123 );
buf ( n1312 , n239 );
buf ( n1313 , n298 );
buf ( n1314 , n382 );
buf ( n1315 , n21 );
buf ( n1316 , n457 );
buf ( n1317 , n146 );
buf ( n1318 , n106 );
buf ( n1319 , n416 );
buf ( n1320 , n120 );
buf ( n1321 , n369 );
buf ( n1322 , n474 );
buf ( n1323 , n72 );
buf ( n1324 , n269 );
buf ( n1325 , n203 );
buf ( n1326 , n490 );
buf ( n1327 , n422 );
buf ( n1328 , n233 );
buf ( n1329 , n177 );
buf ( n1330 , n94 );
buf ( n1331 , n485 );
buf ( n1332 , n294 );
buf ( n1333 , n132 );
buf ( n1334 , n419 );
buf ( n1335 , n74 );
buf ( n1336 , n60 );
buf ( n1337 , n430 );
buf ( n1338 , n150 );
buf ( n1339 , n197 );
buf ( n1340 , n283 );
buf ( n1341 , n254 );
buf ( n1342 , n375 );
buf ( n1343 , n505 );
buf ( n1344 , n443 );
buf ( n1345 , n290 );
buf ( n1346 , n365 );
buf ( n1347 , n139 );
buf ( n1348 , n256 );
buf ( n1349 , n19 );
buf ( n1350 , n53 );
buf ( n1351 , n452 );
buf ( n1352 , n479 );
buf ( n1353 , n381 );
buf ( n1354 , n346 );
buf ( n1355 , n178 );
buf ( n1356 , n272 );
buf ( n1357 , n234 );
buf ( n1358 , n12 );
buf ( n1359 , n67 );
buf ( n1360 , n386 );
buf ( n1361 , n282 );
buf ( n1362 , n509 );
buf ( n1363 , n164 );
buf ( n1364 , n297 );
buf ( n1365 , n211 );
buf ( n1366 , n274 );
buf ( n1367 , n425 );
buf ( n1368 , n113 );
buf ( n1369 , n345 );
buf ( n1370 , n66 );
buf ( n1371 , n317 );
buf ( n1372 , n341 );
buf ( n1373 , n496 );
buf ( n1374 , n358 );
buf ( n1375 , n80 );
buf ( n1376 , n268 );
buf ( n1377 , n108 );
buf ( n1378 , n22 );
buf ( n1379 , n96 );
buf ( n1380 , n159 );
buf ( n1381 , n189 );
buf ( n1382 , n361 );
buf ( n1383 , n107 );
buf ( n1384 , n370 );
buf ( n1385 , n315 );
buf ( n1386 , n409 );
buf ( n1387 , n35 );
buf ( n1388 , n305 );
buf ( n1389 , n175 );
buf ( n1390 , n423 );
buf ( n1391 , n155 );
buf ( n1392 , n200 );
buf ( n1393 , n385 );
buf ( n1394 , n344 );
buf ( n1395 , n208 );
buf ( n1396 , n227 );
buf ( n1397 , n441 );
buf ( n1398 , n69 );
buf ( n1399 , n95 );
buf ( n1400 , n251 );
buf ( n1401 , n506 );
buf ( n1402 , n503 );
buf ( n1403 , n508 );
buf ( n1404 , n156 );
buf ( n1405 , n418 );
buf ( n1406 , n510 );
buf ( n1407 , n275 );
buf ( n1408 , n97 );
buf ( n1409 , n289 );
buf ( n1410 , n184 );
buf ( n1411 , n308 );
buf ( n1412 , n259 );
buf ( n1413 , n210 );
buf ( n1414 , n507 );
buf ( n1415 , n41 );
buf ( n1416 , n323 );
buf ( n1417 , n488 );
buf ( n1418 , n128 );
buf ( n1419 , n504 );
buf ( n1420 , n333 );
buf ( n1421 , n347 );
buf ( n1422 , n406 );
buf ( n1423 , n245 );
buf ( n1424 , n213 );
buf ( n1425 , n141 );
buf ( n1426 , n270 );
buf ( n1427 , n363 );
buf ( n1428 , n236 );
buf ( n1429 , n444 );
buf ( n1430 , n28 );
buf ( n1431 , n300 );
buf ( n1432 , n288 );
buf ( n1433 , n102 );
buf ( n1434 , n329 );
buf ( n1435 , n207 );
buf ( n1436 , n176 );
buf ( n1437 , n442 );
buf ( n1438 , n43 );
buf ( n1439 , n83 );
buf ( n1440 , n417 );
buf ( n1441 , n376 );
buf ( n1442 , n456 );
buf ( n1443 , n58 );
buf ( n1444 , n480 );
buf ( n1445 , n46 );
buf ( n1446 , n492 );
buf ( n1447 , n125 );
buf ( n1448 , n413 );
buf ( n1449 , n433 );
buf ( n1450 , n318 );
buf ( n1451 , n412 );
buf ( n1452 , n484 );
buf ( n1453 , n397 );
buf ( n1454 , n158 );
buf ( n1455 , n343 );
buf ( n1456 , n242 );
buf ( n1457 , n330 );
buf ( n1458 , n198 );
buf ( n1459 , n195 );
buf ( n1460 , n187 );
buf ( n1461 , n352 );
buf ( n1462 , n101 );
buf ( n1463 , n354 );
buf ( n1464 , n379 );
buf ( n1465 , n88 );
buf ( n1466 , n332 );
buf ( n1467 , n331 );
buf ( n1468 , n491 );
buf ( n1469 , n378 );
buf ( n1470 , n489 );
buf ( n1471 , n360 );
buf ( n1472 , n147 );
buf ( n1473 , n104 );
buf ( n1474 , n89 );
buf ( n1475 , n82 );
buf ( n1476 , n446 );
buf ( n1477 , n205 );
buf ( n1478 , n216 );
buf ( n1479 , n296 );
buf ( n1480 , n84 );
buf ( n1481 , n75 );
buf ( n1482 , n5 );
buf ( n1483 , n1 );
buf ( n1484 , n192 );
buf ( n1485 , n383 );
buf ( n1486 , n117 );
buf ( n1487 , n450 );
buf ( n1488 , n45 );
buf ( n1489 , n71 );
buf ( n1490 , n498 );
buf ( n1491 , n48 );
buf ( n1492 , n301 );
buf ( n1493 , n440 );
buf ( n1494 , n111 );
buf ( n1495 , n152 );
buf ( n1496 , n428 );
buf ( n1497 , n47 );
buf ( n1498 , n193 );
buf ( n1499 , n351 );
buf ( n1500 , n131 );
buf ( n1501 , n404 );
buf ( n1502 , n399 );
buf ( n1503 , n252 );
buf ( n1504 , n458 );
buf ( n1505 , n105 );
buf ( n1506 , n231 );
buf ( n1507 , n273 );
buf ( n1508 , n266 );
buf ( n1509 , n255 );
buf ( n1510 , n185 );
buf ( n1511 , n56 );
buf ( n1512 , n248 );
buf ( n1513 , n438 );
buf ( n1514 , n261 );
buf ( n1515 , n468 );
buf ( n1516 , n23 );
buf ( n1517 , n311 );
buf ( n1518 , n279 );
buf ( n1519 , n338 );
buf ( n1520 , n79 );
buf ( n1521 , n285 );
buf ( n1522 , n222 );
buf ( n1523 , n73 );
buf ( n1524 , n116 );
buf ( n1525 , n225 );
buf ( n1526 , n209 );
buf ( n1527 , n157 );
buf ( n1528 , n319 );
buf ( n1529 , n391 );
buf ( n1530 , n134 );
buf ( n1531 , n462 );
buf ( n1532 , n374 );
buf ( n1533 , n322 );
buf ( n1534 , n186 );
buf ( n1535 , n486 );
buf ( n1536 , n465 );
buf ( n1537 , n11 );
buf ( n1538 , n1026 );
buf ( n1539 , n1282 );
xor ( n1540 , n1538 , n1539 );
buf ( n1541 , n1027 );
buf ( n1542 , n1283 );
and ( n1543 , n1541 , n1542 );
buf ( n1544 , n1028 );
buf ( n1545 , n1284 );
and ( n1546 , n1544 , n1545 );
buf ( n1547 , n1029 );
buf ( n1548 , n1285 );
and ( n1549 , n1547 , n1548 );
buf ( n1550 , n1030 );
buf ( n1551 , n1286 );
and ( n1552 , n1550 , n1551 );
buf ( n1553 , n1031 );
buf ( n1554 , n1287 );
and ( n1555 , n1553 , n1554 );
buf ( n1556 , n1032 );
buf ( n1557 , n1288 );
and ( n1558 , n1556 , n1557 );
buf ( n1559 , n1033 );
buf ( n1560 , n1289 );
and ( n1561 , n1559 , n1560 );
buf ( n1562 , n1034 );
buf ( n1563 , n1290 );
and ( n1564 , n1562 , n1563 );
buf ( n1565 , n1035 );
buf ( n1566 , n1291 );
and ( n1567 , n1565 , n1566 );
buf ( n1568 , n1036 );
buf ( n1569 , n1292 );
and ( n1570 , n1568 , n1569 );
buf ( n1571 , n1037 );
buf ( n1572 , n1293 );
and ( n1573 , n1571 , n1572 );
buf ( n1574 , n1038 );
buf ( n1575 , n1294 );
and ( n1576 , n1574 , n1575 );
buf ( n1577 , n1039 );
buf ( n1578 , n1295 );
and ( n1579 , n1577 , n1578 );
buf ( n1580 , n1040 );
buf ( n1581 , n1296 );
and ( n1582 , n1580 , n1581 );
buf ( n1583 , n1041 );
buf ( n1584 , n1297 );
and ( n1585 , n1583 , n1584 );
buf ( n1586 , n1042 );
buf ( n1587 , n1298 );
and ( n1588 , n1586 , n1587 );
buf ( n1589 , n1043 );
buf ( n1590 , n1299 );
and ( n1591 , n1589 , n1590 );
buf ( n1592 , n1044 );
buf ( n1593 , n1300 );
and ( n1594 , n1592 , n1593 );
buf ( n1595 , n1045 );
buf ( n1596 , n1301 );
and ( n1597 , n1595 , n1596 );
buf ( n1598 , n1046 );
buf ( n1599 , n1302 );
and ( n1600 , n1598 , n1599 );
buf ( n1601 , n1047 );
buf ( n1602 , n1303 );
and ( n1603 , n1601 , n1602 );
buf ( n1604 , n1048 );
buf ( n1605 , n1304 );
and ( n1606 , n1604 , n1605 );
buf ( n1607 , n1049 );
buf ( n1608 , n1305 );
and ( n1609 , n1607 , n1608 );
buf ( n1610 , n1050 );
buf ( n1611 , n1306 );
and ( n1612 , n1610 , n1611 );
buf ( n1613 , n1051 );
buf ( n1614 , n1307 );
and ( n1615 , n1613 , n1614 );
buf ( n1616 , n1052 );
buf ( n1617 , n1308 );
and ( n1618 , n1616 , n1617 );
buf ( n1619 , n1053 );
buf ( n1620 , n1309 );
and ( n1621 , n1619 , n1620 );
buf ( n1622 , n1054 );
buf ( n1623 , n1310 );
and ( n1624 , n1622 , n1623 );
buf ( n1625 , n1055 );
buf ( n1626 , n1311 );
and ( n1627 , n1625 , n1626 );
buf ( n1628 , n1056 );
buf ( n1629 , n1312 );
and ( n1630 , n1628 , n1629 );
buf ( n1631 , n1057 );
buf ( n1632 , n1313 );
and ( n1633 , n1631 , n1632 );
buf ( n1634 , n1058 );
buf ( n1635 , n1314 );
and ( n1636 , n1634 , n1635 );
buf ( n1637 , n1059 );
buf ( n1638 , n1315 );
and ( n1639 , n1637 , n1638 );
buf ( n1640 , n1060 );
buf ( n1641 , n1316 );
and ( n1642 , n1640 , n1641 );
buf ( n1643 , n1061 );
buf ( n1644 , n1317 );
and ( n1645 , n1643 , n1644 );
buf ( n1646 , n1062 );
buf ( n1647 , n1318 );
and ( n1648 , n1646 , n1647 );
buf ( n1649 , n1063 );
buf ( n1650 , n1319 );
and ( n1651 , n1649 , n1650 );
buf ( n1652 , n1064 );
buf ( n1653 , n1320 );
and ( n1654 , n1652 , n1653 );
buf ( n1655 , n1065 );
buf ( n1656 , n1321 );
and ( n1657 , n1655 , n1656 );
buf ( n1658 , n1066 );
buf ( n1659 , n1322 );
and ( n1660 , n1658 , n1659 );
buf ( n1661 , n1067 );
buf ( n1662 , n1323 );
and ( n1663 , n1661 , n1662 );
buf ( n1664 , n1068 );
buf ( n1665 , n1324 );
and ( n1666 , n1664 , n1665 );
buf ( n1667 , n1069 );
buf ( n1668 , n1325 );
and ( n1669 , n1667 , n1668 );
buf ( n1670 , n1070 );
buf ( n1671 , n1326 );
and ( n1672 , n1670 , n1671 );
buf ( n1673 , n1071 );
buf ( n1674 , n1327 );
and ( n1675 , n1673 , n1674 );
buf ( n1676 , n1072 );
buf ( n1677 , n1328 );
and ( n1678 , n1676 , n1677 );
buf ( n1679 , n1073 );
buf ( n1680 , n1329 );
and ( n1681 , n1679 , n1680 );
buf ( n1682 , n1074 );
buf ( n1683 , n1330 );
and ( n1684 , n1682 , n1683 );
buf ( n1685 , n1075 );
buf ( n1686 , n1331 );
and ( n1687 , n1685 , n1686 );
buf ( n1688 , n1076 );
buf ( n1689 , n1332 );
and ( n1690 , n1688 , n1689 );
buf ( n1691 , n1077 );
buf ( n1692 , n1333 );
and ( n1693 , n1691 , n1692 );
buf ( n1694 , n1078 );
buf ( n1695 , n1334 );
and ( n1696 , n1694 , n1695 );
buf ( n1697 , n1079 );
buf ( n1698 , n1335 );
and ( n1699 , n1697 , n1698 );
buf ( n1700 , n1080 );
buf ( n1701 , n1336 );
and ( n1702 , n1700 , n1701 );
buf ( n1703 , n1081 );
buf ( n1704 , n1337 );
and ( n1705 , n1703 , n1704 );
buf ( n1706 , n1082 );
buf ( n1707 , n1338 );
and ( n1708 , n1706 , n1707 );
buf ( n1709 , n1083 );
buf ( n1710 , n1339 );
and ( n1711 , n1709 , n1710 );
buf ( n1712 , n1084 );
buf ( n1713 , n1340 );
and ( n1714 , n1712 , n1713 );
buf ( n1715 , n1085 );
buf ( n1716 , n1341 );
and ( n1717 , n1715 , n1716 );
buf ( n1718 , n1086 );
buf ( n1719 , n1342 );
and ( n1720 , n1718 , n1719 );
buf ( n1721 , n1087 );
buf ( n1722 , n1343 );
and ( n1723 , n1721 , n1722 );
buf ( n1724 , n1088 );
buf ( n1725 , n1344 );
and ( n1726 , n1724 , n1725 );
buf ( n1727 , n1089 );
buf ( n1728 , n1345 );
and ( n1729 , n1727 , n1728 );
buf ( n1730 , n1090 );
buf ( n1731 , n1346 );
and ( n1732 , n1730 , n1731 );
buf ( n1733 , n1091 );
buf ( n1734 , n1347 );
and ( n1735 , n1733 , n1734 );
buf ( n1736 , n1092 );
buf ( n1737 , n1348 );
and ( n1738 , n1736 , n1737 );
buf ( n1739 , n1093 );
buf ( n1740 , n1349 );
and ( n1741 , n1739 , n1740 );
buf ( n1742 , n1094 );
buf ( n1743 , n1350 );
and ( n1744 , n1742 , n1743 );
buf ( n1745 , n1095 );
buf ( n1746 , n1351 );
and ( n1747 , n1745 , n1746 );
buf ( n1748 , n1096 );
buf ( n1749 , n1352 );
and ( n1750 , n1748 , n1749 );
buf ( n1751 , n1097 );
buf ( n1752 , n1353 );
and ( n1753 , n1751 , n1752 );
buf ( n1754 , n1098 );
buf ( n1755 , n1354 );
and ( n1756 , n1754 , n1755 );
buf ( n1757 , n1099 );
buf ( n1758 , n1355 );
and ( n1759 , n1757 , n1758 );
buf ( n1760 , n1100 );
buf ( n1761 , n1356 );
and ( n1762 , n1760 , n1761 );
buf ( n1763 , n1101 );
buf ( n1764 , n1357 );
and ( n1765 , n1763 , n1764 );
buf ( n1766 , n1102 );
buf ( n1767 , n1358 );
and ( n1768 , n1766 , n1767 );
buf ( n1769 , n1103 );
buf ( n1770 , n1359 );
and ( n1771 , n1769 , n1770 );
buf ( n1772 , n1104 );
buf ( n1773 , n1360 );
and ( n1774 , n1772 , n1773 );
buf ( n1775 , n1105 );
buf ( n1776 , n1361 );
and ( n1777 , n1775 , n1776 );
buf ( n1778 , n1106 );
buf ( n1779 , n1362 );
and ( n1780 , n1778 , n1779 );
buf ( n1781 , n1107 );
buf ( n1782 , n1363 );
and ( n1783 , n1781 , n1782 );
buf ( n1784 , n1108 );
buf ( n1785 , n1364 );
and ( n1786 , n1784 , n1785 );
buf ( n1787 , n1109 );
buf ( n1788 , n1365 );
and ( n1789 , n1787 , n1788 );
buf ( n1790 , n1110 );
buf ( n1791 , n1366 );
and ( n1792 , n1790 , n1791 );
buf ( n1793 , n1111 );
buf ( n1794 , n1367 );
and ( n1795 , n1793 , n1794 );
buf ( n1796 , n1112 );
buf ( n1797 , n1368 );
and ( n1798 , n1796 , n1797 );
buf ( n1799 , n1113 );
buf ( n1800 , n1369 );
and ( n1801 , n1799 , n1800 );
buf ( n1802 , n1114 );
buf ( n1803 , n1370 );
and ( n1804 , n1802 , n1803 );
buf ( n1805 , n1115 );
buf ( n1806 , n1371 );
and ( n1807 , n1805 , n1806 );
buf ( n1808 , n1116 );
buf ( n1809 , n1372 );
and ( n1810 , n1808 , n1809 );
buf ( n1811 , n1117 );
buf ( n1812 , n1373 );
and ( n1813 , n1811 , n1812 );
buf ( n1814 , n1118 );
buf ( n1815 , n1374 );
and ( n1816 , n1814 , n1815 );
buf ( n1817 , n1119 );
buf ( n1818 , n1375 );
and ( n1819 , n1817 , n1818 );
buf ( n1820 , n1120 );
buf ( n1821 , n1376 );
and ( n1822 , n1820 , n1821 );
buf ( n1823 , n1121 );
buf ( n1824 , n1377 );
and ( n1825 , n1823 , n1824 );
buf ( n1826 , n1122 );
buf ( n1827 , n1378 );
and ( n1828 , n1826 , n1827 );
buf ( n1829 , n1123 );
buf ( n1830 , n1379 );
and ( n1831 , n1829 , n1830 );
buf ( n1832 , n1124 );
buf ( n1833 , n1380 );
and ( n1834 , n1832 , n1833 );
buf ( n1835 , n1125 );
buf ( n1836 , n1381 );
and ( n1837 , n1835 , n1836 );
buf ( n1838 , n1126 );
buf ( n1839 , n1382 );
and ( n1840 , n1838 , n1839 );
buf ( n1841 , n1127 );
buf ( n1842 , n1383 );
and ( n1843 , n1841 , n1842 );
buf ( n1844 , n1128 );
buf ( n1845 , n1384 );
and ( n1846 , n1844 , n1845 );
buf ( n1847 , n1129 );
buf ( n1848 , n1385 );
and ( n1849 , n1847 , n1848 );
buf ( n1850 , n1130 );
buf ( n1851 , n1386 );
and ( n1852 , n1850 , n1851 );
buf ( n1853 , n1131 );
buf ( n1854 , n1387 );
and ( n1855 , n1853 , n1854 );
buf ( n1856 , n1132 );
buf ( n1857 , n1388 );
and ( n1858 , n1856 , n1857 );
buf ( n1859 , n1133 );
buf ( n1860 , n1389 );
and ( n1861 , n1859 , n1860 );
buf ( n1862 , n1134 );
buf ( n1863 , n1390 );
and ( n1864 , n1862 , n1863 );
buf ( n1865 , n1135 );
buf ( n1866 , n1391 );
and ( n1867 , n1865 , n1866 );
buf ( n1868 , n1136 );
buf ( n1869 , n1392 );
and ( n1870 , n1868 , n1869 );
buf ( n1871 , n1137 );
buf ( n1872 , n1393 );
and ( n1873 , n1871 , n1872 );
buf ( n1874 , n1138 );
buf ( n1875 , n1394 );
and ( n1876 , n1874 , n1875 );
buf ( n1877 , n1139 );
buf ( n1878 , n1395 );
and ( n1879 , n1877 , n1878 );
buf ( n1880 , n1140 );
buf ( n1881 , n1396 );
and ( n1882 , n1880 , n1881 );
buf ( n1883 , n1141 );
buf ( n1884 , n1397 );
and ( n1885 , n1883 , n1884 );
buf ( n1886 , n1142 );
buf ( n1887 , n1398 );
and ( n1888 , n1886 , n1887 );
buf ( n1889 , n1143 );
buf ( n1890 , n1399 );
and ( n1891 , n1889 , n1890 );
buf ( n1892 , n1144 );
buf ( n1893 , n1400 );
and ( n1894 , n1892 , n1893 );
buf ( n1895 , n1145 );
buf ( n1896 , n1401 );
and ( n1897 , n1895 , n1896 );
buf ( n1898 , n1146 );
buf ( n1899 , n1402 );
and ( n1900 , n1898 , n1899 );
buf ( n1901 , n1147 );
buf ( n1902 , n1403 );
and ( n1903 , n1901 , n1902 );
buf ( n1904 , n1148 );
buf ( n1905 , n1404 );
and ( n1906 , n1904 , n1905 );
buf ( n1907 , n1149 );
buf ( n1908 , n1405 );
and ( n1909 , n1907 , n1908 );
buf ( n1910 , n1150 );
buf ( n1911 , n1406 );
and ( n1912 , n1910 , n1911 );
buf ( n1913 , n1151 );
buf ( n1914 , n1407 );
and ( n1915 , n1913 , n1914 );
buf ( n1916 , n1152 );
buf ( n1917 , n1408 );
and ( n1918 , n1916 , n1917 );
buf ( n1919 , n1153 );
buf ( n1920 , n1409 );
and ( n1921 , n1919 , n1920 );
buf ( n1922 , n1154 );
buf ( n1923 , n1410 );
and ( n1924 , n1922 , n1923 );
buf ( n1925 , n1155 );
buf ( n1926 , n1411 );
and ( n1927 , n1925 , n1926 );
buf ( n1928 , n1156 );
buf ( n1929 , n1412 );
and ( n1930 , n1928 , n1929 );
buf ( n1931 , n1157 );
buf ( n1932 , n1413 );
and ( n1933 , n1931 , n1932 );
buf ( n1934 , n1158 );
buf ( n1935 , n1414 );
and ( n1936 , n1934 , n1935 );
buf ( n1937 , n1159 );
buf ( n1938 , n1415 );
and ( n1939 , n1937 , n1938 );
buf ( n1940 , n1160 );
buf ( n1941 , n1416 );
and ( n1942 , n1940 , n1941 );
buf ( n1943 , n1161 );
buf ( n1944 , n1417 );
and ( n1945 , n1943 , n1944 );
buf ( n1946 , n1162 );
buf ( n1947 , n1418 );
and ( n1948 , n1946 , n1947 );
buf ( n1949 , n1163 );
buf ( n1950 , n1419 );
and ( n1951 , n1949 , n1950 );
buf ( n1952 , n1164 );
buf ( n1953 , n1420 );
and ( n1954 , n1952 , n1953 );
buf ( n1955 , n1165 );
buf ( n1956 , n1421 );
and ( n1957 , n1955 , n1956 );
buf ( n1958 , n1166 );
buf ( n1959 , n1422 );
and ( n1960 , n1958 , n1959 );
buf ( n1961 , n1167 );
buf ( n1962 , n1423 );
and ( n1963 , n1961 , n1962 );
buf ( n1964 , n1168 );
buf ( n1965 , n1424 );
and ( n1966 , n1964 , n1965 );
buf ( n1967 , n1169 );
buf ( n1968 , n1425 );
and ( n1969 , n1967 , n1968 );
buf ( n1970 , n1170 );
buf ( n1971 , n1426 );
and ( n1972 , n1970 , n1971 );
buf ( n1973 , n1171 );
buf ( n1974 , n1427 );
and ( n1975 , n1973 , n1974 );
buf ( n1976 , n1172 );
buf ( n1977 , n1428 );
and ( n1978 , n1976 , n1977 );
buf ( n1979 , n1173 );
buf ( n1980 , n1429 );
and ( n1981 , n1979 , n1980 );
buf ( n1982 , n1174 );
buf ( n1983 , n1430 );
and ( n1984 , n1982 , n1983 );
buf ( n1985 , n1175 );
buf ( n1986 , n1431 );
and ( n1987 , n1985 , n1986 );
buf ( n1988 , n1176 );
buf ( n1989 , n1432 );
and ( n1990 , n1988 , n1989 );
buf ( n1991 , n1177 );
buf ( n1992 , n1433 );
and ( n1993 , n1991 , n1992 );
buf ( n1994 , n1178 );
buf ( n1995 , n1434 );
and ( n1996 , n1994 , n1995 );
buf ( n1997 , n1179 );
buf ( n1998 , n1435 );
and ( n1999 , n1997 , n1998 );
buf ( n2000 , n1180 );
buf ( n2001 , n1436 );
and ( n2002 , n2000 , n2001 );
buf ( n2003 , n1181 );
buf ( n2004 , n1437 );
and ( n2005 , n2003 , n2004 );
buf ( n2006 , n1182 );
buf ( n2007 , n1438 );
and ( n2008 , n2006 , n2007 );
buf ( n2009 , n1183 );
buf ( n2010 , n1439 );
and ( n2011 , n2009 , n2010 );
buf ( n2012 , n1184 );
buf ( n2013 , n1440 );
and ( n2014 , n2012 , n2013 );
buf ( n2015 , n1185 );
buf ( n2016 , n1441 );
and ( n2017 , n2015 , n2016 );
buf ( n2018 , n1186 );
buf ( n2019 , n1442 );
and ( n2020 , n2018 , n2019 );
buf ( n2021 , n1187 );
buf ( n2022 , n1443 );
and ( n2023 , n2021 , n2022 );
buf ( n2024 , n1188 );
buf ( n2025 , n1444 );
and ( n2026 , n2024 , n2025 );
buf ( n2027 , n1189 );
buf ( n2028 , n1445 );
and ( n2029 , n2027 , n2028 );
buf ( n2030 , n1190 );
buf ( n2031 , n1446 );
and ( n2032 , n2030 , n2031 );
buf ( n2033 , n1191 );
buf ( n2034 , n1447 );
and ( n2035 , n2033 , n2034 );
buf ( n2036 , n1192 );
buf ( n2037 , n1448 );
and ( n2038 , n2036 , n2037 );
buf ( n2039 , n1193 );
buf ( n2040 , n1449 );
and ( n2041 , n2039 , n2040 );
buf ( n2042 , n1194 );
buf ( n2043 , n1450 );
and ( n2044 , n2042 , n2043 );
buf ( n2045 , n1195 );
buf ( n2046 , n1451 );
and ( n2047 , n2045 , n2046 );
buf ( n2048 , n1196 );
buf ( n2049 , n1452 );
and ( n2050 , n2048 , n2049 );
buf ( n2051 , n1197 );
buf ( n2052 , n1453 );
and ( n2053 , n2051 , n2052 );
buf ( n2054 , n1198 );
buf ( n2055 , n1454 );
and ( n2056 , n2054 , n2055 );
buf ( n2057 , n1199 );
buf ( n2058 , n1455 );
and ( n2059 , n2057 , n2058 );
buf ( n2060 , n1200 );
buf ( n2061 , n1456 );
and ( n2062 , n2060 , n2061 );
buf ( n2063 , n1201 );
buf ( n2064 , n1457 );
and ( n2065 , n2063 , n2064 );
buf ( n2066 , n1202 );
buf ( n2067 , n1458 );
and ( n2068 , n2066 , n2067 );
buf ( n2069 , n1203 );
buf ( n2070 , n1459 );
and ( n2071 , n2069 , n2070 );
buf ( n2072 , n1204 );
buf ( n2073 , n1460 );
and ( n2074 , n2072 , n2073 );
buf ( n2075 , n1205 );
buf ( n2076 , n1461 );
and ( n2077 , n2075 , n2076 );
buf ( n2078 , n1206 );
buf ( n2079 , n1462 );
and ( n2080 , n2078 , n2079 );
buf ( n2081 , n1207 );
buf ( n2082 , n1463 );
and ( n2083 , n2081 , n2082 );
buf ( n2084 , n1208 );
buf ( n2085 , n1464 );
and ( n2086 , n2084 , n2085 );
buf ( n2087 , n1209 );
buf ( n2088 , n1465 );
and ( n2089 , n2087 , n2088 );
buf ( n2090 , n1210 );
buf ( n2091 , n1466 );
and ( n2092 , n2090 , n2091 );
buf ( n2093 , n1211 );
buf ( n2094 , n1467 );
and ( n2095 , n2093 , n2094 );
buf ( n2096 , n1212 );
buf ( n2097 , n1468 );
and ( n2098 , n2096 , n2097 );
buf ( n2099 , n1213 );
buf ( n2100 , n1469 );
and ( n2101 , n2099 , n2100 );
buf ( n2102 , n1214 );
buf ( n2103 , n1470 );
and ( n2104 , n2102 , n2103 );
buf ( n2105 , n1215 );
buf ( n2106 , n1471 );
and ( n2107 , n2105 , n2106 );
buf ( n2108 , n1216 );
buf ( n2109 , n1472 );
and ( n2110 , n2108 , n2109 );
buf ( n2111 , n1217 );
buf ( n2112 , n1473 );
and ( n2113 , n2111 , n2112 );
buf ( n2114 , n1218 );
buf ( n2115 , n1474 );
and ( n2116 , n2114 , n2115 );
buf ( n2117 , n1219 );
buf ( n2118 , n1475 );
and ( n2119 , n2117 , n2118 );
buf ( n2120 , n1220 );
buf ( n2121 , n1476 );
and ( n2122 , n2120 , n2121 );
buf ( n2123 , n1221 );
buf ( n2124 , n1477 );
and ( n2125 , n2123 , n2124 );
buf ( n2126 , n1222 );
buf ( n2127 , n1478 );
and ( n2128 , n2126 , n2127 );
buf ( n2129 , n1223 );
buf ( n2130 , n1479 );
and ( n2131 , n2129 , n2130 );
buf ( n2132 , n1224 );
buf ( n2133 , n1480 );
and ( n2134 , n2132 , n2133 );
buf ( n2135 , n1225 );
buf ( n2136 , n1481 );
and ( n2137 , n2135 , n2136 );
buf ( n2138 , n1226 );
buf ( n2139 , n1482 );
and ( n2140 , n2138 , n2139 );
buf ( n2141 , n1227 );
buf ( n2142 , n1483 );
and ( n2143 , n2141 , n2142 );
buf ( n2144 , n1228 );
buf ( n2145 , n1484 );
and ( n2146 , n2144 , n2145 );
buf ( n2147 , n1229 );
buf ( n2148 , n1485 );
and ( n2149 , n2147 , n2148 );
buf ( n2150 , n1230 );
buf ( n2151 , n1486 );
and ( n2152 , n2150 , n2151 );
buf ( n2153 , n1231 );
buf ( n2154 , n1487 );
and ( n2155 , n2153 , n2154 );
buf ( n2156 , n1232 );
buf ( n2157 , n1488 );
and ( n2158 , n2156 , n2157 );
buf ( n2159 , n1233 );
buf ( n2160 , n1489 );
and ( n2161 , n2159 , n2160 );
buf ( n2162 , n1234 );
buf ( n2163 , n1490 );
and ( n2164 , n2162 , n2163 );
buf ( n2165 , n1235 );
buf ( n2166 , n1491 );
and ( n2167 , n2165 , n2166 );
buf ( n2168 , n1236 );
buf ( n2169 , n1492 );
and ( n2170 , n2168 , n2169 );
buf ( n2171 , n1237 );
buf ( n2172 , n1493 );
and ( n2173 , n2171 , n2172 );
buf ( n2174 , n1238 );
buf ( n2175 , n1494 );
and ( n2176 , n2174 , n2175 );
buf ( n2177 , n1239 );
buf ( n2178 , n1495 );
and ( n2179 , n2177 , n2178 );
buf ( n2180 , n1240 );
buf ( n2181 , n1496 );
and ( n2182 , n2180 , n2181 );
buf ( n2183 , n1241 );
buf ( n2184 , n1497 );
and ( n2185 , n2183 , n2184 );
buf ( n2186 , n1242 );
buf ( n2187 , n1498 );
and ( n2188 , n2186 , n2187 );
buf ( n2189 , n1243 );
buf ( n2190 , n1499 );
and ( n2191 , n2189 , n2190 );
buf ( n2192 , n1244 );
buf ( n2193 , n1500 );
and ( n2194 , n2192 , n2193 );
buf ( n2195 , n1245 );
buf ( n2196 , n1501 );
and ( n2197 , n2195 , n2196 );
buf ( n2198 , n1246 );
buf ( n2199 , n1502 );
and ( n2200 , n2198 , n2199 );
buf ( n2201 , n1247 );
buf ( n2202 , n1503 );
and ( n2203 , n2201 , n2202 );
buf ( n2204 , n1248 );
buf ( n2205 , n1504 );
and ( n2206 , n2204 , n2205 );
buf ( n2207 , n1249 );
buf ( n2208 , n1505 );
and ( n2209 , n2207 , n2208 );
buf ( n2210 , n1250 );
buf ( n2211 , n1506 );
and ( n2212 , n2210 , n2211 );
buf ( n2213 , n1251 );
buf ( n2214 , n1507 );
and ( n2215 , n2213 , n2214 );
buf ( n2216 , n1252 );
buf ( n2217 , n1508 );
and ( n2218 , n2216 , n2217 );
buf ( n2219 , n1253 );
buf ( n2220 , n1509 );
and ( n2221 , n2219 , n2220 );
buf ( n2222 , n1254 );
buf ( n2223 , n1510 );
and ( n2224 , n2222 , n2223 );
buf ( n2225 , n1255 );
buf ( n2226 , n1511 );
and ( n2227 , n2225 , n2226 );
buf ( n2228 , n1256 );
buf ( n2229 , n1512 );
and ( n2230 , n2228 , n2229 );
buf ( n2231 , n1257 );
buf ( n2232 , n1513 );
and ( n2233 , n2231 , n2232 );
buf ( n2234 , n1258 );
buf ( n2235 , n2234 );
buf ( n2236 , n1259 );
buf ( n2237 , n1515 );
and ( n2238 , n2236 , n2237 );
buf ( n2239 , n1260 );
buf ( n2240 , n1516 );
and ( n2241 , n2239 , n2240 );
buf ( n2242 , n2240 );
buf ( n2243 , n2239 );
or ( n2244 , n2241 , n2242 , n2243 );
and ( n2245 , n2237 , n2244 );
and ( n2246 , n2236 , n2244 );
or ( n2247 , n2238 , n2245 , n2246 );
buf ( n2248 , n2247 );
and ( n2249 , n2234 , n2247 );
or ( n2250 , n2235 , n2248 , n2249 );
and ( n2251 , n2232 , n2250 );
and ( n2252 , n2231 , n2250 );
or ( n2253 , n2233 , n2251 , n2252 );
and ( n2254 , n2229 , n2253 );
and ( n2255 , n2228 , n2253 );
or ( n2256 , n2230 , n2254 , n2255 );
and ( n2257 , n2226 , n2256 );
and ( n2258 , n2225 , n2256 );
or ( n2259 , n2227 , n2257 , n2258 );
and ( n2260 , n2223 , n2259 );
and ( n2261 , n2222 , n2259 );
or ( n2262 , n2224 , n2260 , n2261 );
and ( n2263 , n2220 , n2262 );
and ( n2264 , n2219 , n2262 );
or ( n2265 , n2221 , n2263 , n2264 );
and ( n2266 , n2217 , n2265 );
and ( n2267 , n2216 , n2265 );
or ( n2268 , n2218 , n2266 , n2267 );
and ( n2269 , n2214 , n2268 );
and ( n2270 , n2213 , n2268 );
or ( n2271 , n2215 , n2269 , n2270 );
and ( n2272 , n2211 , n2271 );
and ( n2273 , n2210 , n2271 );
or ( n2274 , n2212 , n2272 , n2273 );
and ( n2275 , n2208 , n2274 );
and ( n2276 , n2207 , n2274 );
or ( n2277 , n2209 , n2275 , n2276 );
and ( n2278 , n2205 , n2277 );
and ( n2279 , n2204 , n2277 );
or ( n2280 , n2206 , n2278 , n2279 );
and ( n2281 , n2202 , n2280 );
and ( n2282 , n2201 , n2280 );
or ( n2283 , n2203 , n2281 , n2282 );
and ( n2284 , n2199 , n2283 );
and ( n2285 , n2198 , n2283 );
or ( n2286 , n2200 , n2284 , n2285 );
and ( n2287 , n2196 , n2286 );
and ( n2288 , n2195 , n2286 );
or ( n2289 , n2197 , n2287 , n2288 );
and ( n2290 , n2193 , n2289 );
and ( n2291 , n2192 , n2289 );
or ( n2292 , n2194 , n2290 , n2291 );
and ( n2293 , n2190 , n2292 );
and ( n2294 , n2189 , n2292 );
or ( n2295 , n2191 , n2293 , n2294 );
and ( n2296 , n2187 , n2295 );
and ( n2297 , n2186 , n2295 );
or ( n2298 , n2188 , n2296 , n2297 );
and ( n2299 , n2184 , n2298 );
and ( n2300 , n2183 , n2298 );
or ( n2301 , n2185 , n2299 , n2300 );
and ( n2302 , n2181 , n2301 );
and ( n2303 , n2180 , n2301 );
or ( n2304 , n2182 , n2302 , n2303 );
and ( n2305 , n2178 , n2304 );
and ( n2306 , n2177 , n2304 );
or ( n2307 , n2179 , n2305 , n2306 );
and ( n2308 , n2175 , n2307 );
and ( n2309 , n2174 , n2307 );
or ( n2310 , n2176 , n2308 , n2309 );
and ( n2311 , n2172 , n2310 );
and ( n2312 , n2171 , n2310 );
or ( n2313 , n2173 , n2311 , n2312 );
and ( n2314 , n2169 , n2313 );
and ( n2315 , n2168 , n2313 );
or ( n2316 , n2170 , n2314 , n2315 );
and ( n2317 , n2166 , n2316 );
and ( n2318 , n2165 , n2316 );
or ( n2319 , n2167 , n2317 , n2318 );
and ( n2320 , n2163 , n2319 );
and ( n2321 , n2162 , n2319 );
or ( n2322 , n2164 , n2320 , n2321 );
and ( n2323 , n2160 , n2322 );
and ( n2324 , n2159 , n2322 );
or ( n2325 , n2161 , n2323 , n2324 );
and ( n2326 , n2157 , n2325 );
and ( n2327 , n2156 , n2325 );
or ( n2328 , n2158 , n2326 , n2327 );
and ( n2329 , n2154 , n2328 );
and ( n2330 , n2153 , n2328 );
or ( n2331 , n2155 , n2329 , n2330 );
and ( n2332 , n2151 , n2331 );
and ( n2333 , n2150 , n2331 );
or ( n2334 , n2152 , n2332 , n2333 );
and ( n2335 , n2148 , n2334 );
and ( n2336 , n2147 , n2334 );
or ( n2337 , n2149 , n2335 , n2336 );
and ( n2338 , n2145 , n2337 );
and ( n2339 , n2144 , n2337 );
or ( n2340 , n2146 , n2338 , n2339 );
and ( n2341 , n2142 , n2340 );
and ( n2342 , n2141 , n2340 );
or ( n2343 , n2143 , n2341 , n2342 );
and ( n2344 , n2139 , n2343 );
and ( n2345 , n2138 , n2343 );
or ( n2346 , n2140 , n2344 , n2345 );
and ( n2347 , n2136 , n2346 );
and ( n2348 , n2135 , n2346 );
or ( n2349 , n2137 , n2347 , n2348 );
and ( n2350 , n2133 , n2349 );
and ( n2351 , n2132 , n2349 );
or ( n2352 , n2134 , n2350 , n2351 );
and ( n2353 , n2130 , n2352 );
and ( n2354 , n2129 , n2352 );
or ( n2355 , n2131 , n2353 , n2354 );
and ( n2356 , n2127 , n2355 );
and ( n2357 , n2126 , n2355 );
or ( n2358 , n2128 , n2356 , n2357 );
and ( n2359 , n2124 , n2358 );
and ( n2360 , n2123 , n2358 );
or ( n2361 , n2125 , n2359 , n2360 );
and ( n2362 , n2121 , n2361 );
and ( n2363 , n2120 , n2361 );
or ( n2364 , n2122 , n2362 , n2363 );
and ( n2365 , n2118 , n2364 );
and ( n2366 , n2117 , n2364 );
or ( n2367 , n2119 , n2365 , n2366 );
and ( n2368 , n2115 , n2367 );
and ( n2369 , n2114 , n2367 );
or ( n2370 , n2116 , n2368 , n2369 );
and ( n2371 , n2112 , n2370 );
and ( n2372 , n2111 , n2370 );
or ( n2373 , n2113 , n2371 , n2372 );
and ( n2374 , n2109 , n2373 );
and ( n2375 , n2108 , n2373 );
or ( n2376 , n2110 , n2374 , n2375 );
and ( n2377 , n2106 , n2376 );
and ( n2378 , n2105 , n2376 );
or ( n2379 , n2107 , n2377 , n2378 );
and ( n2380 , n2103 , n2379 );
and ( n2381 , n2102 , n2379 );
or ( n2382 , n2104 , n2380 , n2381 );
and ( n2383 , n2100 , n2382 );
and ( n2384 , n2099 , n2382 );
or ( n2385 , n2101 , n2383 , n2384 );
and ( n2386 , n2097 , n2385 );
and ( n2387 , n2096 , n2385 );
or ( n2388 , n2098 , n2386 , n2387 );
and ( n2389 , n2094 , n2388 );
and ( n2390 , n2093 , n2388 );
or ( n2391 , n2095 , n2389 , n2390 );
and ( n2392 , n2091 , n2391 );
and ( n2393 , n2090 , n2391 );
or ( n2394 , n2092 , n2392 , n2393 );
and ( n2395 , n2088 , n2394 );
and ( n2396 , n2087 , n2394 );
or ( n2397 , n2089 , n2395 , n2396 );
and ( n2398 , n2085 , n2397 );
and ( n2399 , n2084 , n2397 );
or ( n2400 , n2086 , n2398 , n2399 );
and ( n2401 , n2082 , n2400 );
and ( n2402 , n2081 , n2400 );
or ( n2403 , n2083 , n2401 , n2402 );
and ( n2404 , n2079 , n2403 );
and ( n2405 , n2078 , n2403 );
or ( n2406 , n2080 , n2404 , n2405 );
and ( n2407 , n2076 , n2406 );
and ( n2408 , n2075 , n2406 );
or ( n2409 , n2077 , n2407 , n2408 );
and ( n2410 , n2073 , n2409 );
and ( n2411 , n2072 , n2409 );
or ( n2412 , n2074 , n2410 , n2411 );
and ( n2413 , n2070 , n2412 );
and ( n2414 , n2069 , n2412 );
or ( n2415 , n2071 , n2413 , n2414 );
and ( n2416 , n2067 , n2415 );
and ( n2417 , n2066 , n2415 );
or ( n2418 , n2068 , n2416 , n2417 );
and ( n2419 , n2064 , n2418 );
and ( n2420 , n2063 , n2418 );
or ( n2421 , n2065 , n2419 , n2420 );
and ( n2422 , n2061 , n2421 );
and ( n2423 , n2060 , n2421 );
or ( n2424 , n2062 , n2422 , n2423 );
and ( n2425 , n2058 , n2424 );
and ( n2426 , n2057 , n2424 );
or ( n2427 , n2059 , n2425 , n2426 );
and ( n2428 , n2055 , n2427 );
and ( n2429 , n2054 , n2427 );
or ( n2430 , n2056 , n2428 , n2429 );
and ( n2431 , n2052 , n2430 );
and ( n2432 , n2051 , n2430 );
or ( n2433 , n2053 , n2431 , n2432 );
and ( n2434 , n2049 , n2433 );
and ( n2435 , n2048 , n2433 );
or ( n2436 , n2050 , n2434 , n2435 );
and ( n2437 , n2046 , n2436 );
and ( n2438 , n2045 , n2436 );
or ( n2439 , n2047 , n2437 , n2438 );
and ( n2440 , n2043 , n2439 );
and ( n2441 , n2042 , n2439 );
or ( n2442 , n2044 , n2440 , n2441 );
and ( n2443 , n2040 , n2442 );
and ( n2444 , n2039 , n2442 );
or ( n2445 , n2041 , n2443 , n2444 );
and ( n2446 , n2037 , n2445 );
and ( n2447 , n2036 , n2445 );
or ( n2448 , n2038 , n2446 , n2447 );
and ( n2449 , n2034 , n2448 );
and ( n2450 , n2033 , n2448 );
or ( n2451 , n2035 , n2449 , n2450 );
and ( n2452 , n2031 , n2451 );
and ( n2453 , n2030 , n2451 );
or ( n2454 , n2032 , n2452 , n2453 );
and ( n2455 , n2028 , n2454 );
and ( n2456 , n2027 , n2454 );
or ( n2457 , n2029 , n2455 , n2456 );
and ( n2458 , n2025 , n2457 );
and ( n2459 , n2024 , n2457 );
or ( n2460 , n2026 , n2458 , n2459 );
and ( n2461 , n2022 , n2460 );
and ( n2462 , n2021 , n2460 );
or ( n2463 , n2023 , n2461 , n2462 );
and ( n2464 , n2019 , n2463 );
and ( n2465 , n2018 , n2463 );
or ( n2466 , n2020 , n2464 , n2465 );
and ( n2467 , n2016 , n2466 );
and ( n2468 , n2015 , n2466 );
or ( n2469 , n2017 , n2467 , n2468 );
and ( n2470 , n2013 , n2469 );
and ( n2471 , n2012 , n2469 );
or ( n2472 , n2014 , n2470 , n2471 );
and ( n2473 , n2010 , n2472 );
and ( n2474 , n2009 , n2472 );
or ( n2475 , n2011 , n2473 , n2474 );
and ( n2476 , n2007 , n2475 );
and ( n2477 , n2006 , n2475 );
or ( n2478 , n2008 , n2476 , n2477 );
and ( n2479 , n2004 , n2478 );
and ( n2480 , n2003 , n2478 );
or ( n2481 , n2005 , n2479 , n2480 );
and ( n2482 , n2001 , n2481 );
and ( n2483 , n2000 , n2481 );
or ( n2484 , n2002 , n2482 , n2483 );
and ( n2485 , n1998 , n2484 );
and ( n2486 , n1997 , n2484 );
or ( n2487 , n1999 , n2485 , n2486 );
and ( n2488 , n1995 , n2487 );
and ( n2489 , n1994 , n2487 );
or ( n2490 , n1996 , n2488 , n2489 );
and ( n2491 , n1992 , n2490 );
and ( n2492 , n1991 , n2490 );
or ( n2493 , n1993 , n2491 , n2492 );
and ( n2494 , n1989 , n2493 );
and ( n2495 , n1988 , n2493 );
or ( n2496 , n1990 , n2494 , n2495 );
and ( n2497 , n1986 , n2496 );
and ( n2498 , n1985 , n2496 );
or ( n2499 , n1987 , n2497 , n2498 );
and ( n2500 , n1983 , n2499 );
and ( n2501 , n1982 , n2499 );
or ( n2502 , n1984 , n2500 , n2501 );
and ( n2503 , n1980 , n2502 );
and ( n2504 , n1979 , n2502 );
or ( n2505 , n1981 , n2503 , n2504 );
and ( n2506 , n1977 , n2505 );
and ( n2507 , n1976 , n2505 );
or ( n2508 , n1978 , n2506 , n2507 );
and ( n2509 , n1974 , n2508 );
and ( n2510 , n1973 , n2508 );
or ( n2511 , n1975 , n2509 , n2510 );
and ( n2512 , n1971 , n2511 );
and ( n2513 , n1970 , n2511 );
or ( n2514 , n1972 , n2512 , n2513 );
and ( n2515 , n1968 , n2514 );
and ( n2516 , n1967 , n2514 );
or ( n2517 , n1969 , n2515 , n2516 );
and ( n2518 , n1965 , n2517 );
and ( n2519 , n1964 , n2517 );
or ( n2520 , n1966 , n2518 , n2519 );
and ( n2521 , n1962 , n2520 );
and ( n2522 , n1961 , n2520 );
or ( n2523 , n1963 , n2521 , n2522 );
and ( n2524 , n1959 , n2523 );
and ( n2525 , n1958 , n2523 );
or ( n2526 , n1960 , n2524 , n2525 );
and ( n2527 , n1956 , n2526 );
and ( n2528 , n1955 , n2526 );
or ( n2529 , n1957 , n2527 , n2528 );
and ( n2530 , n1953 , n2529 );
and ( n2531 , n1952 , n2529 );
or ( n2532 , n1954 , n2530 , n2531 );
and ( n2533 , n1950 , n2532 );
and ( n2534 , n1949 , n2532 );
or ( n2535 , n1951 , n2533 , n2534 );
and ( n2536 , n1947 , n2535 );
and ( n2537 , n1946 , n2535 );
or ( n2538 , n1948 , n2536 , n2537 );
and ( n2539 , n1944 , n2538 );
and ( n2540 , n1943 , n2538 );
or ( n2541 , n1945 , n2539 , n2540 );
and ( n2542 , n1941 , n2541 );
and ( n2543 , n1940 , n2541 );
or ( n2544 , n1942 , n2542 , n2543 );
and ( n2545 , n1938 , n2544 );
and ( n2546 , n1937 , n2544 );
or ( n2547 , n1939 , n2545 , n2546 );
and ( n2548 , n1935 , n2547 );
and ( n2549 , n1934 , n2547 );
or ( n2550 , n1936 , n2548 , n2549 );
and ( n2551 , n1932 , n2550 );
and ( n2552 , n1931 , n2550 );
or ( n2553 , n1933 , n2551 , n2552 );
and ( n2554 , n1929 , n2553 );
and ( n2555 , n1928 , n2553 );
or ( n2556 , n1930 , n2554 , n2555 );
and ( n2557 , n1926 , n2556 );
and ( n2558 , n1925 , n2556 );
or ( n2559 , n1927 , n2557 , n2558 );
and ( n2560 , n1923 , n2559 );
and ( n2561 , n1922 , n2559 );
or ( n2562 , n1924 , n2560 , n2561 );
and ( n2563 , n1920 , n2562 );
and ( n2564 , n1919 , n2562 );
or ( n2565 , n1921 , n2563 , n2564 );
and ( n2566 , n1917 , n2565 );
and ( n2567 , n1916 , n2565 );
or ( n2568 , n1918 , n2566 , n2567 );
and ( n2569 , n1914 , n2568 );
and ( n2570 , n1913 , n2568 );
or ( n2571 , n1915 , n2569 , n2570 );
and ( n2572 , n1911 , n2571 );
and ( n2573 , n1910 , n2571 );
or ( n2574 , n1912 , n2572 , n2573 );
and ( n2575 , n1908 , n2574 );
and ( n2576 , n1907 , n2574 );
or ( n2577 , n1909 , n2575 , n2576 );
and ( n2578 , n1905 , n2577 );
and ( n2579 , n1904 , n2577 );
or ( n2580 , n1906 , n2578 , n2579 );
and ( n2581 , n1902 , n2580 );
and ( n2582 , n1901 , n2580 );
or ( n2583 , n1903 , n2581 , n2582 );
and ( n2584 , n1899 , n2583 );
and ( n2585 , n1898 , n2583 );
or ( n2586 , n1900 , n2584 , n2585 );
and ( n2587 , n1896 , n2586 );
and ( n2588 , n1895 , n2586 );
or ( n2589 , n1897 , n2587 , n2588 );
and ( n2590 , n1893 , n2589 );
and ( n2591 , n1892 , n2589 );
or ( n2592 , n1894 , n2590 , n2591 );
and ( n2593 , n1890 , n2592 );
and ( n2594 , n1889 , n2592 );
or ( n2595 , n1891 , n2593 , n2594 );
and ( n2596 , n1887 , n2595 );
and ( n2597 , n1886 , n2595 );
or ( n2598 , n1888 , n2596 , n2597 );
and ( n2599 , n1884 , n2598 );
and ( n2600 , n1883 , n2598 );
or ( n2601 , n1885 , n2599 , n2600 );
and ( n2602 , n1881 , n2601 );
and ( n2603 , n1880 , n2601 );
or ( n2604 , n1882 , n2602 , n2603 );
and ( n2605 , n1878 , n2604 );
and ( n2606 , n1877 , n2604 );
or ( n2607 , n1879 , n2605 , n2606 );
and ( n2608 , n1875 , n2607 );
and ( n2609 , n1874 , n2607 );
or ( n2610 , n1876 , n2608 , n2609 );
and ( n2611 , n1872 , n2610 );
and ( n2612 , n1871 , n2610 );
or ( n2613 , n1873 , n2611 , n2612 );
and ( n2614 , n1869 , n2613 );
and ( n2615 , n1868 , n2613 );
or ( n2616 , n1870 , n2614 , n2615 );
and ( n2617 , n1866 , n2616 );
and ( n2618 , n1865 , n2616 );
or ( n2619 , n1867 , n2617 , n2618 );
and ( n2620 , n1863 , n2619 );
and ( n2621 , n1862 , n2619 );
or ( n2622 , n1864 , n2620 , n2621 );
and ( n2623 , n1860 , n2622 );
and ( n2624 , n1859 , n2622 );
or ( n2625 , n1861 , n2623 , n2624 );
and ( n2626 , n1857 , n2625 );
and ( n2627 , n1856 , n2625 );
or ( n2628 , n1858 , n2626 , n2627 );
and ( n2629 , n1854 , n2628 );
and ( n2630 , n1853 , n2628 );
or ( n2631 , n1855 , n2629 , n2630 );
and ( n2632 , n1851 , n2631 );
and ( n2633 , n1850 , n2631 );
or ( n2634 , n1852 , n2632 , n2633 );
and ( n2635 , n1848 , n2634 );
and ( n2636 , n1847 , n2634 );
or ( n2637 , n1849 , n2635 , n2636 );
and ( n2638 , n1845 , n2637 );
and ( n2639 , n1844 , n2637 );
or ( n2640 , n1846 , n2638 , n2639 );
and ( n2641 , n1842 , n2640 );
and ( n2642 , n1841 , n2640 );
or ( n2643 , n1843 , n2641 , n2642 );
and ( n2644 , n1839 , n2643 );
and ( n2645 , n1838 , n2643 );
or ( n2646 , n1840 , n2644 , n2645 );
and ( n2647 , n1836 , n2646 );
and ( n2648 , n1835 , n2646 );
or ( n2649 , n1837 , n2647 , n2648 );
and ( n2650 , n1833 , n2649 );
and ( n2651 , n1832 , n2649 );
or ( n2652 , n1834 , n2650 , n2651 );
and ( n2653 , n1830 , n2652 );
and ( n2654 , n1829 , n2652 );
or ( n2655 , n1831 , n2653 , n2654 );
and ( n2656 , n1827 , n2655 );
and ( n2657 , n1826 , n2655 );
or ( n2658 , n1828 , n2656 , n2657 );
and ( n2659 , n1824 , n2658 );
and ( n2660 , n1823 , n2658 );
or ( n2661 , n1825 , n2659 , n2660 );
and ( n2662 , n1821 , n2661 );
and ( n2663 , n1820 , n2661 );
or ( n2664 , n1822 , n2662 , n2663 );
and ( n2665 , n1818 , n2664 );
and ( n2666 , n1817 , n2664 );
or ( n2667 , n1819 , n2665 , n2666 );
and ( n2668 , n1815 , n2667 );
and ( n2669 , n1814 , n2667 );
or ( n2670 , n1816 , n2668 , n2669 );
and ( n2671 , n1812 , n2670 );
and ( n2672 , n1811 , n2670 );
or ( n2673 , n1813 , n2671 , n2672 );
and ( n2674 , n1809 , n2673 );
and ( n2675 , n1808 , n2673 );
or ( n2676 , n1810 , n2674 , n2675 );
and ( n2677 , n1806 , n2676 );
and ( n2678 , n1805 , n2676 );
or ( n2679 , n1807 , n2677 , n2678 );
and ( n2680 , n1803 , n2679 );
and ( n2681 , n1802 , n2679 );
or ( n2682 , n1804 , n2680 , n2681 );
and ( n2683 , n1800 , n2682 );
and ( n2684 , n1799 , n2682 );
or ( n2685 , n1801 , n2683 , n2684 );
and ( n2686 , n1797 , n2685 );
and ( n2687 , n1796 , n2685 );
or ( n2688 , n1798 , n2686 , n2687 );
and ( n2689 , n1794 , n2688 );
and ( n2690 , n1793 , n2688 );
or ( n2691 , n1795 , n2689 , n2690 );
and ( n2692 , n1791 , n2691 );
and ( n2693 , n1790 , n2691 );
or ( n2694 , n1792 , n2692 , n2693 );
and ( n2695 , n1788 , n2694 );
and ( n2696 , n1787 , n2694 );
or ( n2697 , n1789 , n2695 , n2696 );
and ( n2698 , n1785 , n2697 );
and ( n2699 , n1784 , n2697 );
or ( n2700 , n1786 , n2698 , n2699 );
and ( n2701 , n1782 , n2700 );
and ( n2702 , n1781 , n2700 );
or ( n2703 , n1783 , n2701 , n2702 );
and ( n2704 , n1779 , n2703 );
and ( n2705 , n1778 , n2703 );
or ( n2706 , n1780 , n2704 , n2705 );
and ( n2707 , n1776 , n2706 );
and ( n2708 , n1775 , n2706 );
or ( n2709 , n1777 , n2707 , n2708 );
and ( n2710 , n1773 , n2709 );
and ( n2711 , n1772 , n2709 );
or ( n2712 , n1774 , n2710 , n2711 );
and ( n2713 , n1770 , n2712 );
and ( n2714 , n1769 , n2712 );
or ( n2715 , n1771 , n2713 , n2714 );
and ( n2716 , n1767 , n2715 );
and ( n2717 , n1766 , n2715 );
or ( n2718 , n1768 , n2716 , n2717 );
and ( n2719 , n1764 , n2718 );
and ( n2720 , n1763 , n2718 );
or ( n2721 , n1765 , n2719 , n2720 );
and ( n2722 , n1761 , n2721 );
and ( n2723 , n1760 , n2721 );
or ( n2724 , n1762 , n2722 , n2723 );
and ( n2725 , n1758 , n2724 );
and ( n2726 , n1757 , n2724 );
or ( n2727 , n1759 , n2725 , n2726 );
and ( n2728 , n1755 , n2727 );
and ( n2729 , n1754 , n2727 );
or ( n2730 , n1756 , n2728 , n2729 );
and ( n2731 , n1752 , n2730 );
and ( n2732 , n1751 , n2730 );
or ( n2733 , n1753 , n2731 , n2732 );
and ( n2734 , n1749 , n2733 );
and ( n2735 , n1748 , n2733 );
or ( n2736 , n1750 , n2734 , n2735 );
and ( n2737 , n1746 , n2736 );
and ( n2738 , n1745 , n2736 );
or ( n2739 , n1747 , n2737 , n2738 );
and ( n2740 , n1743 , n2739 );
and ( n2741 , n1742 , n2739 );
or ( n2742 , n1744 , n2740 , n2741 );
and ( n2743 , n1740 , n2742 );
and ( n2744 , n1739 , n2742 );
or ( n2745 , n1741 , n2743 , n2744 );
and ( n2746 , n1737 , n2745 );
and ( n2747 , n1736 , n2745 );
or ( n2748 , n1738 , n2746 , n2747 );
and ( n2749 , n1734 , n2748 );
and ( n2750 , n1733 , n2748 );
or ( n2751 , n1735 , n2749 , n2750 );
and ( n2752 , n1731 , n2751 );
and ( n2753 , n1730 , n2751 );
or ( n2754 , n1732 , n2752 , n2753 );
and ( n2755 , n1728 , n2754 );
and ( n2756 , n1727 , n2754 );
or ( n2757 , n1729 , n2755 , n2756 );
and ( n2758 , n1725 , n2757 );
and ( n2759 , n1724 , n2757 );
or ( n2760 , n1726 , n2758 , n2759 );
and ( n2761 , n1722 , n2760 );
and ( n2762 , n1721 , n2760 );
or ( n2763 , n1723 , n2761 , n2762 );
and ( n2764 , n1719 , n2763 );
and ( n2765 , n1718 , n2763 );
or ( n2766 , n1720 , n2764 , n2765 );
and ( n2767 , n1716 , n2766 );
and ( n2768 , n1715 , n2766 );
or ( n2769 , n1717 , n2767 , n2768 );
and ( n2770 , n1713 , n2769 );
and ( n2771 , n1712 , n2769 );
or ( n2772 , n1714 , n2770 , n2771 );
and ( n2773 , n1710 , n2772 );
and ( n2774 , n1709 , n2772 );
or ( n2775 , n1711 , n2773 , n2774 );
and ( n2776 , n1707 , n2775 );
and ( n2777 , n1706 , n2775 );
or ( n2778 , n1708 , n2776 , n2777 );
and ( n2779 , n1704 , n2778 );
and ( n2780 , n1703 , n2778 );
or ( n2781 , n1705 , n2779 , n2780 );
and ( n2782 , n1701 , n2781 );
and ( n2783 , n1700 , n2781 );
or ( n2784 , n1702 , n2782 , n2783 );
and ( n2785 , n1698 , n2784 );
and ( n2786 , n1697 , n2784 );
or ( n2787 , n1699 , n2785 , n2786 );
and ( n2788 , n1695 , n2787 );
and ( n2789 , n1694 , n2787 );
or ( n2790 , n1696 , n2788 , n2789 );
and ( n2791 , n1692 , n2790 );
and ( n2792 , n1691 , n2790 );
or ( n2793 , n1693 , n2791 , n2792 );
and ( n2794 , n1689 , n2793 );
and ( n2795 , n1688 , n2793 );
or ( n2796 , n1690 , n2794 , n2795 );
and ( n2797 , n1686 , n2796 );
and ( n2798 , n1685 , n2796 );
or ( n2799 , n1687 , n2797 , n2798 );
and ( n2800 , n1683 , n2799 );
and ( n2801 , n1682 , n2799 );
or ( n2802 , n1684 , n2800 , n2801 );
and ( n2803 , n1680 , n2802 );
and ( n2804 , n1679 , n2802 );
or ( n2805 , n1681 , n2803 , n2804 );
and ( n2806 , n1677 , n2805 );
and ( n2807 , n1676 , n2805 );
or ( n2808 , n1678 , n2806 , n2807 );
and ( n2809 , n1674 , n2808 );
and ( n2810 , n1673 , n2808 );
or ( n2811 , n1675 , n2809 , n2810 );
and ( n2812 , n1671 , n2811 );
and ( n2813 , n1670 , n2811 );
or ( n2814 , n1672 , n2812 , n2813 );
and ( n2815 , n1668 , n2814 );
and ( n2816 , n1667 , n2814 );
or ( n2817 , n1669 , n2815 , n2816 );
and ( n2818 , n1665 , n2817 );
and ( n2819 , n1664 , n2817 );
or ( n2820 , n1666 , n2818 , n2819 );
and ( n2821 , n1662 , n2820 );
and ( n2822 , n1661 , n2820 );
or ( n2823 , n1663 , n2821 , n2822 );
and ( n2824 , n1659 , n2823 );
and ( n2825 , n1658 , n2823 );
or ( n2826 , n1660 , n2824 , n2825 );
and ( n2827 , n1656 , n2826 );
and ( n2828 , n1655 , n2826 );
or ( n2829 , n1657 , n2827 , n2828 );
and ( n2830 , n1653 , n2829 );
and ( n2831 , n1652 , n2829 );
or ( n2832 , n1654 , n2830 , n2831 );
and ( n2833 , n1650 , n2832 );
and ( n2834 , n1649 , n2832 );
or ( n2835 , n1651 , n2833 , n2834 );
and ( n2836 , n1647 , n2835 );
and ( n2837 , n1646 , n2835 );
or ( n2838 , n1648 , n2836 , n2837 );
and ( n2839 , n1644 , n2838 );
and ( n2840 , n1643 , n2838 );
or ( n2841 , n1645 , n2839 , n2840 );
and ( n2842 , n1641 , n2841 );
and ( n2843 , n1640 , n2841 );
or ( n2844 , n1642 , n2842 , n2843 );
and ( n2845 , n1638 , n2844 );
and ( n2846 , n1637 , n2844 );
or ( n2847 , n1639 , n2845 , n2846 );
and ( n2848 , n1635 , n2847 );
and ( n2849 , n1634 , n2847 );
or ( n2850 , n1636 , n2848 , n2849 );
and ( n2851 , n1632 , n2850 );
and ( n2852 , n1631 , n2850 );
or ( n2853 , n1633 , n2851 , n2852 );
and ( n2854 , n1629 , n2853 );
and ( n2855 , n1628 , n2853 );
or ( n2856 , n1630 , n2854 , n2855 );
and ( n2857 , n1626 , n2856 );
and ( n2858 , n1625 , n2856 );
or ( n2859 , n1627 , n2857 , n2858 );
and ( n2860 , n1623 , n2859 );
and ( n2861 , n1622 , n2859 );
or ( n2862 , n1624 , n2860 , n2861 );
and ( n2863 , n1620 , n2862 );
and ( n2864 , n1619 , n2862 );
or ( n2865 , n1621 , n2863 , n2864 );
and ( n2866 , n1617 , n2865 );
and ( n2867 , n1616 , n2865 );
or ( n2868 , n1618 , n2866 , n2867 );
and ( n2869 , n1614 , n2868 );
and ( n2870 , n1613 , n2868 );
or ( n2871 , n1615 , n2869 , n2870 );
and ( n2872 , n1611 , n2871 );
and ( n2873 , n1610 , n2871 );
or ( n2874 , n1612 , n2872 , n2873 );
and ( n2875 , n1608 , n2874 );
and ( n2876 , n1607 , n2874 );
or ( n2877 , n1609 , n2875 , n2876 );
and ( n2878 , n1605 , n2877 );
and ( n2879 , n1604 , n2877 );
or ( n2880 , n1606 , n2878 , n2879 );
and ( n2881 , n1602 , n2880 );
and ( n2882 , n1601 , n2880 );
or ( n2883 , n1603 , n2881 , n2882 );
and ( n2884 , n1599 , n2883 );
and ( n2885 , n1598 , n2883 );
or ( n2886 , n1600 , n2884 , n2885 );
and ( n2887 , n1596 , n2886 );
and ( n2888 , n1595 , n2886 );
or ( n2889 , n1597 , n2887 , n2888 );
and ( n2890 , n1593 , n2889 );
and ( n2891 , n1592 , n2889 );
or ( n2892 , n1594 , n2890 , n2891 );
and ( n2893 , n1590 , n2892 );
and ( n2894 , n1589 , n2892 );
or ( n2895 , n1591 , n2893 , n2894 );
and ( n2896 , n1587 , n2895 );
and ( n2897 , n1586 , n2895 );
or ( n2898 , n1588 , n2896 , n2897 );
and ( n2899 , n1584 , n2898 );
and ( n2900 , n1583 , n2898 );
or ( n2901 , n1585 , n2899 , n2900 );
and ( n2902 , n1581 , n2901 );
and ( n2903 , n1580 , n2901 );
or ( n2904 , n1582 , n2902 , n2903 );
and ( n2905 , n1578 , n2904 );
and ( n2906 , n1577 , n2904 );
or ( n2907 , n1579 , n2905 , n2906 );
and ( n2908 , n1575 , n2907 );
and ( n2909 , n1574 , n2907 );
or ( n2910 , n1576 , n2908 , n2909 );
and ( n2911 , n1572 , n2910 );
and ( n2912 , n1571 , n2910 );
or ( n2913 , n1573 , n2911 , n2912 );
and ( n2914 , n1569 , n2913 );
and ( n2915 , n1568 , n2913 );
or ( n2916 , n1570 , n2914 , n2915 );
and ( n2917 , n1566 , n2916 );
and ( n2918 , n1565 , n2916 );
or ( n2919 , n1567 , n2917 , n2918 );
and ( n2920 , n1563 , n2919 );
and ( n2921 , n1562 , n2919 );
or ( n2922 , n1564 , n2920 , n2921 );
and ( n2923 , n1560 , n2922 );
and ( n2924 , n1559 , n2922 );
or ( n2925 , n1561 , n2923 , n2924 );
and ( n2926 , n1557 , n2925 );
and ( n2927 , n1556 , n2925 );
or ( n2928 , n1558 , n2926 , n2927 );
and ( n2929 , n1554 , n2928 );
and ( n2930 , n1553 , n2928 );
or ( n2931 , n1555 , n2929 , n2930 );
and ( n2932 , n1551 , n2931 );
and ( n2933 , n1550 , n2931 );
or ( n2934 , n1552 , n2932 , n2933 );
and ( n2935 , n1548 , n2934 );
and ( n2936 , n1547 , n2934 );
or ( n2937 , n1549 , n2935 , n2936 );
and ( n2938 , n1545 , n2937 );
and ( n2939 , n1544 , n2937 );
or ( n2940 , n1546 , n2938 , n2939 );
and ( n2941 , n1542 , n2940 );
and ( n2942 , n1541 , n2940 );
or ( n2943 , n1543 , n2941 , n2942 );
xor ( n2944 , n1540 , n2943 );
buf ( n2945 , n2944 );
xor ( n2946 , n1541 , n1542 );
xor ( n2947 , n2946 , n2940 );
buf ( n2948 , n2947 );
xor ( n2949 , n2945 , n2948 );
xor ( n2950 , n1544 , n1545 );
xor ( n2951 , n2950 , n2937 );
buf ( n2952 , n2951 );
xor ( n2953 , n1547 , n1548 );
xor ( n2954 , n2953 , n2934 );
buf ( n2955 , n2954 );
xor ( n2956 , n2952 , n2955 );
xor ( n2957 , n2949 , n2956 );
xor ( n2958 , n1550 , n1551 );
xor ( n2959 , n2958 , n2931 );
buf ( n2960 , n2959 );
xor ( n2961 , n1553 , n1554 );
xor ( n2962 , n2961 , n2928 );
buf ( n2963 , n2962 );
xor ( n2964 , n2960 , n2963 );
xor ( n2965 , n1556 , n1557 );
xor ( n2966 , n2965 , n2925 );
buf ( n2967 , n2966 );
xor ( n2968 , n1559 , n1560 );
xor ( n2969 , n2968 , n2922 );
buf ( n2970 , n2969 );
xor ( n2971 , n2967 , n2970 );
xor ( n2972 , n2964 , n2971 );
xor ( n2973 , n2957 , n2972 );
xor ( n2974 , n1562 , n1563 );
xor ( n2975 , n2974 , n2919 );
buf ( n2976 , n2975 );
xor ( n2977 , n1565 , n1566 );
xor ( n2978 , n2977 , n2916 );
buf ( n2979 , n2978 );
xor ( n2980 , n2976 , n2979 );
xor ( n2981 , n1568 , n1569 );
xor ( n2982 , n2981 , n2913 );
buf ( n2983 , n2982 );
xor ( n2984 , n1571 , n1572 );
xor ( n2985 , n2984 , n2910 );
buf ( n2986 , n2985 );
xor ( n2987 , n2983 , n2986 );
xor ( n2988 , n2980 , n2987 );
xor ( n2989 , n1574 , n1575 );
xor ( n2990 , n2989 , n2907 );
buf ( n2991 , n2990 );
xor ( n2992 , n1577 , n1578 );
xor ( n2993 , n2992 , n2904 );
buf ( n2994 , n2993 );
xor ( n2995 , n2991 , n2994 );
xor ( n2996 , n1580 , n1581 );
xor ( n2997 , n2996 , n2901 );
buf ( n2998 , n2997 );
xor ( n2999 , n1583 , n1584 );
xor ( n3000 , n2999 , n2898 );
buf ( n3001 , n3000 );
xor ( n3002 , n2998 , n3001 );
xor ( n3003 , n2995 , n3002 );
xor ( n3004 , n2988 , n3003 );
xor ( n3005 , n2973 , n3004 );
xor ( n3006 , n1586 , n1587 );
xor ( n3007 , n3006 , n2895 );
buf ( n3008 , n3007 );
xor ( n3009 , n1589 , n1590 );
xor ( n3010 , n3009 , n2892 );
buf ( n3011 , n3010 );
xor ( n3012 , n3008 , n3011 );
xor ( n3013 , n1592 , n1593 );
xor ( n3014 , n3013 , n2889 );
buf ( n3015 , n3014 );
xor ( n3016 , n1595 , n1596 );
xor ( n3017 , n3016 , n2886 );
buf ( n3018 , n3017 );
xor ( n3019 , n3015 , n3018 );
xor ( n3020 , n3012 , n3019 );
xor ( n3021 , n1598 , n1599 );
xor ( n3022 , n3021 , n2883 );
buf ( n3023 , n3022 );
xor ( n3024 , n1601 , n1602 );
xor ( n3025 , n3024 , n2880 );
buf ( n3026 , n3025 );
xor ( n3027 , n3023 , n3026 );
xor ( n3028 , n1604 , n1605 );
xor ( n3029 , n3028 , n2877 );
buf ( n3030 , n3029 );
xor ( n3031 , n1607 , n1608 );
xor ( n3032 , n3031 , n2874 );
buf ( n3033 , n3032 );
xor ( n3034 , n3030 , n3033 );
xor ( n3035 , n3027 , n3034 );
xor ( n3036 , n3020 , n3035 );
xor ( n3037 , n1610 , n1611 );
xor ( n3038 , n3037 , n2871 );
buf ( n3039 , n3038 );
xor ( n3040 , n1613 , n1614 );
xor ( n3041 , n3040 , n2868 );
buf ( n3042 , n3041 );
xor ( n3043 , n3039 , n3042 );
xor ( n3044 , n1616 , n1617 );
xor ( n3045 , n3044 , n2865 );
buf ( n3046 , n3045 );
xor ( n3047 , n1619 , n1620 );
xor ( n3048 , n3047 , n2862 );
buf ( n3049 , n3048 );
xor ( n3050 , n3046 , n3049 );
xor ( n3051 , n3043 , n3050 );
xor ( n3052 , n1622 , n1623 );
xor ( n3053 , n3052 , n2859 );
buf ( n3054 , n3053 );
xor ( n3055 , n1625 , n1626 );
xor ( n3056 , n3055 , n2856 );
buf ( n3057 , n3056 );
xor ( n3058 , n3054 , n3057 );
xor ( n3059 , n1628 , n1629 );
xor ( n3060 , n3059 , n2853 );
buf ( n3061 , n3060 );
xor ( n3062 , n1631 , n1632 );
xor ( n3063 , n3062 , n2850 );
buf ( n3064 , n3063 );
xor ( n3065 , n3061 , n3064 );
xor ( n3066 , n3058 , n3065 );
xor ( n3067 , n3051 , n3066 );
xor ( n3068 , n3036 , n3067 );
xor ( n3069 , n3005 , n3068 );
xor ( n3070 , n1634 , n1635 );
xor ( n3071 , n3070 , n2847 );
buf ( n3072 , n3071 );
xor ( n3073 , n1637 , n1638 );
xor ( n3074 , n3073 , n2844 );
buf ( n3075 , n3074 );
xor ( n3076 , n3072 , n3075 );
xor ( n3077 , n1640 , n1641 );
xor ( n3078 , n3077 , n2841 );
buf ( n3079 , n3078 );
xor ( n3080 , n1643 , n1644 );
xor ( n3081 , n3080 , n2838 );
buf ( n3082 , n3081 );
xor ( n3083 , n3079 , n3082 );
xor ( n3084 , n3076 , n3083 );
xor ( n3085 , n1646 , n1647 );
xor ( n3086 , n3085 , n2835 );
buf ( n3087 , n3086 );
xor ( n3088 , n1649 , n1650 );
xor ( n3089 , n3088 , n2832 );
buf ( n3090 , n3089 );
xor ( n3091 , n3087 , n3090 );
xor ( n3092 , n1652 , n1653 );
xor ( n3093 , n3092 , n2829 );
buf ( n3094 , n3093 );
xor ( n3095 , n1655 , n1656 );
xor ( n3096 , n3095 , n2826 );
buf ( n3097 , n3096 );
xor ( n3098 , n3094 , n3097 );
xor ( n3099 , n3091 , n3098 );
xor ( n3100 , n3084 , n3099 );
xor ( n3101 , n1658 , n1659 );
xor ( n3102 , n3101 , n2823 );
buf ( n3103 , n3102 );
xor ( n3104 , n1661 , n1662 );
xor ( n3105 , n3104 , n2820 );
buf ( n3106 , n3105 );
xor ( n3107 , n3103 , n3106 );
xor ( n3108 , n1664 , n1665 );
xor ( n3109 , n3108 , n2817 );
buf ( n3110 , n3109 );
xor ( n3111 , n1667 , n1668 );
xor ( n3112 , n3111 , n2814 );
buf ( n3113 , n3112 );
xor ( n3114 , n3110 , n3113 );
xor ( n3115 , n3107 , n3114 );
xor ( n3116 , n1670 , n1671 );
xor ( n3117 , n3116 , n2811 );
buf ( n3118 , n3117 );
xor ( n3119 , n1673 , n1674 );
xor ( n3120 , n3119 , n2808 );
buf ( n3121 , n3120 );
xor ( n3122 , n3118 , n3121 );
xor ( n3123 , n1676 , n1677 );
xor ( n3124 , n3123 , n2805 );
buf ( n3125 , n3124 );
xor ( n3126 , n1679 , n1680 );
xor ( n3127 , n3126 , n2802 );
buf ( n3128 , n3127 );
xor ( n3129 , n3125 , n3128 );
xor ( n3130 , n3122 , n3129 );
xor ( n3131 , n3115 , n3130 );
xor ( n3132 , n3100 , n3131 );
xor ( n3133 , n1682 , n1683 );
xor ( n3134 , n3133 , n2799 );
buf ( n3135 , n3134 );
xor ( n3136 , n1685 , n1686 );
xor ( n3137 , n3136 , n2796 );
buf ( n3138 , n3137 );
xor ( n3139 , n3135 , n3138 );
xor ( n3140 , n1688 , n1689 );
xor ( n3141 , n3140 , n2793 );
buf ( n3142 , n3141 );
xor ( n3143 , n1691 , n1692 );
xor ( n3144 , n3143 , n2790 );
buf ( n3145 , n3144 );
xor ( n3146 , n3142 , n3145 );
xor ( n3147 , n3139 , n3146 );
xor ( n3148 , n1694 , n1695 );
xor ( n3149 , n3148 , n2787 );
buf ( n3150 , n3149 );
xor ( n3151 , n1697 , n1698 );
xor ( n3152 , n3151 , n2784 );
buf ( n3153 , n3152 );
xor ( n3154 , n3150 , n3153 );
xor ( n3155 , n1700 , n1701 );
xor ( n3156 , n3155 , n2781 );
buf ( n3157 , n3156 );
xor ( n3158 , n1703 , n1704 );
xor ( n3159 , n3158 , n2778 );
buf ( n3160 , n3159 );
xor ( n3161 , n3157 , n3160 );
xor ( n3162 , n3154 , n3161 );
xor ( n3163 , n3147 , n3162 );
xor ( n3164 , n1706 , n1707 );
xor ( n3165 , n3164 , n2775 );
buf ( n3166 , n3165 );
xor ( n3167 , n1709 , n1710 );
xor ( n3168 , n3167 , n2772 );
buf ( n3169 , n3168 );
xor ( n3170 , n3166 , n3169 );
xor ( n3171 , n1712 , n1713 );
xor ( n3172 , n3171 , n2769 );
buf ( n3173 , n3172 );
xor ( n3174 , n1715 , n1716 );
xor ( n3175 , n3174 , n2766 );
buf ( n3176 , n3175 );
xor ( n3177 , n3173 , n3176 );
xor ( n3178 , n3170 , n3177 );
xor ( n3179 , n1718 , n1719 );
xor ( n3180 , n3179 , n2763 );
buf ( n3181 , n3180 );
xor ( n3182 , n1721 , n1722 );
xor ( n3183 , n3182 , n2760 );
buf ( n3184 , n3183 );
xor ( n3185 , n3181 , n3184 );
xor ( n3186 , n1724 , n1725 );
xor ( n3187 , n3186 , n2757 );
buf ( n3188 , n3187 );
xor ( n3189 , n1727 , n1728 );
xor ( n3190 , n3189 , n2754 );
buf ( n3191 , n3190 );
xor ( n3192 , n3188 , n3191 );
xor ( n3193 , n3185 , n3192 );
xor ( n3194 , n3178 , n3193 );
xor ( n3195 , n3163 , n3194 );
xor ( n3196 , n3132 , n3195 );
xor ( n3197 , n3069 , n3196 );
xor ( n3198 , n1730 , n1731 );
xor ( n3199 , n3198 , n2751 );
buf ( n3200 , n3199 );
xor ( n3201 , n1733 , n1734 );
xor ( n3202 , n3201 , n2748 );
buf ( n3203 , n3202 );
xor ( n3204 , n3200 , n3203 );
xor ( n3205 , n1736 , n1737 );
xor ( n3206 , n3205 , n2745 );
buf ( n3207 , n3206 );
xor ( n3208 , n1739 , n1740 );
xor ( n3209 , n3208 , n2742 );
buf ( n3210 , n3209 );
xor ( n3211 , n3207 , n3210 );
xor ( n3212 , n3204 , n3211 );
xor ( n3213 , n1742 , n1743 );
xor ( n3214 , n3213 , n2739 );
buf ( n3215 , n3214 );
xor ( n3216 , n1745 , n1746 );
xor ( n3217 , n3216 , n2736 );
buf ( n3218 , n3217 );
xor ( n3219 , n3215 , n3218 );
xor ( n3220 , n1748 , n1749 );
xor ( n3221 , n3220 , n2733 );
buf ( n3222 , n3221 );
xor ( n3223 , n1751 , n1752 );
xor ( n3224 , n3223 , n2730 );
buf ( n3225 , n3224 );
xor ( n3226 , n3222 , n3225 );
xor ( n3227 , n3219 , n3226 );
xor ( n3228 , n3212 , n3227 );
xor ( n3229 , n1754 , n1755 );
xor ( n3230 , n3229 , n2727 );
buf ( n3231 , n3230 );
xor ( n3232 , n1757 , n1758 );
xor ( n3233 , n3232 , n2724 );
buf ( n3234 , n3233 );
xor ( n3235 , n3231 , n3234 );
xor ( n3236 , n1760 , n1761 );
xor ( n3237 , n3236 , n2721 );
buf ( n3238 , n3237 );
xor ( n3239 , n1763 , n1764 );
xor ( n3240 , n3239 , n2718 );
buf ( n3241 , n3240 );
xor ( n3242 , n3238 , n3241 );
xor ( n3243 , n3235 , n3242 );
xor ( n3244 , n1766 , n1767 );
xor ( n3245 , n3244 , n2715 );
buf ( n3246 , n3245 );
xor ( n3247 , n1769 , n1770 );
xor ( n3248 , n3247 , n2712 );
buf ( n3249 , n3248 );
xor ( n3250 , n3246 , n3249 );
xor ( n3251 , n1772 , n1773 );
xor ( n3252 , n3251 , n2709 );
buf ( n3253 , n3252 );
xor ( n3254 , n1775 , n1776 );
xor ( n3255 , n3254 , n2706 );
buf ( n3256 , n3255 );
xor ( n3257 , n3253 , n3256 );
xor ( n3258 , n3250 , n3257 );
xor ( n3259 , n3243 , n3258 );
xor ( n3260 , n3228 , n3259 );
xor ( n3261 , n1778 , n1779 );
xor ( n3262 , n3261 , n2703 );
buf ( n3263 , n3262 );
xor ( n3264 , n1781 , n1782 );
xor ( n3265 , n3264 , n2700 );
buf ( n3266 , n3265 );
xor ( n3267 , n3263 , n3266 );
xor ( n3268 , n1784 , n1785 );
xor ( n3269 , n3268 , n2697 );
buf ( n3270 , n3269 );
xor ( n3271 , n1787 , n1788 );
xor ( n3272 , n3271 , n2694 );
buf ( n3273 , n3272 );
xor ( n3274 , n3270 , n3273 );
xor ( n3275 , n3267 , n3274 );
xor ( n3276 , n1790 , n1791 );
xor ( n3277 , n3276 , n2691 );
buf ( n3278 , n3277 );
xor ( n3279 , n1793 , n1794 );
xor ( n3280 , n3279 , n2688 );
buf ( n3281 , n3280 );
xor ( n3282 , n3278 , n3281 );
xor ( n3283 , n1796 , n1797 );
xor ( n3284 , n3283 , n2685 );
buf ( n3285 , n3284 );
xor ( n3286 , n1799 , n1800 );
xor ( n3287 , n3286 , n2682 );
buf ( n3288 , n3287 );
xor ( n3289 , n3285 , n3288 );
xor ( n3290 , n3282 , n3289 );
xor ( n3291 , n3275 , n3290 );
xor ( n3292 , n1802 , n1803 );
xor ( n3293 , n3292 , n2679 );
buf ( n3294 , n3293 );
xor ( n3295 , n1805 , n1806 );
xor ( n3296 , n3295 , n2676 );
buf ( n3297 , n3296 );
xor ( n3298 , n3294 , n3297 );
xor ( n3299 , n1808 , n1809 );
xor ( n3300 , n3299 , n2673 );
buf ( n3301 , n3300 );
xor ( n3302 , n1811 , n1812 );
xor ( n3303 , n3302 , n2670 );
buf ( n3304 , n3303 );
xor ( n3305 , n3301 , n3304 );
xor ( n3306 , n3298 , n3305 );
xor ( n3307 , n1814 , n1815 );
xor ( n3308 , n3307 , n2667 );
buf ( n3309 , n3308 );
xor ( n3310 , n1817 , n1818 );
xor ( n3311 , n3310 , n2664 );
buf ( n3312 , n3311 );
xor ( n3313 , n3309 , n3312 );
xor ( n3314 , n1820 , n1821 );
xor ( n3315 , n3314 , n2661 );
buf ( n3316 , n3315 );
xor ( n3317 , n1823 , n1824 );
xor ( n3318 , n3317 , n2658 );
buf ( n3319 , n3318 );
xor ( n3320 , n3316 , n3319 );
xor ( n3321 , n3313 , n3320 );
xor ( n3322 , n3306 , n3321 );
xor ( n3323 , n3291 , n3322 );
xor ( n3324 , n3260 , n3323 );
xor ( n3325 , n1826 , n1827 );
xor ( n3326 , n3325 , n2655 );
buf ( n3327 , n3326 );
xor ( n3328 , n1829 , n1830 );
xor ( n3329 , n3328 , n2652 );
buf ( n3330 , n3329 );
xor ( n3331 , n3327 , n3330 );
xor ( n3332 , n1832 , n1833 );
xor ( n3333 , n3332 , n2649 );
buf ( n3334 , n3333 );
xor ( n3335 , n1835 , n1836 );
xor ( n3336 , n3335 , n2646 );
buf ( n3337 , n3336 );
xor ( n3338 , n3334 , n3337 );
xor ( n3339 , n3331 , n3338 );
xor ( n3340 , n1838 , n1839 );
xor ( n3341 , n3340 , n2643 );
buf ( n3342 , n3341 );
xor ( n3343 , n1841 , n1842 );
xor ( n3344 , n3343 , n2640 );
buf ( n3345 , n3344 );
xor ( n3346 , n3342 , n3345 );
xor ( n3347 , n1844 , n1845 );
xor ( n3348 , n3347 , n2637 );
buf ( n3349 , n3348 );
xor ( n3350 , n1847 , n1848 );
xor ( n3351 , n3350 , n2634 );
buf ( n3352 , n3351 );
xor ( n3353 , n3349 , n3352 );
xor ( n3354 , n3346 , n3353 );
xor ( n3355 , n3339 , n3354 );
xor ( n3356 , n1850 , n1851 );
xor ( n3357 , n3356 , n2631 );
buf ( n3358 , n3357 );
xor ( n3359 , n1853 , n1854 );
xor ( n3360 , n3359 , n2628 );
buf ( n3361 , n3360 );
xor ( n3362 , n3358 , n3361 );
xor ( n3363 , n1856 , n1857 );
xor ( n3364 , n3363 , n2625 );
buf ( n3365 , n3364 );
xor ( n3366 , n1859 , n1860 );
xor ( n3367 , n3366 , n2622 );
buf ( n3368 , n3367 );
xor ( n3369 , n3365 , n3368 );
xor ( n3370 , n3362 , n3369 );
xor ( n3371 , n1862 , n1863 );
xor ( n3372 , n3371 , n2619 );
buf ( n3373 , n3372 );
xor ( n3374 , n1865 , n1866 );
xor ( n3375 , n3374 , n2616 );
buf ( n3376 , n3375 );
xor ( n3377 , n3373 , n3376 );
xor ( n3378 , n1868 , n1869 );
xor ( n3379 , n3378 , n2613 );
buf ( n3380 , n3379 );
xor ( n3381 , n1871 , n1872 );
xor ( n3382 , n3381 , n2610 );
buf ( n3383 , n3382 );
xor ( n3384 , n3380 , n3383 );
xor ( n3385 , n3377 , n3384 );
xor ( n3386 , n3370 , n3385 );
xor ( n3387 , n3355 , n3386 );
xor ( n3388 , n1874 , n1875 );
xor ( n3389 , n3388 , n2607 );
buf ( n3390 , n3389 );
xor ( n3391 , n1877 , n1878 );
xor ( n3392 , n3391 , n2604 );
buf ( n3393 , n3392 );
xor ( n3394 , n3390 , n3393 );
xor ( n3395 , n1880 , n1881 );
xor ( n3396 , n3395 , n2601 );
buf ( n3397 , n3396 );
xor ( n3398 , n1883 , n1884 );
xor ( n3399 , n3398 , n2598 );
buf ( n3400 , n3399 );
xor ( n3401 , n3397 , n3400 );
xor ( n3402 , n3394 , n3401 );
xor ( n3403 , n1886 , n1887 );
xor ( n3404 , n3403 , n2595 );
buf ( n3405 , n3404 );
xor ( n3406 , n1889 , n1890 );
xor ( n3407 , n3406 , n2592 );
buf ( n3408 , n3407 );
xor ( n3409 , n3405 , n3408 );
xor ( n3410 , n1892 , n1893 );
xor ( n3411 , n3410 , n2589 );
buf ( n3412 , n3411 );
xor ( n3413 , n1895 , n1896 );
xor ( n3414 , n3413 , n2586 );
buf ( n3415 , n3414 );
xor ( n3416 , n3412 , n3415 );
xor ( n3417 , n3409 , n3416 );
xor ( n3418 , n3402 , n3417 );
xor ( n3419 , n1898 , n1899 );
xor ( n3420 , n3419 , n2583 );
buf ( n3421 , n3420 );
xor ( n3422 , n1901 , n1902 );
xor ( n3423 , n3422 , n2580 );
buf ( n3424 , n3423 );
xor ( n3425 , n3421 , n3424 );
xor ( n3426 , n1904 , n1905 );
xor ( n3427 , n3426 , n2577 );
buf ( n3428 , n3427 );
xor ( n3429 , n1907 , n1908 );
xor ( n3430 , n3429 , n2574 );
buf ( n3431 , n3430 );
xor ( n3432 , n3428 , n3431 );
xor ( n3433 , n3425 , n3432 );
xor ( n3434 , n1910 , n1911 );
xor ( n3435 , n3434 , n2571 );
buf ( n3436 , n3435 );
xor ( n3437 , n1913 , n1914 );
xor ( n3438 , n3437 , n2568 );
buf ( n3439 , n3438 );
xor ( n3440 , n3436 , n3439 );
xor ( n3441 , n1916 , n1917 );
xor ( n3442 , n3441 , n2565 );
buf ( n3443 , n3442 );
xor ( n3444 , n1919 , n1920 );
xor ( n3445 , n3444 , n2562 );
buf ( n3446 , n3445 );
xor ( n3447 , n3443 , n3446 );
xor ( n3448 , n3440 , n3447 );
xor ( n3449 , n3433 , n3448 );
xor ( n3450 , n3418 , n3449 );
xor ( n3451 , n3387 , n3450 );
xor ( n3452 , n3324 , n3451 );
xor ( n3453 , n3197 , n3452 );
xor ( n3454 , n1922 , n1923 );
xor ( n3455 , n3454 , n2559 );
buf ( n3456 , n3455 );
xor ( n3457 , n1925 , n1926 );
xor ( n3458 , n3457 , n2556 );
buf ( n3459 , n3458 );
xor ( n3460 , n3456 , n3459 );
xor ( n3461 , n1928 , n1929 );
xor ( n3462 , n3461 , n2553 );
buf ( n3463 , n3462 );
xor ( n3464 , n1931 , n1932 );
xor ( n3465 , n3464 , n2550 );
buf ( n3466 , n3465 );
xor ( n3467 , n3463 , n3466 );
xor ( n3468 , n3460 , n3467 );
xor ( n3469 , n1934 , n1935 );
xor ( n3470 , n3469 , n2547 );
buf ( n3471 , n3470 );
xor ( n3472 , n1937 , n1938 );
xor ( n3473 , n3472 , n2544 );
buf ( n3474 , n3473 );
xor ( n3475 , n3471 , n3474 );
xor ( n3476 , n1940 , n1941 );
xor ( n3477 , n3476 , n2541 );
buf ( n3478 , n3477 );
xor ( n3479 , n1943 , n1944 );
xor ( n3480 , n3479 , n2538 );
buf ( n3481 , n3480 );
xor ( n3482 , n3478 , n3481 );
xor ( n3483 , n3475 , n3482 );
xor ( n3484 , n3468 , n3483 );
xor ( n3485 , n1946 , n1947 );
xor ( n3486 , n3485 , n2535 );
buf ( n3487 , n3486 );
xor ( n3488 , n1949 , n1950 );
xor ( n3489 , n3488 , n2532 );
buf ( n3490 , n3489 );
xor ( n3491 , n3487 , n3490 );
xor ( n3492 , n1952 , n1953 );
xor ( n3493 , n3492 , n2529 );
buf ( n3494 , n3493 );
xor ( n3495 , n1955 , n1956 );
xor ( n3496 , n3495 , n2526 );
buf ( n3497 , n3496 );
xor ( n3498 , n3494 , n3497 );
xor ( n3499 , n3491 , n3498 );
xor ( n3500 , n1958 , n1959 );
xor ( n3501 , n3500 , n2523 );
buf ( n3502 , n3501 );
xor ( n3503 , n1961 , n1962 );
xor ( n3504 , n3503 , n2520 );
buf ( n3505 , n3504 );
xor ( n3506 , n3502 , n3505 );
xor ( n3507 , n1964 , n1965 );
xor ( n3508 , n3507 , n2517 );
buf ( n3509 , n3508 );
xor ( n3510 , n1967 , n1968 );
xor ( n3511 , n3510 , n2514 );
buf ( n3512 , n3511 );
xor ( n3513 , n3509 , n3512 );
xor ( n3514 , n3506 , n3513 );
xor ( n3515 , n3499 , n3514 );
xor ( n3516 , n3484 , n3515 );
xor ( n3517 , n1970 , n1971 );
xor ( n3518 , n3517 , n2511 );
buf ( n3519 , n3518 );
xor ( n3520 , n1973 , n1974 );
xor ( n3521 , n3520 , n2508 );
buf ( n3522 , n3521 );
xor ( n3523 , n3519 , n3522 );
xor ( n3524 , n1976 , n1977 );
xor ( n3525 , n3524 , n2505 );
buf ( n3526 , n3525 );
xor ( n3527 , n1979 , n1980 );
xor ( n3528 , n3527 , n2502 );
buf ( n3529 , n3528 );
xor ( n3530 , n3526 , n3529 );
xor ( n3531 , n3523 , n3530 );
xor ( n3532 , n1982 , n1983 );
xor ( n3533 , n3532 , n2499 );
buf ( n3534 , n3533 );
xor ( n3535 , n1985 , n1986 );
xor ( n3536 , n3535 , n2496 );
buf ( n3537 , n3536 );
xor ( n3538 , n3534 , n3537 );
xor ( n3539 , n1988 , n1989 );
xor ( n3540 , n3539 , n2493 );
buf ( n3541 , n3540 );
xor ( n3542 , n1991 , n1992 );
xor ( n3543 , n3542 , n2490 );
buf ( n3544 , n3543 );
xor ( n3545 , n3541 , n3544 );
xor ( n3546 , n3538 , n3545 );
xor ( n3547 , n3531 , n3546 );
xor ( n3548 , n1994 , n1995 );
xor ( n3549 , n3548 , n2487 );
buf ( n3550 , n3549 );
xor ( n3551 , n1997 , n1998 );
xor ( n3552 , n3551 , n2484 );
buf ( n3553 , n3552 );
xor ( n3554 , n3550 , n3553 );
xor ( n3555 , n2000 , n2001 );
xor ( n3556 , n3555 , n2481 );
buf ( n3557 , n3556 );
xor ( n3558 , n2003 , n2004 );
xor ( n3559 , n3558 , n2478 );
buf ( n3560 , n3559 );
xor ( n3561 , n3557 , n3560 );
xor ( n3562 , n3554 , n3561 );
xor ( n3563 , n2006 , n2007 );
xor ( n3564 , n3563 , n2475 );
buf ( n3565 , n3564 );
xor ( n3566 , n2009 , n2010 );
xor ( n3567 , n3566 , n2472 );
buf ( n3568 , n3567 );
xor ( n3569 , n3565 , n3568 );
xor ( n3570 , n2012 , n2013 );
xor ( n3571 , n3570 , n2469 );
buf ( n3572 , n3571 );
xor ( n3573 , n2015 , n2016 );
xor ( n3574 , n3573 , n2466 );
buf ( n3575 , n3574 );
xor ( n3576 , n3572 , n3575 );
xor ( n3577 , n3569 , n3576 );
xor ( n3578 , n3562 , n3577 );
xor ( n3579 , n3547 , n3578 );
xor ( n3580 , n3516 , n3579 );
xor ( n3581 , n2018 , n2019 );
xor ( n3582 , n3581 , n2463 );
buf ( n3583 , n3582 );
xor ( n3584 , n2021 , n2022 );
xor ( n3585 , n3584 , n2460 );
buf ( n3586 , n3585 );
xor ( n3587 , n3583 , n3586 );
xor ( n3588 , n2024 , n2025 );
xor ( n3589 , n3588 , n2457 );
buf ( n3590 , n3589 );
xor ( n3591 , n2027 , n2028 );
xor ( n3592 , n3591 , n2454 );
buf ( n3593 , n3592 );
xor ( n3594 , n3590 , n3593 );
xor ( n3595 , n3587 , n3594 );
xor ( n3596 , n2030 , n2031 );
xor ( n3597 , n3596 , n2451 );
buf ( n3598 , n3597 );
xor ( n3599 , n2033 , n2034 );
xor ( n3600 , n3599 , n2448 );
buf ( n3601 , n3600 );
xor ( n3602 , n3598 , n3601 );
xor ( n3603 , n2036 , n2037 );
xor ( n3604 , n3603 , n2445 );
buf ( n3605 , n3604 );
xor ( n3606 , n2039 , n2040 );
xor ( n3607 , n3606 , n2442 );
buf ( n3608 , n3607 );
xor ( n3609 , n3605 , n3608 );
xor ( n3610 , n3602 , n3609 );
xor ( n3611 , n3595 , n3610 );
xor ( n3612 , n2042 , n2043 );
xor ( n3613 , n3612 , n2439 );
buf ( n3614 , n3613 );
xor ( n3615 , n2045 , n2046 );
xor ( n3616 , n3615 , n2436 );
buf ( n3617 , n3616 );
xor ( n3618 , n3614 , n3617 );
xor ( n3619 , n2048 , n2049 );
xor ( n3620 , n3619 , n2433 );
buf ( n3621 , n3620 );
xor ( n3622 , n2051 , n2052 );
xor ( n3623 , n3622 , n2430 );
buf ( n3624 , n3623 );
xor ( n3625 , n3621 , n3624 );
xor ( n3626 , n3618 , n3625 );
xor ( n3627 , n2054 , n2055 );
xor ( n3628 , n3627 , n2427 );
buf ( n3629 , n3628 );
xor ( n3630 , n2057 , n2058 );
xor ( n3631 , n3630 , n2424 );
buf ( n3632 , n3631 );
xor ( n3633 , n3629 , n3632 );
xor ( n3634 , n2060 , n2061 );
xor ( n3635 , n3634 , n2421 );
buf ( n3636 , n3635 );
xor ( n3637 , n2063 , n2064 );
xor ( n3638 , n3637 , n2418 );
buf ( n3639 , n3638 );
xor ( n3640 , n3636 , n3639 );
xor ( n3641 , n3633 , n3640 );
xor ( n3642 , n3626 , n3641 );
xor ( n3643 , n3611 , n3642 );
xor ( n3644 , n2066 , n2067 );
xor ( n3645 , n3644 , n2415 );
buf ( n3646 , n3645 );
xor ( n3647 , n2069 , n2070 );
xor ( n3648 , n3647 , n2412 );
buf ( n3649 , n3648 );
xor ( n3650 , n3646 , n3649 );
xor ( n3651 , n2072 , n2073 );
xor ( n3652 , n3651 , n2409 );
buf ( n3653 , n3652 );
xor ( n3654 , n2075 , n2076 );
xor ( n3655 , n3654 , n2406 );
buf ( n3656 , n3655 );
xor ( n3657 , n3653 , n3656 );
xor ( n3658 , n3650 , n3657 );
xor ( n3659 , n2078 , n2079 );
xor ( n3660 , n3659 , n2403 );
buf ( n3661 , n3660 );
xor ( n3662 , n2081 , n2082 );
xor ( n3663 , n3662 , n2400 );
buf ( n3664 , n3663 );
xor ( n3665 , n3661 , n3664 );
xor ( n3666 , n2084 , n2085 );
xor ( n3667 , n3666 , n2397 );
buf ( n3668 , n3667 );
xor ( n3669 , n2087 , n2088 );
xor ( n3670 , n3669 , n2394 );
buf ( n3671 , n3670 );
xor ( n3672 , n3668 , n3671 );
xor ( n3673 , n3665 , n3672 );
xor ( n3674 , n3658 , n3673 );
xor ( n3675 , n2090 , n2091 );
xor ( n3676 , n3675 , n2391 );
buf ( n3677 , n3676 );
xor ( n3678 , n2093 , n2094 );
xor ( n3679 , n3678 , n2388 );
buf ( n3680 , n3679 );
xor ( n3681 , n3677 , n3680 );
xor ( n3682 , n2096 , n2097 );
xor ( n3683 , n3682 , n2385 );
buf ( n3684 , n3683 );
xor ( n3685 , n2099 , n2100 );
xor ( n3686 , n3685 , n2382 );
buf ( n3687 , n3686 );
xor ( n3688 , n3684 , n3687 );
xor ( n3689 , n3681 , n3688 );
xor ( n3690 , n2102 , n2103 );
xor ( n3691 , n3690 , n2379 );
buf ( n3692 , n3691 );
xor ( n3693 , n2105 , n2106 );
xor ( n3694 , n3693 , n2376 );
buf ( n3695 , n3694 );
xor ( n3696 , n3692 , n3695 );
xor ( n3697 , n2108 , n2109 );
xor ( n3698 , n3697 , n2373 );
buf ( n3699 , n3698 );
xor ( n3700 , n2111 , n2112 );
xor ( n3701 , n3700 , n2370 );
buf ( n3702 , n3701 );
xor ( n3703 , n3699 , n3702 );
xor ( n3704 , n3696 , n3703 );
xor ( n3705 , n3689 , n3704 );
xor ( n3706 , n3674 , n3705 );
xor ( n3707 , n3643 , n3706 );
xor ( n3708 , n3580 , n3707 );
xor ( n3709 , n2114 , n2115 );
xor ( n3710 , n3709 , n2367 );
buf ( n3711 , n3710 );
xor ( n3712 , n2117 , n2118 );
xor ( n3713 , n3712 , n2364 );
buf ( n3714 , n3713 );
xor ( n3715 , n3711 , n3714 );
xor ( n3716 , n2120 , n2121 );
xor ( n3717 , n3716 , n2361 );
buf ( n3718 , n3717 );
xor ( n3719 , n2123 , n2124 );
xor ( n3720 , n3719 , n2358 );
buf ( n3721 , n3720 );
xor ( n3722 , n3718 , n3721 );
xor ( n3723 , n3715 , n3722 );
xor ( n3724 , n2126 , n2127 );
xor ( n3725 , n3724 , n2355 );
buf ( n3726 , n3725 );
xor ( n3727 , n2129 , n2130 );
xor ( n3728 , n3727 , n2352 );
buf ( n3729 , n3728 );
xor ( n3730 , n3726 , n3729 );
xor ( n3731 , n2132 , n2133 );
xor ( n3732 , n3731 , n2349 );
buf ( n3733 , n3732 );
xor ( n3734 , n2135 , n2136 );
xor ( n3735 , n3734 , n2346 );
buf ( n3736 , n3735 );
xor ( n3737 , n3733 , n3736 );
xor ( n3738 , n3730 , n3737 );
xor ( n3739 , n3723 , n3738 );
xor ( n3740 , n2138 , n2139 );
xor ( n3741 , n3740 , n2343 );
buf ( n3742 , n3741 );
xor ( n3743 , n2141 , n2142 );
xor ( n3744 , n3743 , n2340 );
buf ( n3745 , n3744 );
xor ( n3746 , n3742 , n3745 );
xor ( n3747 , n2144 , n2145 );
xor ( n3748 , n3747 , n2337 );
buf ( n3749 , n3748 );
xor ( n3750 , n2147 , n2148 );
xor ( n3751 , n3750 , n2334 );
buf ( n3752 , n3751 );
xor ( n3753 , n3749 , n3752 );
xor ( n3754 , n3746 , n3753 );
xor ( n3755 , n2150 , n2151 );
xor ( n3756 , n3755 , n2331 );
buf ( n3757 , n3756 );
xor ( n3758 , n2153 , n2154 );
xor ( n3759 , n3758 , n2328 );
buf ( n3760 , n3759 );
xor ( n3761 , n3757 , n3760 );
xor ( n3762 , n2156 , n2157 );
xor ( n3763 , n3762 , n2325 );
buf ( n3764 , n3763 );
xor ( n3765 , n2159 , n2160 );
xor ( n3766 , n3765 , n2322 );
buf ( n3767 , n3766 );
xor ( n3768 , n3764 , n3767 );
xor ( n3769 , n3761 , n3768 );
xor ( n3770 , n3754 , n3769 );
xor ( n3771 , n3739 , n3770 );
xor ( n3772 , n2162 , n2163 );
xor ( n3773 , n3772 , n2319 );
buf ( n3774 , n3773 );
xor ( n3775 , n2165 , n2166 );
xor ( n3776 , n3775 , n2316 );
buf ( n3777 , n3776 );
xor ( n3778 , n3774 , n3777 );
xor ( n3779 , n2168 , n2169 );
xor ( n3780 , n3779 , n2313 );
buf ( n3781 , n3780 );
xor ( n3782 , n2171 , n2172 );
xor ( n3783 , n3782 , n2310 );
buf ( n3784 , n3783 );
xor ( n3785 , n3781 , n3784 );
xor ( n3786 , n3778 , n3785 );
xor ( n3787 , n2174 , n2175 );
xor ( n3788 , n3787 , n2307 );
buf ( n3789 , n3788 );
xor ( n3790 , n2177 , n2178 );
xor ( n3791 , n3790 , n2304 );
buf ( n3792 , n3791 );
xor ( n3793 , n3789 , n3792 );
xor ( n3794 , n2180 , n2181 );
xor ( n3795 , n3794 , n2301 );
buf ( n3796 , n3795 );
xor ( n3797 , n2183 , n2184 );
xor ( n3798 , n3797 , n2298 );
buf ( n3799 , n3798 );
xor ( n3800 , n3796 , n3799 );
xor ( n3801 , n3793 , n3800 );
xor ( n3802 , n3786 , n3801 );
xor ( n3803 , n2186 , n2187 );
xor ( n3804 , n3803 , n2295 );
buf ( n3805 , n3804 );
xor ( n3806 , n2189 , n2190 );
xor ( n3807 , n3806 , n2292 );
buf ( n3808 , n3807 );
xor ( n3809 , n3805 , n3808 );
xor ( n3810 , n2192 , n2193 );
xor ( n3811 , n3810 , n2289 );
buf ( n3812 , n3811 );
xor ( n3813 , n2195 , n2196 );
xor ( n3814 , n3813 , n2286 );
buf ( n3815 , n3814 );
xor ( n3816 , n3812 , n3815 );
xor ( n3817 , n3809 , n3816 );
xor ( n3818 , n2198 , n2199 );
xor ( n3819 , n3818 , n2283 );
buf ( n3820 , n3819 );
xor ( n3821 , n2201 , n2202 );
xor ( n3822 , n3821 , n2280 );
buf ( n3823 , n3822 );
xor ( n3824 , n3820 , n3823 );
xor ( n3825 , n2204 , n2205 );
xor ( n3826 , n3825 , n2277 );
buf ( n3827 , n3826 );
xor ( n3828 , n2207 , n2208 );
xor ( n3829 , n3828 , n2274 );
buf ( n3830 , n3829 );
xor ( n3831 , n3827 , n3830 );
xor ( n3832 , n3824 , n3831 );
xor ( n3833 , n3817 , n3832 );
xor ( n3834 , n3802 , n3833 );
xor ( n3835 , n3771 , n3834 );
xor ( n3836 , n2210 , n2211 );
xor ( n3837 , n3836 , n2271 );
buf ( n3838 , n3837 );
xor ( n3839 , n2213 , n2214 );
xor ( n3840 , n3839 , n2268 );
buf ( n3841 , n3840 );
xor ( n3842 , n3838 , n3841 );
xor ( n3843 , n2216 , n2217 );
xor ( n3844 , n3843 , n2265 );
buf ( n3845 , n3844 );
xor ( n3846 , n2219 , n2220 );
xor ( n3847 , n3846 , n2262 );
buf ( n3848 , n3847 );
xor ( n3849 , n3845 , n3848 );
xor ( n3850 , n3842 , n3849 );
xor ( n3851 , n2222 , n2223 );
xor ( n3852 , n3851 , n2259 );
buf ( n3853 , n3852 );
xor ( n3854 , n2225 , n2226 );
xor ( n3855 , n3854 , n2256 );
buf ( n3856 , n3855 );
xor ( n3857 , n3853 , n3856 );
xor ( n3858 , n2228 , n2229 );
xor ( n3859 , n3858 , n2253 );
buf ( n3860 , n3859 );
xor ( n3861 , n2231 , n2232 );
xor ( n3862 , n3861 , n2250 );
buf ( n3863 , n3862 );
xor ( n3864 , n3860 , n3863 );
xor ( n3865 , n3857 , n3864 );
xor ( n3866 , n3850 , n3865 );
not ( n3867 , n2234 );
xor ( n3868 , n3867 , n2247 );
buf ( n3869 , n3868 );
xor ( n3870 , n2236 , n2237 );
xor ( n3871 , n3870 , n2244 );
buf ( n3872 , n3871 );
xor ( n3873 , n3869 , n3872 );
xor ( n3874 , n2239 , n2240 );
not ( n3875 , n3874 );
buf ( n3876 , n3875 );
buf ( n3877 , n1262 );
buf ( n3878 , n1518 );
and ( n3879 , n3877 , n3878 );
buf ( n3880 , n3878 );
buf ( n3881 , n3877 );
or ( n3882 , n3879 , n3880 , n3881 );
buf ( n3883 , n3882 );
buf ( n3884 , n3883 );
xor ( n3885 , n3876 , n3884 );
xor ( n3886 , n3873 , n3885 );
xor ( n3887 , n3877 , n3878 );
not ( n3888 , n3887 );
buf ( n3889 , n3888 );
buf ( n3890 , n1263 );
not ( n3891 , n3890 );
not ( n3892 , n3891 );
buf ( n3893 , n3892 );
xor ( n3894 , n3889 , n3893 );
buf ( n3895 , n1265 );
buf ( n3896 , n1521 );
and ( n3897 , n3895 , n3896 );
buf ( n3898 , n3896 );
buf ( n3899 , n3895 );
or ( n3900 , n3897 , n3898 , n3899 );
buf ( n3901 , n3900 );
buf ( n3902 , n3901 );
xor ( n3903 , n3895 , n3896 );
not ( n3904 , n3903 );
buf ( n3905 , n3904 );
xor ( n3906 , n3902 , n3905 );
xor ( n3907 , n3894 , n3906 );
xor ( n3908 , n3886 , n3907 );
xor ( n3909 , n3866 , n3908 );
buf ( n3910 , n1523 );
not ( n3911 , n3910 );
not ( n3912 , n3911 );
buf ( n3913 , n3912 );
not ( n3914 , n3913 );
buf ( n3915 , n1268 );
not ( n3916 , n3915 );
not ( n3917 , n3916 );
buf ( n3918 , n3917 );
buf ( n3919 , n1270 );
buf ( n3920 , n1526 );
and ( n3921 , n3919 , n3920 );
buf ( n3922 , n3920 );
buf ( n3923 , n3919 );
or ( n3924 , n3921 , n3922 , n3923 );
buf ( n3925 , n3924 );
buf ( n3926 , n3925 );
xor ( n3927 , n3918 , n3926 );
xor ( n3928 , n3914 , n3927 );
xor ( n3929 , n3919 , n3920 );
not ( n3930 , n3929 );
buf ( n3931 , n3930 );
buf ( n3932 , n1528 );
buf ( n3933 , n3932 );
buf ( n3934 , n1273 );
buf ( n3935 , n1529 );
and ( n3936 , n3934 , n3935 );
buf ( n3937 , n1530 );
buf ( n3938 , n3937 );
buf ( n3939 , n1275 );
buf ( n3940 , n1531 );
and ( n3941 , n3939 , n3940 );
buf ( n3942 , n3940 );
buf ( n3943 , n3939 );
or ( n3944 , n3941 , n3942 , n3943 );
and ( n3945 , n3937 , n3944 );
buf ( n3946 , n3944 );
or ( n3947 , n3938 , n3945 , n3946 );
and ( n3948 , n3935 , n3947 );
and ( n3949 , n3934 , n3947 );
or ( n3950 , n3936 , n3948 , n3949 );
and ( n3951 , n3932 , n3950 );
buf ( n3952 , n3950 );
or ( n3953 , n3933 , n3951 , n3952 );
buf ( n3954 , n3953 );
buf ( n3955 , n3954 );
xor ( n3956 , n3931 , n3955 );
not ( n3957 , n3932 );
xor ( n3958 , n3957 , n3950 );
buf ( n3959 , n3958 );
xor ( n3960 , n3934 , n3935 );
xor ( n3961 , n3960 , n3947 );
buf ( n3962 , n3961 );
xor ( n3963 , n3959 , n3962 );
xor ( n3964 , n3956 , n3963 );
xor ( n3965 , n3928 , n3964 );
not ( n3966 , n3937 );
xor ( n3967 , n3966 , n3944 );
buf ( n3968 , n3967 );
xor ( n3969 , n3939 , n3940 );
not ( n3970 , n3969 );
buf ( n3971 , n3970 );
xor ( n3972 , n3968 , n3971 );
buf ( n3973 , n1276 );
not ( n3974 , n3973 );
not ( n3975 , n3974 );
buf ( n3976 , n3975 );
buf ( n3977 , n1277 );
not ( n3978 , n3977 );
not ( n3979 , n3978 );
buf ( n3980 , n3979 );
xor ( n3981 , n3976 , n3980 );
xor ( n3982 , n3972 , n3981 );
buf ( n3983 , n1278 );
not ( n3984 , n3983 );
not ( n3985 , n3984 );
buf ( n3986 , n3985 );
not ( n3987 , n3986 );
not ( n3988 , n3987 );
xor ( n3989 , n3982 , n3988 );
xor ( n3990 , n3965 , n3989 );
xor ( n3991 , n3909 , n3990 );
xor ( n3992 , n3835 , n3991 );
xor ( n3993 , n3708 , n3992 );
xor ( n3994 , n3453 , n3993 );
buf ( n3995 , n3994 );
buf ( n3996 , n3995 );
buf ( n3997 , n1026 );
buf ( n3998 , n1282 );
not ( n3999 , n3998 );
xor ( n4000 , n3997 , n3999 );
buf ( n4001 , n1027 );
buf ( n4002 , n1283 );
not ( n4003 , n4002 );
and ( n4004 , n4001 , n4003 );
buf ( n4005 , n1028 );
buf ( n4006 , n1284 );
not ( n4007 , n4006 );
and ( n4008 , n4005 , n4007 );
buf ( n4009 , n1029 );
buf ( n4010 , n1285 );
not ( n4011 , n4010 );
and ( n4012 , n4009 , n4011 );
buf ( n4013 , n1030 );
buf ( n4014 , n1286 );
not ( n4015 , n4014 );
and ( n4016 , n4013 , n4015 );
buf ( n4017 , n1031 );
buf ( n4018 , n1287 );
not ( n4019 , n4018 );
and ( n4020 , n4017 , n4019 );
buf ( n4021 , n1032 );
buf ( n4022 , n1288 );
not ( n4023 , n4022 );
and ( n4024 , n4021 , n4023 );
buf ( n4025 , n1033 );
buf ( n4026 , n1289 );
not ( n4027 , n4026 );
and ( n4028 , n4025 , n4027 );
buf ( n4029 , n1034 );
buf ( n4030 , n1290 );
not ( n4031 , n4030 );
and ( n4032 , n4029 , n4031 );
buf ( n4033 , n1035 );
buf ( n4034 , n1291 );
not ( n4035 , n4034 );
and ( n4036 , n4033 , n4035 );
buf ( n4037 , n1036 );
buf ( n4038 , n1292 );
not ( n4039 , n4038 );
and ( n4040 , n4037 , n4039 );
buf ( n4041 , n1037 );
buf ( n4042 , n1293 );
not ( n4043 , n4042 );
and ( n4044 , n4041 , n4043 );
buf ( n4045 , n1038 );
buf ( n4046 , n1294 );
not ( n4047 , n4046 );
and ( n4048 , n4045 , n4047 );
buf ( n4049 , n1039 );
buf ( n4050 , n1295 );
not ( n4051 , n4050 );
and ( n4052 , n4049 , n4051 );
buf ( n4053 , n1040 );
buf ( n4054 , n1296 );
not ( n4055 , n4054 );
and ( n4056 , n4053 , n4055 );
buf ( n4057 , n1041 );
buf ( n4058 , n1297 );
not ( n4059 , n4058 );
and ( n4060 , n4057 , n4059 );
buf ( n4061 , n1042 );
buf ( n4062 , n1298 );
not ( n4063 , n4062 );
and ( n4064 , n4061 , n4063 );
buf ( n4065 , n1043 );
buf ( n4066 , n1299 );
not ( n4067 , n4066 );
and ( n4068 , n4065 , n4067 );
buf ( n4069 , n1044 );
buf ( n4070 , n1300 );
not ( n4071 , n4070 );
and ( n4072 , n4069 , n4071 );
buf ( n4073 , n1045 );
buf ( n4074 , n1301 );
not ( n4075 , n4074 );
and ( n4076 , n4073 , n4075 );
buf ( n4077 , n1046 );
buf ( n4078 , n1302 );
not ( n4079 , n4078 );
and ( n4080 , n4077 , n4079 );
buf ( n4081 , n1047 );
buf ( n4082 , n1303 );
not ( n4083 , n4082 );
and ( n4084 , n4081 , n4083 );
buf ( n4085 , n1048 );
buf ( n4086 , n1304 );
not ( n4087 , n4086 );
and ( n4088 , n4085 , n4087 );
buf ( n4089 , n1049 );
buf ( n4090 , n1305 );
not ( n4091 , n4090 );
and ( n4092 , n4089 , n4091 );
buf ( n4093 , n1050 );
buf ( n4094 , n1306 );
not ( n4095 , n4094 );
and ( n4096 , n4093 , n4095 );
buf ( n4097 , n1051 );
buf ( n4098 , n1307 );
not ( n4099 , n4098 );
and ( n4100 , n4097 , n4099 );
buf ( n4101 , n1052 );
buf ( n4102 , n1308 );
not ( n4103 , n4102 );
and ( n4104 , n4101 , n4103 );
buf ( n4105 , n1053 );
buf ( n4106 , n1309 );
not ( n4107 , n4106 );
and ( n4108 , n4105 , n4107 );
buf ( n4109 , n1054 );
buf ( n4110 , n1310 );
not ( n4111 , n4110 );
and ( n4112 , n4109 , n4111 );
buf ( n4113 , n1055 );
buf ( n4114 , n1311 );
not ( n4115 , n4114 );
and ( n4116 , n4113 , n4115 );
buf ( n4117 , n1056 );
buf ( n4118 , n1312 );
not ( n4119 , n4118 );
and ( n4120 , n4117 , n4119 );
buf ( n4121 , n1057 );
buf ( n4122 , n1313 );
not ( n4123 , n4122 );
and ( n4124 , n4121 , n4123 );
buf ( n4125 , n1058 );
buf ( n4126 , n1314 );
not ( n4127 , n4126 );
and ( n4128 , n4125 , n4127 );
buf ( n4129 , n1059 );
buf ( n4130 , n1315 );
not ( n4131 , n4130 );
and ( n4132 , n4129 , n4131 );
buf ( n4133 , n1060 );
buf ( n4134 , n1316 );
not ( n4135 , n4134 );
and ( n4136 , n4133 , n4135 );
buf ( n4137 , n1061 );
buf ( n4138 , n1317 );
not ( n4139 , n4138 );
and ( n4140 , n4137 , n4139 );
buf ( n4141 , n1062 );
buf ( n4142 , n1318 );
not ( n4143 , n4142 );
and ( n4144 , n4141 , n4143 );
buf ( n4145 , n1063 );
buf ( n4146 , n1319 );
not ( n4147 , n4146 );
and ( n4148 , n4145 , n4147 );
buf ( n4149 , n1064 );
buf ( n4150 , n1320 );
not ( n4151 , n4150 );
and ( n4152 , n4149 , n4151 );
buf ( n4153 , n1065 );
buf ( n4154 , n1321 );
not ( n4155 , n4154 );
and ( n4156 , n4153 , n4155 );
buf ( n4157 , n1066 );
buf ( n4158 , n1322 );
not ( n4159 , n4158 );
and ( n4160 , n4157 , n4159 );
buf ( n4161 , n1067 );
buf ( n4162 , n1323 );
not ( n4163 , n4162 );
and ( n4164 , n4161 , n4163 );
buf ( n4165 , n1068 );
buf ( n4166 , n1324 );
not ( n4167 , n4166 );
and ( n4168 , n4165 , n4167 );
buf ( n4169 , n1069 );
buf ( n4170 , n1325 );
not ( n4171 , n4170 );
and ( n4172 , n4169 , n4171 );
buf ( n4173 , n1070 );
buf ( n4174 , n1326 );
not ( n4175 , n4174 );
and ( n4176 , n4173 , n4175 );
buf ( n4177 , n1071 );
buf ( n4178 , n1327 );
not ( n4179 , n4178 );
and ( n4180 , n4177 , n4179 );
buf ( n4181 , n1072 );
buf ( n4182 , n1328 );
not ( n4183 , n4182 );
and ( n4184 , n4181 , n4183 );
buf ( n4185 , n1073 );
buf ( n4186 , n1329 );
not ( n4187 , n4186 );
and ( n4188 , n4185 , n4187 );
buf ( n4189 , n1074 );
buf ( n4190 , n1330 );
not ( n4191 , n4190 );
and ( n4192 , n4189 , n4191 );
buf ( n4193 , n1075 );
buf ( n4194 , n1331 );
not ( n4195 , n4194 );
and ( n4196 , n4193 , n4195 );
buf ( n4197 , n1076 );
buf ( n4198 , n1332 );
not ( n4199 , n4198 );
and ( n4200 , n4197 , n4199 );
buf ( n4201 , n1077 );
buf ( n4202 , n1333 );
not ( n4203 , n4202 );
and ( n4204 , n4201 , n4203 );
buf ( n4205 , n1078 );
buf ( n4206 , n1334 );
not ( n4207 , n4206 );
and ( n4208 , n4205 , n4207 );
buf ( n4209 , n1079 );
buf ( n4210 , n1335 );
not ( n4211 , n4210 );
and ( n4212 , n4209 , n4211 );
buf ( n4213 , n1080 );
buf ( n4214 , n1336 );
not ( n4215 , n4214 );
and ( n4216 , n4213 , n4215 );
buf ( n4217 , n1081 );
buf ( n4218 , n1337 );
not ( n4219 , n4218 );
and ( n4220 , n4217 , n4219 );
buf ( n4221 , n1082 );
buf ( n4222 , n1338 );
not ( n4223 , n4222 );
and ( n4224 , n4221 , n4223 );
buf ( n4225 , n1083 );
buf ( n4226 , n1339 );
not ( n4227 , n4226 );
and ( n4228 , n4225 , n4227 );
buf ( n4229 , n1084 );
buf ( n4230 , n1340 );
not ( n4231 , n4230 );
and ( n4232 , n4229 , n4231 );
buf ( n4233 , n1085 );
buf ( n4234 , n1341 );
not ( n4235 , n4234 );
and ( n4236 , n4233 , n4235 );
buf ( n4237 , n1086 );
buf ( n4238 , n1342 );
not ( n4239 , n4238 );
and ( n4240 , n4237 , n4239 );
buf ( n4241 , n1087 );
buf ( n4242 , n1343 );
not ( n4243 , n4242 );
and ( n4244 , n4241 , n4243 );
buf ( n4245 , n1088 );
buf ( n4246 , n1344 );
not ( n4247 , n4246 );
and ( n4248 , n4245 , n4247 );
buf ( n4249 , n1089 );
buf ( n4250 , n1345 );
not ( n4251 , n4250 );
and ( n4252 , n4249 , n4251 );
buf ( n4253 , n1090 );
buf ( n4254 , n1346 );
not ( n4255 , n4254 );
and ( n4256 , n4253 , n4255 );
buf ( n4257 , n1091 );
buf ( n4258 , n1347 );
not ( n4259 , n4258 );
and ( n4260 , n4257 , n4259 );
buf ( n4261 , n1092 );
buf ( n4262 , n1348 );
not ( n4263 , n4262 );
and ( n4264 , n4261 , n4263 );
buf ( n4265 , n1093 );
buf ( n4266 , n1349 );
not ( n4267 , n4266 );
and ( n4268 , n4265 , n4267 );
buf ( n4269 , n1094 );
buf ( n4270 , n1350 );
not ( n4271 , n4270 );
and ( n4272 , n4269 , n4271 );
buf ( n4273 , n1095 );
buf ( n4274 , n1351 );
not ( n4275 , n4274 );
and ( n4276 , n4273 , n4275 );
buf ( n4277 , n1096 );
buf ( n4278 , n1352 );
not ( n4279 , n4278 );
and ( n4280 , n4277 , n4279 );
buf ( n4281 , n1097 );
buf ( n4282 , n1353 );
not ( n4283 , n4282 );
and ( n4284 , n4281 , n4283 );
buf ( n4285 , n1098 );
buf ( n4286 , n1354 );
not ( n4287 , n4286 );
and ( n4288 , n4285 , n4287 );
buf ( n4289 , n1099 );
buf ( n4290 , n1355 );
not ( n4291 , n4290 );
and ( n4292 , n4289 , n4291 );
buf ( n4293 , n1100 );
buf ( n4294 , n1356 );
not ( n4295 , n4294 );
and ( n4296 , n4293 , n4295 );
buf ( n4297 , n1101 );
buf ( n4298 , n1357 );
not ( n4299 , n4298 );
and ( n4300 , n4297 , n4299 );
buf ( n4301 , n1102 );
buf ( n4302 , n1358 );
not ( n4303 , n4302 );
and ( n4304 , n4301 , n4303 );
buf ( n4305 , n1103 );
buf ( n4306 , n1359 );
not ( n4307 , n4306 );
and ( n4308 , n4305 , n4307 );
buf ( n4309 , n1104 );
buf ( n4310 , n1360 );
not ( n4311 , n4310 );
and ( n4312 , n4309 , n4311 );
buf ( n4313 , n1105 );
buf ( n4314 , n1361 );
not ( n4315 , n4314 );
and ( n4316 , n4313 , n4315 );
buf ( n4317 , n1106 );
buf ( n4318 , n1362 );
not ( n4319 , n4318 );
and ( n4320 , n4317 , n4319 );
buf ( n4321 , n1107 );
buf ( n4322 , n1363 );
not ( n4323 , n4322 );
and ( n4324 , n4321 , n4323 );
buf ( n4325 , n1108 );
buf ( n4326 , n1364 );
not ( n4327 , n4326 );
and ( n4328 , n4325 , n4327 );
buf ( n4329 , n1109 );
buf ( n4330 , n1365 );
not ( n4331 , n4330 );
and ( n4332 , n4329 , n4331 );
buf ( n4333 , n1110 );
buf ( n4334 , n1366 );
not ( n4335 , n4334 );
and ( n4336 , n4333 , n4335 );
buf ( n4337 , n1111 );
buf ( n4338 , n1367 );
not ( n4339 , n4338 );
and ( n4340 , n4337 , n4339 );
buf ( n4341 , n1112 );
buf ( n4342 , n1368 );
not ( n4343 , n4342 );
and ( n4344 , n4341 , n4343 );
buf ( n4345 , n1113 );
buf ( n4346 , n1369 );
not ( n4347 , n4346 );
and ( n4348 , n4345 , n4347 );
buf ( n4349 , n1114 );
buf ( n4350 , n1370 );
not ( n4351 , n4350 );
and ( n4352 , n4349 , n4351 );
buf ( n4353 , n1115 );
buf ( n4354 , n1371 );
not ( n4355 , n4354 );
and ( n4356 , n4353 , n4355 );
buf ( n4357 , n1116 );
buf ( n4358 , n1372 );
not ( n4359 , n4358 );
and ( n4360 , n4357 , n4359 );
buf ( n4361 , n1117 );
buf ( n4362 , n1373 );
not ( n4363 , n4362 );
and ( n4364 , n4361 , n4363 );
buf ( n4365 , n1118 );
buf ( n4366 , n1374 );
not ( n4367 , n4366 );
and ( n4368 , n4365 , n4367 );
buf ( n4369 , n1119 );
buf ( n4370 , n1375 );
not ( n4371 , n4370 );
and ( n4372 , n4369 , n4371 );
buf ( n4373 , n1120 );
buf ( n4374 , n1376 );
not ( n4375 , n4374 );
and ( n4376 , n4373 , n4375 );
buf ( n4377 , n1121 );
buf ( n4378 , n1377 );
not ( n4379 , n4378 );
and ( n4380 , n4377 , n4379 );
buf ( n4381 , n1122 );
buf ( n4382 , n1378 );
not ( n4383 , n4382 );
and ( n4384 , n4381 , n4383 );
buf ( n4385 , n1123 );
buf ( n4386 , n1379 );
not ( n4387 , n4386 );
and ( n4388 , n4385 , n4387 );
buf ( n4389 , n1124 );
buf ( n4390 , n1380 );
not ( n4391 , n4390 );
and ( n4392 , n4389 , n4391 );
buf ( n4393 , n1125 );
buf ( n4394 , n1381 );
not ( n4395 , n4394 );
and ( n4396 , n4393 , n4395 );
buf ( n4397 , n1126 );
buf ( n4398 , n1382 );
not ( n4399 , n4398 );
and ( n4400 , n4397 , n4399 );
buf ( n4401 , n1127 );
buf ( n4402 , n1383 );
not ( n4403 , n4402 );
and ( n4404 , n4401 , n4403 );
buf ( n4405 , n1128 );
buf ( n4406 , n1384 );
not ( n4407 , n4406 );
and ( n4408 , n4405 , n4407 );
buf ( n4409 , n1129 );
buf ( n4410 , n1385 );
not ( n4411 , n4410 );
and ( n4412 , n4409 , n4411 );
buf ( n4413 , n1130 );
buf ( n4414 , n1386 );
not ( n4415 , n4414 );
and ( n4416 , n4413 , n4415 );
buf ( n4417 , n1131 );
buf ( n4418 , n1387 );
not ( n4419 , n4418 );
and ( n4420 , n4417 , n4419 );
buf ( n4421 , n1132 );
buf ( n4422 , n1388 );
not ( n4423 , n4422 );
and ( n4424 , n4421 , n4423 );
buf ( n4425 , n1133 );
buf ( n4426 , n1389 );
not ( n4427 , n4426 );
and ( n4428 , n4425 , n4427 );
buf ( n4429 , n1134 );
buf ( n4430 , n1390 );
not ( n4431 , n4430 );
and ( n4432 , n4429 , n4431 );
buf ( n4433 , n1135 );
buf ( n4434 , n1391 );
not ( n4435 , n4434 );
and ( n4436 , n4433 , n4435 );
buf ( n4437 , n1136 );
buf ( n4438 , n1392 );
not ( n4439 , n4438 );
and ( n4440 , n4437 , n4439 );
buf ( n4441 , n1137 );
buf ( n4442 , n1393 );
not ( n4443 , n4442 );
and ( n4444 , n4441 , n4443 );
buf ( n4445 , n1138 );
buf ( n4446 , n1394 );
not ( n4447 , n4446 );
and ( n4448 , n4445 , n4447 );
buf ( n4449 , n1139 );
buf ( n4450 , n1395 );
not ( n4451 , n4450 );
and ( n4452 , n4449 , n4451 );
buf ( n4453 , n1140 );
buf ( n4454 , n1396 );
not ( n4455 , n4454 );
and ( n4456 , n4453 , n4455 );
buf ( n4457 , n1141 );
buf ( n4458 , n1397 );
not ( n4459 , n4458 );
and ( n4460 , n4457 , n4459 );
buf ( n4461 , n1142 );
buf ( n4462 , n1398 );
not ( n4463 , n4462 );
and ( n4464 , n4461 , n4463 );
buf ( n4465 , n1143 );
buf ( n4466 , n1399 );
not ( n4467 , n4466 );
and ( n4468 , n4465 , n4467 );
buf ( n4469 , n1144 );
buf ( n4470 , n1400 );
not ( n4471 , n4470 );
and ( n4472 , n4469 , n4471 );
buf ( n4473 , n1145 );
buf ( n4474 , n1401 );
not ( n4475 , n4474 );
and ( n4476 , n4473 , n4475 );
buf ( n4477 , n1146 );
buf ( n4478 , n1402 );
not ( n4479 , n4478 );
and ( n4480 , n4477 , n4479 );
buf ( n4481 , n1147 );
buf ( n4482 , n1403 );
not ( n4483 , n4482 );
and ( n4484 , n4481 , n4483 );
buf ( n4485 , n1148 );
buf ( n4486 , n1404 );
not ( n4487 , n4486 );
and ( n4488 , n4485 , n4487 );
buf ( n4489 , n1149 );
buf ( n4490 , n1405 );
not ( n4491 , n4490 );
and ( n4492 , n4489 , n4491 );
buf ( n4493 , n1150 );
buf ( n4494 , n1406 );
not ( n4495 , n4494 );
and ( n4496 , n4493 , n4495 );
buf ( n4497 , n1151 );
buf ( n4498 , n1407 );
not ( n4499 , n4498 );
and ( n4500 , n4497 , n4499 );
buf ( n4501 , n1152 );
buf ( n4502 , n1408 );
not ( n4503 , n4502 );
and ( n4504 , n4501 , n4503 );
buf ( n4505 , n1153 );
buf ( n4506 , n1409 );
not ( n4507 , n4506 );
and ( n4508 , n4505 , n4507 );
buf ( n4509 , n1154 );
buf ( n4510 , n1410 );
not ( n4511 , n4510 );
and ( n4512 , n4509 , n4511 );
buf ( n4513 , n1155 );
buf ( n4514 , n1411 );
not ( n4515 , n4514 );
and ( n4516 , n4513 , n4515 );
buf ( n4517 , n1156 );
buf ( n4518 , n1412 );
not ( n4519 , n4518 );
and ( n4520 , n4517 , n4519 );
buf ( n4521 , n1157 );
buf ( n4522 , n1413 );
not ( n4523 , n4522 );
and ( n4524 , n4521 , n4523 );
buf ( n4525 , n1158 );
buf ( n4526 , n1414 );
not ( n4527 , n4526 );
and ( n4528 , n4525 , n4527 );
buf ( n4529 , n1159 );
buf ( n4530 , n1415 );
not ( n4531 , n4530 );
and ( n4532 , n4529 , n4531 );
buf ( n4533 , n1160 );
buf ( n4534 , n1416 );
not ( n4535 , n4534 );
and ( n4536 , n4533 , n4535 );
buf ( n4537 , n1161 );
buf ( n4538 , n1417 );
not ( n4539 , n4538 );
and ( n4540 , n4537 , n4539 );
buf ( n4541 , n1162 );
buf ( n4542 , n1418 );
not ( n4543 , n4542 );
and ( n4544 , n4541 , n4543 );
buf ( n4545 , n1163 );
buf ( n4546 , n1419 );
not ( n4547 , n4546 );
and ( n4548 , n4545 , n4547 );
buf ( n4549 , n1164 );
buf ( n4550 , n1420 );
not ( n4551 , n4550 );
and ( n4552 , n4549 , n4551 );
buf ( n4553 , n1165 );
buf ( n4554 , n1421 );
not ( n4555 , n4554 );
and ( n4556 , n4553 , n4555 );
buf ( n4557 , n1166 );
buf ( n4558 , n1422 );
not ( n4559 , n4558 );
and ( n4560 , n4557 , n4559 );
buf ( n4561 , n1167 );
buf ( n4562 , n1423 );
not ( n4563 , n4562 );
and ( n4564 , n4561 , n4563 );
buf ( n4565 , n1168 );
buf ( n4566 , n1424 );
not ( n4567 , n4566 );
and ( n4568 , n4565 , n4567 );
buf ( n4569 , n1169 );
buf ( n4570 , n1425 );
not ( n4571 , n4570 );
and ( n4572 , n4569 , n4571 );
buf ( n4573 , n1170 );
buf ( n4574 , n1426 );
not ( n4575 , n4574 );
and ( n4576 , n4573 , n4575 );
buf ( n4577 , n1171 );
buf ( n4578 , n1427 );
not ( n4579 , n4578 );
and ( n4580 , n4577 , n4579 );
buf ( n4581 , n1172 );
buf ( n4582 , n1428 );
not ( n4583 , n4582 );
and ( n4584 , n4581 , n4583 );
buf ( n4585 , n1173 );
buf ( n4586 , n1429 );
not ( n4587 , n4586 );
and ( n4588 , n4585 , n4587 );
buf ( n4589 , n1174 );
buf ( n4590 , n1430 );
not ( n4591 , n4590 );
and ( n4592 , n4589 , n4591 );
buf ( n4593 , n1175 );
buf ( n4594 , n1431 );
not ( n4595 , n4594 );
and ( n4596 , n4593 , n4595 );
buf ( n4597 , n1176 );
buf ( n4598 , n1432 );
not ( n4599 , n4598 );
and ( n4600 , n4597 , n4599 );
buf ( n4601 , n1177 );
buf ( n4602 , n1433 );
not ( n4603 , n4602 );
and ( n4604 , n4601 , n4603 );
buf ( n4605 , n1178 );
buf ( n4606 , n1434 );
not ( n4607 , n4606 );
and ( n4608 , n4605 , n4607 );
buf ( n4609 , n1179 );
buf ( n4610 , n1435 );
not ( n4611 , n4610 );
and ( n4612 , n4609 , n4611 );
buf ( n4613 , n1180 );
buf ( n4614 , n1436 );
not ( n4615 , n4614 );
and ( n4616 , n4613 , n4615 );
buf ( n4617 , n1181 );
buf ( n4618 , n1437 );
not ( n4619 , n4618 );
and ( n4620 , n4617 , n4619 );
buf ( n4621 , n1182 );
buf ( n4622 , n1438 );
not ( n4623 , n4622 );
and ( n4624 , n4621 , n4623 );
buf ( n4625 , n1183 );
buf ( n4626 , n1439 );
not ( n4627 , n4626 );
and ( n4628 , n4625 , n4627 );
buf ( n4629 , n1184 );
buf ( n4630 , n1440 );
not ( n4631 , n4630 );
and ( n4632 , n4629 , n4631 );
buf ( n4633 , n1185 );
buf ( n4634 , n1441 );
not ( n4635 , n4634 );
and ( n4636 , n4633 , n4635 );
buf ( n4637 , n1186 );
buf ( n4638 , n1442 );
not ( n4639 , n4638 );
and ( n4640 , n4637 , n4639 );
buf ( n4641 , n1187 );
buf ( n4642 , n1443 );
not ( n4643 , n4642 );
and ( n4644 , n4641 , n4643 );
buf ( n4645 , n1188 );
buf ( n4646 , n1444 );
not ( n4647 , n4646 );
and ( n4648 , n4645 , n4647 );
buf ( n4649 , n1189 );
buf ( n4650 , n1445 );
not ( n4651 , n4650 );
and ( n4652 , n4649 , n4651 );
buf ( n4653 , n1190 );
buf ( n4654 , n1446 );
not ( n4655 , n4654 );
and ( n4656 , n4653 , n4655 );
buf ( n4657 , n1191 );
buf ( n4658 , n1447 );
not ( n4659 , n4658 );
and ( n4660 , n4657 , n4659 );
buf ( n4661 , n1192 );
buf ( n4662 , n1448 );
not ( n4663 , n4662 );
and ( n4664 , n4661 , n4663 );
buf ( n4665 , n1193 );
buf ( n4666 , n1449 );
not ( n4667 , n4666 );
and ( n4668 , n4665 , n4667 );
buf ( n4669 , n1194 );
buf ( n4670 , n1450 );
not ( n4671 , n4670 );
and ( n4672 , n4669 , n4671 );
buf ( n4673 , n1195 );
buf ( n4674 , n1451 );
not ( n4675 , n4674 );
and ( n4676 , n4673 , n4675 );
buf ( n4677 , n1196 );
buf ( n4678 , n1452 );
not ( n4679 , n4678 );
and ( n4680 , n4677 , n4679 );
buf ( n4681 , n1197 );
buf ( n4682 , n1453 );
not ( n4683 , n4682 );
and ( n4684 , n4681 , n4683 );
buf ( n4685 , n1198 );
buf ( n4686 , n1454 );
not ( n4687 , n4686 );
and ( n4688 , n4685 , n4687 );
buf ( n4689 , n1199 );
buf ( n4690 , n1455 );
not ( n4691 , n4690 );
and ( n4692 , n4689 , n4691 );
buf ( n4693 , n1200 );
buf ( n4694 , n1456 );
not ( n4695 , n4694 );
and ( n4696 , n4693 , n4695 );
buf ( n4697 , n1201 );
buf ( n4698 , n1457 );
not ( n4699 , n4698 );
and ( n4700 , n4697 , n4699 );
buf ( n4701 , n1202 );
buf ( n4702 , n1458 );
not ( n4703 , n4702 );
and ( n4704 , n4701 , n4703 );
buf ( n4705 , n1203 );
buf ( n4706 , n1459 );
not ( n4707 , n4706 );
and ( n4708 , n4705 , n4707 );
buf ( n4709 , n1204 );
buf ( n4710 , n1460 );
not ( n4711 , n4710 );
and ( n4712 , n4709 , n4711 );
buf ( n4713 , n1205 );
buf ( n4714 , n1461 );
not ( n4715 , n4714 );
and ( n4716 , n4713 , n4715 );
buf ( n4717 , n1206 );
buf ( n4718 , n1462 );
not ( n4719 , n4718 );
and ( n4720 , n4717 , n4719 );
buf ( n4721 , n1207 );
buf ( n4722 , n1463 );
not ( n4723 , n4722 );
and ( n4724 , n4721 , n4723 );
buf ( n4725 , n1208 );
buf ( n4726 , n1464 );
not ( n4727 , n4726 );
and ( n4728 , n4725 , n4727 );
buf ( n4729 , n1209 );
buf ( n4730 , n1465 );
not ( n4731 , n4730 );
and ( n4732 , n4729 , n4731 );
buf ( n4733 , n1210 );
buf ( n4734 , n1466 );
not ( n4735 , n4734 );
and ( n4736 , n4733 , n4735 );
buf ( n4737 , n1211 );
buf ( n4738 , n1467 );
not ( n4739 , n4738 );
and ( n4740 , n4737 , n4739 );
buf ( n4741 , n1212 );
buf ( n4742 , n1468 );
not ( n4743 , n4742 );
and ( n4744 , n4741 , n4743 );
buf ( n4745 , n1213 );
buf ( n4746 , n1469 );
not ( n4747 , n4746 );
and ( n4748 , n4745 , n4747 );
buf ( n4749 , n1214 );
buf ( n4750 , n1470 );
not ( n4751 , n4750 );
and ( n4752 , n4749 , n4751 );
buf ( n4753 , n1215 );
buf ( n4754 , n1471 );
not ( n4755 , n4754 );
and ( n4756 , n4753 , n4755 );
buf ( n4757 , n1216 );
buf ( n4758 , n1472 );
not ( n4759 , n4758 );
and ( n4760 , n4757 , n4759 );
buf ( n4761 , n1217 );
buf ( n4762 , n1473 );
not ( n4763 , n4762 );
and ( n4764 , n4761 , n4763 );
buf ( n4765 , n1218 );
buf ( n4766 , n1474 );
not ( n4767 , n4766 );
and ( n4768 , n4765 , n4767 );
buf ( n4769 , n1219 );
buf ( n4770 , n1475 );
not ( n4771 , n4770 );
and ( n4772 , n4769 , n4771 );
buf ( n4773 , n1220 );
buf ( n4774 , n1476 );
not ( n4775 , n4774 );
and ( n4776 , n4773 , n4775 );
buf ( n4777 , n1221 );
buf ( n4778 , n1477 );
not ( n4779 , n4778 );
and ( n4780 , n4777 , n4779 );
buf ( n4781 , n1222 );
buf ( n4782 , n1478 );
not ( n4783 , n4782 );
and ( n4784 , n4781 , n4783 );
buf ( n4785 , n1223 );
buf ( n4786 , n1479 );
not ( n4787 , n4786 );
and ( n4788 , n4785 , n4787 );
buf ( n4789 , n1224 );
buf ( n4790 , n1480 );
not ( n4791 , n4790 );
and ( n4792 , n4789 , n4791 );
buf ( n4793 , n1225 );
buf ( n4794 , n1481 );
not ( n4795 , n4794 );
and ( n4796 , n4793 , n4795 );
buf ( n4797 , n1226 );
buf ( n4798 , n1482 );
not ( n4799 , n4798 );
and ( n4800 , n4797 , n4799 );
buf ( n4801 , n1227 );
buf ( n4802 , n1483 );
not ( n4803 , n4802 );
and ( n4804 , n4801 , n4803 );
buf ( n4805 , n1228 );
buf ( n4806 , n1484 );
not ( n4807 , n4806 );
and ( n4808 , n4805 , n4807 );
buf ( n4809 , n1229 );
buf ( n4810 , n1485 );
not ( n4811 , n4810 );
and ( n4812 , n4809 , n4811 );
buf ( n4813 , n1230 );
buf ( n4814 , n1486 );
not ( n4815 , n4814 );
and ( n4816 , n4813 , n4815 );
buf ( n4817 , n1231 );
buf ( n4818 , n1487 );
not ( n4819 , n4818 );
and ( n4820 , n4817 , n4819 );
buf ( n4821 , n1232 );
buf ( n4822 , n1488 );
not ( n4823 , n4822 );
and ( n4824 , n4821 , n4823 );
buf ( n4825 , n1233 );
buf ( n4826 , n1489 );
not ( n4827 , n4826 );
and ( n4828 , n4825 , n4827 );
buf ( n4829 , n1234 );
buf ( n4830 , n1490 );
not ( n4831 , n4830 );
and ( n4832 , n4829 , n4831 );
buf ( n4833 , n1235 );
buf ( n4834 , n1491 );
not ( n4835 , n4834 );
and ( n4836 , n4833 , n4835 );
buf ( n4837 , n1236 );
buf ( n4838 , n1492 );
not ( n4839 , n4838 );
and ( n4840 , n4837 , n4839 );
buf ( n4841 , n1237 );
buf ( n4842 , n1493 );
not ( n4843 , n4842 );
and ( n4844 , n4841 , n4843 );
buf ( n4845 , n1238 );
buf ( n4846 , n1494 );
not ( n4847 , n4846 );
and ( n4848 , n4845 , n4847 );
buf ( n4849 , n1239 );
buf ( n4850 , n1495 );
not ( n4851 , n4850 );
and ( n4852 , n4849 , n4851 );
buf ( n4853 , n1240 );
buf ( n4854 , n1496 );
not ( n4855 , n4854 );
and ( n4856 , n4853 , n4855 );
buf ( n4857 , n1241 );
buf ( n4858 , n1497 );
not ( n4859 , n4858 );
and ( n4860 , n4857 , n4859 );
buf ( n4861 , n1242 );
buf ( n4862 , n1498 );
not ( n4863 , n4862 );
and ( n4864 , n4861 , n4863 );
buf ( n4865 , n1243 );
buf ( n4866 , n1499 );
not ( n4867 , n4866 );
and ( n4868 , n4865 , n4867 );
buf ( n4869 , n1244 );
buf ( n4870 , n1500 );
not ( n4871 , n4870 );
and ( n4872 , n4869 , n4871 );
buf ( n4873 , n1245 );
buf ( n4874 , n1501 );
not ( n4875 , n4874 );
and ( n4876 , n4873 , n4875 );
buf ( n4877 , n1246 );
buf ( n4878 , n1502 );
not ( n4879 , n4878 );
and ( n4880 , n4877 , n4879 );
buf ( n4881 , n1247 );
buf ( n4882 , n1503 );
not ( n4883 , n4882 );
and ( n4884 , n4881 , n4883 );
buf ( n4885 , n1248 );
buf ( n4886 , n1504 );
not ( n4887 , n4886 );
and ( n4888 , n4885 , n4887 );
buf ( n4889 , n1249 );
buf ( n4890 , n1505 );
not ( n4891 , n4890 );
and ( n4892 , n4889 , n4891 );
buf ( n4893 , n1250 );
buf ( n4894 , n1506 );
not ( n4895 , n4894 );
and ( n4896 , n4893 , n4895 );
buf ( n4897 , n1251 );
buf ( n4898 , n1507 );
not ( n4899 , n4898 );
and ( n4900 , n4897 , n4899 );
buf ( n4901 , n1252 );
buf ( n4902 , n1508 );
not ( n4903 , n4902 );
and ( n4904 , n4901 , n4903 );
buf ( n4905 , n1253 );
buf ( n4906 , n1509 );
not ( n4907 , n4906 );
and ( n4908 , n4905 , n4907 );
buf ( n4909 , n1254 );
buf ( n4910 , n1510 );
not ( n4911 , n4910 );
and ( n4912 , n4909 , n4911 );
buf ( n4913 , n1255 );
buf ( n4914 , n1511 );
not ( n4915 , n4914 );
and ( n4916 , n4913 , n4915 );
buf ( n4917 , n1256 );
buf ( n4918 , n1512 );
not ( n4919 , n4918 );
and ( n4920 , n4917 , n4919 );
buf ( n4921 , n1257 );
buf ( n4922 , n1513 );
not ( n4923 , n4922 );
and ( n4924 , n4921 , n4923 );
buf ( n4925 , n1258 );
buf ( n4926 , n1514 );
not ( n4927 , n4926 );
and ( n4928 , n4925 , n4927 );
buf ( n4929 , n1259 );
buf ( n4930 , n1515 );
not ( n4931 , n4930 );
and ( n4932 , n4929 , n4931 );
buf ( n4933 , n1260 );
buf ( n4934 , n1516 );
not ( n4935 , n4934 );
and ( n4936 , n4933 , n4935 );
buf ( n4937 , n1261 );
buf ( n4938 , n1517 );
not ( n4939 , n4938 );
and ( n4940 , n4937 , n4939 );
buf ( n4941 , n1262 );
buf ( n4942 , n1518 );
not ( n4943 , n4942 );
and ( n4944 , n4941 , n4943 );
buf ( n4945 , n1263 );
buf ( n4946 , n1519 );
not ( n4947 , n4946 );
and ( n4948 , n4945 , n4947 );
buf ( n4949 , n1264 );
buf ( n4950 , n1520 );
not ( n4951 , n4950 );
and ( n4952 , n4949 , n4951 );
buf ( n4953 , n1265 );
buf ( n4954 , n1521 );
not ( n4955 , n4954 );
and ( n4956 , n4953 , n4955 );
buf ( n4957 , n1266 );
buf ( n4958 , n1522 );
not ( n4959 , n4958 );
and ( n4960 , n4957 , n4959 );
buf ( n4961 , n1267 );
buf ( n4962 , n1523 );
not ( n4963 , n4962 );
and ( n4964 , n4961 , n4963 );
buf ( n4965 , n1268 );
buf ( n4966 , n1524 );
not ( n4967 , n4966 );
and ( n4968 , n4965 , n4967 );
buf ( n4969 , n1269 );
buf ( n4970 , n1525 );
not ( n4971 , n4970 );
and ( n4972 , n4969 , n4971 );
buf ( n4973 , n1270 );
buf ( n4974 , n1526 );
not ( n4975 , n4974 );
and ( n4976 , n4973 , n4975 );
buf ( n4977 , n1271 );
buf ( n4978 , n1527 );
not ( n4979 , n4978 );
and ( n4980 , n4977 , n4979 );
buf ( n4981 , n1272 );
buf ( n4982 , n1528 );
not ( n4983 , n4982 );
and ( n4984 , n4981 , n4983 );
buf ( n4985 , n1273 );
buf ( n4986 , n1529 );
not ( n4987 , n4986 );
and ( n4988 , n4985 , n4987 );
buf ( n4989 , n1274 );
buf ( n4990 , n1530 );
not ( n4991 , n4990 );
and ( n4992 , n4989 , n4991 );
buf ( n4993 , n1275 );
buf ( n4994 , n1531 );
not ( n4995 , n4994 );
and ( n4996 , n4993 , n4995 );
buf ( n4997 , n1276 );
buf ( n4998 , n1532 );
not ( n4999 , n4998 );
and ( n5000 , n4997 , n4999 );
buf ( n5001 , n1277 );
buf ( n5002 , n1533 );
not ( n5003 , n5002 );
and ( n5004 , n5001 , n5003 );
buf ( n5005 , n1278 );
buf ( n5006 , n1534 );
not ( n5007 , n5006 );
and ( n5008 , n5005 , n5007 );
buf ( n5009 , n1279 );
buf ( n5010 , n1535 );
not ( n5011 , n5010 );
and ( n5012 , n5009 , n5011 );
buf ( n5013 , n1280 );
buf ( n5014 , n1536 );
not ( n5015 , n5014 );
and ( n5016 , n5013 , n5015 );
buf ( n5017 , n1281 );
buf ( n5018 , n1537 );
not ( n5019 , n5018 );
or ( n5020 , n5017 , n5019 );
and ( n5021 , n5015 , n5020 );
and ( n5022 , n5013 , n5020 );
or ( n5023 , n5016 , n5021 , n5022 );
and ( n5024 , n5011 , n5023 );
and ( n5025 , n5009 , n5023 );
or ( n5026 , n5012 , n5024 , n5025 );
and ( n5027 , n5007 , n5026 );
and ( n5028 , n5005 , n5026 );
or ( n5029 , n5008 , n5027 , n5028 );
and ( n5030 , n5003 , n5029 );
and ( n5031 , n5001 , n5029 );
or ( n5032 , n5004 , n5030 , n5031 );
and ( n5033 , n4999 , n5032 );
and ( n5034 , n4997 , n5032 );
or ( n5035 , n5000 , n5033 , n5034 );
and ( n5036 , n4995 , n5035 );
and ( n5037 , n4993 , n5035 );
or ( n5038 , n4996 , n5036 , n5037 );
and ( n5039 , n4991 , n5038 );
and ( n5040 , n4989 , n5038 );
or ( n5041 , n4992 , n5039 , n5040 );
and ( n5042 , n4987 , n5041 );
and ( n5043 , n4985 , n5041 );
or ( n5044 , n4988 , n5042 , n5043 );
and ( n5045 , n4983 , n5044 );
and ( n5046 , n4981 , n5044 );
or ( n5047 , n4984 , n5045 , n5046 );
and ( n5048 , n4979 , n5047 );
and ( n5049 , n4977 , n5047 );
or ( n5050 , n4980 , n5048 , n5049 );
and ( n5051 , n4975 , n5050 );
and ( n5052 , n4973 , n5050 );
or ( n5053 , n4976 , n5051 , n5052 );
and ( n5054 , n4971 , n5053 );
and ( n5055 , n4969 , n5053 );
or ( n5056 , n4972 , n5054 , n5055 );
and ( n5057 , n4967 , n5056 );
and ( n5058 , n4965 , n5056 );
or ( n5059 , n4968 , n5057 , n5058 );
and ( n5060 , n4963 , n5059 );
and ( n5061 , n4961 , n5059 );
or ( n5062 , n4964 , n5060 , n5061 );
and ( n5063 , n4959 , n5062 );
and ( n5064 , n4957 , n5062 );
or ( n5065 , n4960 , n5063 , n5064 );
and ( n5066 , n4955 , n5065 );
and ( n5067 , n4953 , n5065 );
or ( n5068 , n4956 , n5066 , n5067 );
and ( n5069 , n4951 , n5068 );
and ( n5070 , n4949 , n5068 );
or ( n5071 , n4952 , n5069 , n5070 );
and ( n5072 , n4947 , n5071 );
and ( n5073 , n4945 , n5071 );
or ( n5074 , n4948 , n5072 , n5073 );
and ( n5075 , n4943 , n5074 );
and ( n5076 , n4941 , n5074 );
or ( n5077 , n4944 , n5075 , n5076 );
and ( n5078 , n4939 , n5077 );
and ( n5079 , n4937 , n5077 );
or ( n5080 , n4940 , n5078 , n5079 );
and ( n5081 , n4935 , n5080 );
and ( n5082 , n4933 , n5080 );
or ( n5083 , n4936 , n5081 , n5082 );
and ( n5084 , n4931 , n5083 );
and ( n5085 , n4929 , n5083 );
or ( n5086 , n4932 , n5084 , n5085 );
and ( n5087 , n4927 , n5086 );
and ( n5088 , n4925 , n5086 );
or ( n5089 , n4928 , n5087 , n5088 );
and ( n5090 , n4923 , n5089 );
and ( n5091 , n4921 , n5089 );
or ( n5092 , n4924 , n5090 , n5091 );
and ( n5093 , n4919 , n5092 );
and ( n5094 , n4917 , n5092 );
or ( n5095 , n4920 , n5093 , n5094 );
and ( n5096 , n4915 , n5095 );
and ( n5097 , n4913 , n5095 );
or ( n5098 , n4916 , n5096 , n5097 );
and ( n5099 , n4911 , n5098 );
and ( n5100 , n4909 , n5098 );
or ( n5101 , n4912 , n5099 , n5100 );
and ( n5102 , n4907 , n5101 );
and ( n5103 , n4905 , n5101 );
or ( n5104 , n4908 , n5102 , n5103 );
and ( n5105 , n4903 , n5104 );
and ( n5106 , n4901 , n5104 );
or ( n5107 , n4904 , n5105 , n5106 );
and ( n5108 , n4899 , n5107 );
and ( n5109 , n4897 , n5107 );
or ( n5110 , n4900 , n5108 , n5109 );
and ( n5111 , n4895 , n5110 );
and ( n5112 , n4893 , n5110 );
or ( n5113 , n4896 , n5111 , n5112 );
and ( n5114 , n4891 , n5113 );
and ( n5115 , n4889 , n5113 );
or ( n5116 , n4892 , n5114 , n5115 );
and ( n5117 , n4887 , n5116 );
and ( n5118 , n4885 , n5116 );
or ( n5119 , n4888 , n5117 , n5118 );
and ( n5120 , n4883 , n5119 );
and ( n5121 , n4881 , n5119 );
or ( n5122 , n4884 , n5120 , n5121 );
and ( n5123 , n4879 , n5122 );
and ( n5124 , n4877 , n5122 );
or ( n5125 , n4880 , n5123 , n5124 );
and ( n5126 , n4875 , n5125 );
and ( n5127 , n4873 , n5125 );
or ( n5128 , n4876 , n5126 , n5127 );
and ( n5129 , n4871 , n5128 );
and ( n5130 , n4869 , n5128 );
or ( n5131 , n4872 , n5129 , n5130 );
and ( n5132 , n4867 , n5131 );
and ( n5133 , n4865 , n5131 );
or ( n5134 , n4868 , n5132 , n5133 );
and ( n5135 , n4863 , n5134 );
and ( n5136 , n4861 , n5134 );
or ( n5137 , n4864 , n5135 , n5136 );
and ( n5138 , n4859 , n5137 );
and ( n5139 , n4857 , n5137 );
or ( n5140 , n4860 , n5138 , n5139 );
and ( n5141 , n4855 , n5140 );
and ( n5142 , n4853 , n5140 );
or ( n5143 , n4856 , n5141 , n5142 );
and ( n5144 , n4851 , n5143 );
and ( n5145 , n4849 , n5143 );
or ( n5146 , n4852 , n5144 , n5145 );
and ( n5147 , n4847 , n5146 );
and ( n5148 , n4845 , n5146 );
or ( n5149 , n4848 , n5147 , n5148 );
and ( n5150 , n4843 , n5149 );
and ( n5151 , n4841 , n5149 );
or ( n5152 , n4844 , n5150 , n5151 );
and ( n5153 , n4839 , n5152 );
and ( n5154 , n4837 , n5152 );
or ( n5155 , n4840 , n5153 , n5154 );
and ( n5156 , n4835 , n5155 );
and ( n5157 , n4833 , n5155 );
or ( n5158 , n4836 , n5156 , n5157 );
and ( n5159 , n4831 , n5158 );
and ( n5160 , n4829 , n5158 );
or ( n5161 , n4832 , n5159 , n5160 );
and ( n5162 , n4827 , n5161 );
and ( n5163 , n4825 , n5161 );
or ( n5164 , n4828 , n5162 , n5163 );
and ( n5165 , n4823 , n5164 );
and ( n5166 , n4821 , n5164 );
or ( n5167 , n4824 , n5165 , n5166 );
and ( n5168 , n4819 , n5167 );
and ( n5169 , n4817 , n5167 );
or ( n5170 , n4820 , n5168 , n5169 );
and ( n5171 , n4815 , n5170 );
and ( n5172 , n4813 , n5170 );
or ( n5173 , n4816 , n5171 , n5172 );
and ( n5174 , n4811 , n5173 );
and ( n5175 , n4809 , n5173 );
or ( n5176 , n4812 , n5174 , n5175 );
and ( n5177 , n4807 , n5176 );
and ( n5178 , n4805 , n5176 );
or ( n5179 , n4808 , n5177 , n5178 );
and ( n5180 , n4803 , n5179 );
and ( n5181 , n4801 , n5179 );
or ( n5182 , n4804 , n5180 , n5181 );
and ( n5183 , n4799 , n5182 );
and ( n5184 , n4797 , n5182 );
or ( n5185 , n4800 , n5183 , n5184 );
and ( n5186 , n4795 , n5185 );
and ( n5187 , n4793 , n5185 );
or ( n5188 , n4796 , n5186 , n5187 );
and ( n5189 , n4791 , n5188 );
and ( n5190 , n4789 , n5188 );
or ( n5191 , n4792 , n5189 , n5190 );
and ( n5192 , n4787 , n5191 );
and ( n5193 , n4785 , n5191 );
or ( n5194 , n4788 , n5192 , n5193 );
and ( n5195 , n4783 , n5194 );
and ( n5196 , n4781 , n5194 );
or ( n5197 , n4784 , n5195 , n5196 );
and ( n5198 , n4779 , n5197 );
and ( n5199 , n4777 , n5197 );
or ( n5200 , n4780 , n5198 , n5199 );
and ( n5201 , n4775 , n5200 );
and ( n5202 , n4773 , n5200 );
or ( n5203 , n4776 , n5201 , n5202 );
and ( n5204 , n4771 , n5203 );
and ( n5205 , n4769 , n5203 );
or ( n5206 , n4772 , n5204 , n5205 );
and ( n5207 , n4767 , n5206 );
and ( n5208 , n4765 , n5206 );
or ( n5209 , n4768 , n5207 , n5208 );
and ( n5210 , n4763 , n5209 );
and ( n5211 , n4761 , n5209 );
or ( n5212 , n4764 , n5210 , n5211 );
and ( n5213 , n4759 , n5212 );
and ( n5214 , n4757 , n5212 );
or ( n5215 , n4760 , n5213 , n5214 );
and ( n5216 , n4755 , n5215 );
and ( n5217 , n4753 , n5215 );
or ( n5218 , n4756 , n5216 , n5217 );
and ( n5219 , n4751 , n5218 );
and ( n5220 , n4749 , n5218 );
or ( n5221 , n4752 , n5219 , n5220 );
and ( n5222 , n4747 , n5221 );
and ( n5223 , n4745 , n5221 );
or ( n5224 , n4748 , n5222 , n5223 );
and ( n5225 , n4743 , n5224 );
and ( n5226 , n4741 , n5224 );
or ( n5227 , n4744 , n5225 , n5226 );
and ( n5228 , n4739 , n5227 );
and ( n5229 , n4737 , n5227 );
or ( n5230 , n4740 , n5228 , n5229 );
and ( n5231 , n4735 , n5230 );
and ( n5232 , n4733 , n5230 );
or ( n5233 , n4736 , n5231 , n5232 );
and ( n5234 , n4731 , n5233 );
and ( n5235 , n4729 , n5233 );
or ( n5236 , n4732 , n5234 , n5235 );
and ( n5237 , n4727 , n5236 );
and ( n5238 , n4725 , n5236 );
or ( n5239 , n4728 , n5237 , n5238 );
and ( n5240 , n4723 , n5239 );
and ( n5241 , n4721 , n5239 );
or ( n5242 , n4724 , n5240 , n5241 );
and ( n5243 , n4719 , n5242 );
and ( n5244 , n4717 , n5242 );
or ( n5245 , n4720 , n5243 , n5244 );
and ( n5246 , n4715 , n5245 );
and ( n5247 , n4713 , n5245 );
or ( n5248 , n4716 , n5246 , n5247 );
and ( n5249 , n4711 , n5248 );
and ( n5250 , n4709 , n5248 );
or ( n5251 , n4712 , n5249 , n5250 );
and ( n5252 , n4707 , n5251 );
and ( n5253 , n4705 , n5251 );
or ( n5254 , n4708 , n5252 , n5253 );
and ( n5255 , n4703 , n5254 );
and ( n5256 , n4701 , n5254 );
or ( n5257 , n4704 , n5255 , n5256 );
and ( n5258 , n4699 , n5257 );
and ( n5259 , n4697 , n5257 );
or ( n5260 , n4700 , n5258 , n5259 );
and ( n5261 , n4695 , n5260 );
and ( n5262 , n4693 , n5260 );
or ( n5263 , n4696 , n5261 , n5262 );
and ( n5264 , n4691 , n5263 );
and ( n5265 , n4689 , n5263 );
or ( n5266 , n4692 , n5264 , n5265 );
and ( n5267 , n4687 , n5266 );
and ( n5268 , n4685 , n5266 );
or ( n5269 , n4688 , n5267 , n5268 );
and ( n5270 , n4683 , n5269 );
and ( n5271 , n4681 , n5269 );
or ( n5272 , n4684 , n5270 , n5271 );
and ( n5273 , n4679 , n5272 );
and ( n5274 , n4677 , n5272 );
or ( n5275 , n4680 , n5273 , n5274 );
and ( n5276 , n4675 , n5275 );
and ( n5277 , n4673 , n5275 );
or ( n5278 , n4676 , n5276 , n5277 );
and ( n5279 , n4671 , n5278 );
and ( n5280 , n4669 , n5278 );
or ( n5281 , n4672 , n5279 , n5280 );
and ( n5282 , n4667 , n5281 );
and ( n5283 , n4665 , n5281 );
or ( n5284 , n4668 , n5282 , n5283 );
and ( n5285 , n4663 , n5284 );
and ( n5286 , n4661 , n5284 );
or ( n5287 , n4664 , n5285 , n5286 );
and ( n5288 , n4659 , n5287 );
and ( n5289 , n4657 , n5287 );
or ( n5290 , n4660 , n5288 , n5289 );
and ( n5291 , n4655 , n5290 );
and ( n5292 , n4653 , n5290 );
or ( n5293 , n4656 , n5291 , n5292 );
and ( n5294 , n4651 , n5293 );
and ( n5295 , n4649 , n5293 );
or ( n5296 , n4652 , n5294 , n5295 );
and ( n5297 , n4647 , n5296 );
and ( n5298 , n4645 , n5296 );
or ( n5299 , n4648 , n5297 , n5298 );
and ( n5300 , n4643 , n5299 );
and ( n5301 , n4641 , n5299 );
or ( n5302 , n4644 , n5300 , n5301 );
and ( n5303 , n4639 , n5302 );
and ( n5304 , n4637 , n5302 );
or ( n5305 , n4640 , n5303 , n5304 );
and ( n5306 , n4635 , n5305 );
and ( n5307 , n4633 , n5305 );
or ( n5308 , n4636 , n5306 , n5307 );
and ( n5309 , n4631 , n5308 );
and ( n5310 , n4629 , n5308 );
or ( n5311 , n4632 , n5309 , n5310 );
and ( n5312 , n4627 , n5311 );
and ( n5313 , n4625 , n5311 );
or ( n5314 , n4628 , n5312 , n5313 );
and ( n5315 , n4623 , n5314 );
and ( n5316 , n4621 , n5314 );
or ( n5317 , n4624 , n5315 , n5316 );
and ( n5318 , n4619 , n5317 );
and ( n5319 , n4617 , n5317 );
or ( n5320 , n4620 , n5318 , n5319 );
and ( n5321 , n4615 , n5320 );
and ( n5322 , n4613 , n5320 );
or ( n5323 , n4616 , n5321 , n5322 );
and ( n5324 , n4611 , n5323 );
and ( n5325 , n4609 , n5323 );
or ( n5326 , n4612 , n5324 , n5325 );
and ( n5327 , n4607 , n5326 );
and ( n5328 , n4605 , n5326 );
or ( n5329 , n4608 , n5327 , n5328 );
and ( n5330 , n4603 , n5329 );
and ( n5331 , n4601 , n5329 );
or ( n5332 , n4604 , n5330 , n5331 );
and ( n5333 , n4599 , n5332 );
and ( n5334 , n4597 , n5332 );
or ( n5335 , n4600 , n5333 , n5334 );
and ( n5336 , n4595 , n5335 );
and ( n5337 , n4593 , n5335 );
or ( n5338 , n4596 , n5336 , n5337 );
and ( n5339 , n4591 , n5338 );
and ( n5340 , n4589 , n5338 );
or ( n5341 , n4592 , n5339 , n5340 );
and ( n5342 , n4587 , n5341 );
and ( n5343 , n4585 , n5341 );
or ( n5344 , n4588 , n5342 , n5343 );
and ( n5345 , n4583 , n5344 );
and ( n5346 , n4581 , n5344 );
or ( n5347 , n4584 , n5345 , n5346 );
and ( n5348 , n4579 , n5347 );
and ( n5349 , n4577 , n5347 );
or ( n5350 , n4580 , n5348 , n5349 );
and ( n5351 , n4575 , n5350 );
and ( n5352 , n4573 , n5350 );
or ( n5353 , n4576 , n5351 , n5352 );
and ( n5354 , n4571 , n5353 );
and ( n5355 , n4569 , n5353 );
or ( n5356 , n4572 , n5354 , n5355 );
and ( n5357 , n4567 , n5356 );
and ( n5358 , n4565 , n5356 );
or ( n5359 , n4568 , n5357 , n5358 );
and ( n5360 , n4563 , n5359 );
and ( n5361 , n4561 , n5359 );
or ( n5362 , n4564 , n5360 , n5361 );
and ( n5363 , n4559 , n5362 );
and ( n5364 , n4557 , n5362 );
or ( n5365 , n4560 , n5363 , n5364 );
and ( n5366 , n4555 , n5365 );
and ( n5367 , n4553 , n5365 );
or ( n5368 , n4556 , n5366 , n5367 );
and ( n5369 , n4551 , n5368 );
and ( n5370 , n4549 , n5368 );
or ( n5371 , n4552 , n5369 , n5370 );
and ( n5372 , n4547 , n5371 );
and ( n5373 , n4545 , n5371 );
or ( n5374 , n4548 , n5372 , n5373 );
and ( n5375 , n4543 , n5374 );
and ( n5376 , n4541 , n5374 );
or ( n5377 , n4544 , n5375 , n5376 );
and ( n5378 , n4539 , n5377 );
and ( n5379 , n4537 , n5377 );
or ( n5380 , n4540 , n5378 , n5379 );
and ( n5381 , n4535 , n5380 );
and ( n5382 , n4533 , n5380 );
or ( n5383 , n4536 , n5381 , n5382 );
and ( n5384 , n4531 , n5383 );
and ( n5385 , n4529 , n5383 );
or ( n5386 , n4532 , n5384 , n5385 );
and ( n5387 , n4527 , n5386 );
and ( n5388 , n4525 , n5386 );
or ( n5389 , n4528 , n5387 , n5388 );
and ( n5390 , n4523 , n5389 );
and ( n5391 , n4521 , n5389 );
or ( n5392 , n4524 , n5390 , n5391 );
and ( n5393 , n4519 , n5392 );
and ( n5394 , n4517 , n5392 );
or ( n5395 , n4520 , n5393 , n5394 );
and ( n5396 , n4515 , n5395 );
and ( n5397 , n4513 , n5395 );
or ( n5398 , n4516 , n5396 , n5397 );
and ( n5399 , n4511 , n5398 );
and ( n5400 , n4509 , n5398 );
or ( n5401 , n4512 , n5399 , n5400 );
and ( n5402 , n4507 , n5401 );
and ( n5403 , n4505 , n5401 );
or ( n5404 , n4508 , n5402 , n5403 );
and ( n5405 , n4503 , n5404 );
and ( n5406 , n4501 , n5404 );
or ( n5407 , n4504 , n5405 , n5406 );
and ( n5408 , n4499 , n5407 );
and ( n5409 , n4497 , n5407 );
or ( n5410 , n4500 , n5408 , n5409 );
and ( n5411 , n4495 , n5410 );
and ( n5412 , n4493 , n5410 );
or ( n5413 , n4496 , n5411 , n5412 );
and ( n5414 , n4491 , n5413 );
and ( n5415 , n4489 , n5413 );
or ( n5416 , n4492 , n5414 , n5415 );
and ( n5417 , n4487 , n5416 );
and ( n5418 , n4485 , n5416 );
or ( n5419 , n4488 , n5417 , n5418 );
and ( n5420 , n4483 , n5419 );
and ( n5421 , n4481 , n5419 );
or ( n5422 , n4484 , n5420 , n5421 );
and ( n5423 , n4479 , n5422 );
and ( n5424 , n4477 , n5422 );
or ( n5425 , n4480 , n5423 , n5424 );
and ( n5426 , n4475 , n5425 );
and ( n5427 , n4473 , n5425 );
or ( n5428 , n4476 , n5426 , n5427 );
and ( n5429 , n4471 , n5428 );
and ( n5430 , n4469 , n5428 );
or ( n5431 , n4472 , n5429 , n5430 );
and ( n5432 , n4467 , n5431 );
and ( n5433 , n4465 , n5431 );
or ( n5434 , n4468 , n5432 , n5433 );
and ( n5435 , n4463 , n5434 );
and ( n5436 , n4461 , n5434 );
or ( n5437 , n4464 , n5435 , n5436 );
and ( n5438 , n4459 , n5437 );
and ( n5439 , n4457 , n5437 );
or ( n5440 , n4460 , n5438 , n5439 );
and ( n5441 , n4455 , n5440 );
and ( n5442 , n4453 , n5440 );
or ( n5443 , n4456 , n5441 , n5442 );
and ( n5444 , n4451 , n5443 );
and ( n5445 , n4449 , n5443 );
or ( n5446 , n4452 , n5444 , n5445 );
and ( n5447 , n4447 , n5446 );
and ( n5448 , n4445 , n5446 );
or ( n5449 , n4448 , n5447 , n5448 );
and ( n5450 , n4443 , n5449 );
and ( n5451 , n4441 , n5449 );
or ( n5452 , n4444 , n5450 , n5451 );
and ( n5453 , n4439 , n5452 );
and ( n5454 , n4437 , n5452 );
or ( n5455 , n4440 , n5453 , n5454 );
and ( n5456 , n4435 , n5455 );
and ( n5457 , n4433 , n5455 );
or ( n5458 , n4436 , n5456 , n5457 );
and ( n5459 , n4431 , n5458 );
and ( n5460 , n4429 , n5458 );
or ( n5461 , n4432 , n5459 , n5460 );
and ( n5462 , n4427 , n5461 );
and ( n5463 , n4425 , n5461 );
or ( n5464 , n4428 , n5462 , n5463 );
and ( n5465 , n4423 , n5464 );
and ( n5466 , n4421 , n5464 );
or ( n5467 , n4424 , n5465 , n5466 );
and ( n5468 , n4419 , n5467 );
and ( n5469 , n4417 , n5467 );
or ( n5470 , n4420 , n5468 , n5469 );
and ( n5471 , n4415 , n5470 );
and ( n5472 , n4413 , n5470 );
or ( n5473 , n4416 , n5471 , n5472 );
and ( n5474 , n4411 , n5473 );
and ( n5475 , n4409 , n5473 );
or ( n5476 , n4412 , n5474 , n5475 );
and ( n5477 , n4407 , n5476 );
and ( n5478 , n4405 , n5476 );
or ( n5479 , n4408 , n5477 , n5478 );
and ( n5480 , n4403 , n5479 );
and ( n5481 , n4401 , n5479 );
or ( n5482 , n4404 , n5480 , n5481 );
and ( n5483 , n4399 , n5482 );
and ( n5484 , n4397 , n5482 );
or ( n5485 , n4400 , n5483 , n5484 );
and ( n5486 , n4395 , n5485 );
and ( n5487 , n4393 , n5485 );
or ( n5488 , n4396 , n5486 , n5487 );
and ( n5489 , n4391 , n5488 );
and ( n5490 , n4389 , n5488 );
or ( n5491 , n4392 , n5489 , n5490 );
and ( n5492 , n4387 , n5491 );
and ( n5493 , n4385 , n5491 );
or ( n5494 , n4388 , n5492 , n5493 );
and ( n5495 , n4383 , n5494 );
and ( n5496 , n4381 , n5494 );
or ( n5497 , n4384 , n5495 , n5496 );
and ( n5498 , n4379 , n5497 );
and ( n5499 , n4377 , n5497 );
or ( n5500 , n4380 , n5498 , n5499 );
and ( n5501 , n4375 , n5500 );
and ( n5502 , n4373 , n5500 );
or ( n5503 , n4376 , n5501 , n5502 );
and ( n5504 , n4371 , n5503 );
and ( n5505 , n4369 , n5503 );
or ( n5506 , n4372 , n5504 , n5505 );
and ( n5507 , n4367 , n5506 );
and ( n5508 , n4365 , n5506 );
or ( n5509 , n4368 , n5507 , n5508 );
and ( n5510 , n4363 , n5509 );
and ( n5511 , n4361 , n5509 );
or ( n5512 , n4364 , n5510 , n5511 );
and ( n5513 , n4359 , n5512 );
and ( n5514 , n4357 , n5512 );
or ( n5515 , n4360 , n5513 , n5514 );
and ( n5516 , n4355 , n5515 );
and ( n5517 , n4353 , n5515 );
or ( n5518 , n4356 , n5516 , n5517 );
and ( n5519 , n4351 , n5518 );
and ( n5520 , n4349 , n5518 );
or ( n5521 , n4352 , n5519 , n5520 );
and ( n5522 , n4347 , n5521 );
and ( n5523 , n4345 , n5521 );
or ( n5524 , n4348 , n5522 , n5523 );
and ( n5525 , n4343 , n5524 );
and ( n5526 , n4341 , n5524 );
or ( n5527 , n4344 , n5525 , n5526 );
and ( n5528 , n4339 , n5527 );
and ( n5529 , n4337 , n5527 );
or ( n5530 , n4340 , n5528 , n5529 );
and ( n5531 , n4335 , n5530 );
and ( n5532 , n4333 , n5530 );
or ( n5533 , n4336 , n5531 , n5532 );
and ( n5534 , n4331 , n5533 );
and ( n5535 , n4329 , n5533 );
or ( n5536 , n4332 , n5534 , n5535 );
and ( n5537 , n4327 , n5536 );
and ( n5538 , n4325 , n5536 );
or ( n5539 , n4328 , n5537 , n5538 );
and ( n5540 , n4323 , n5539 );
and ( n5541 , n4321 , n5539 );
or ( n5542 , n4324 , n5540 , n5541 );
and ( n5543 , n4319 , n5542 );
and ( n5544 , n4317 , n5542 );
or ( n5545 , n4320 , n5543 , n5544 );
and ( n5546 , n4315 , n5545 );
and ( n5547 , n4313 , n5545 );
or ( n5548 , n4316 , n5546 , n5547 );
and ( n5549 , n4311 , n5548 );
and ( n5550 , n4309 , n5548 );
or ( n5551 , n4312 , n5549 , n5550 );
and ( n5552 , n4307 , n5551 );
and ( n5553 , n4305 , n5551 );
or ( n5554 , n4308 , n5552 , n5553 );
and ( n5555 , n4303 , n5554 );
and ( n5556 , n4301 , n5554 );
or ( n5557 , n4304 , n5555 , n5556 );
and ( n5558 , n4299 , n5557 );
and ( n5559 , n4297 , n5557 );
or ( n5560 , n4300 , n5558 , n5559 );
and ( n5561 , n4295 , n5560 );
and ( n5562 , n4293 , n5560 );
or ( n5563 , n4296 , n5561 , n5562 );
and ( n5564 , n4291 , n5563 );
and ( n5565 , n4289 , n5563 );
or ( n5566 , n4292 , n5564 , n5565 );
and ( n5567 , n4287 , n5566 );
and ( n5568 , n4285 , n5566 );
or ( n5569 , n4288 , n5567 , n5568 );
and ( n5570 , n4283 , n5569 );
and ( n5571 , n4281 , n5569 );
or ( n5572 , n4284 , n5570 , n5571 );
and ( n5573 , n4279 , n5572 );
and ( n5574 , n4277 , n5572 );
or ( n5575 , n4280 , n5573 , n5574 );
and ( n5576 , n4275 , n5575 );
and ( n5577 , n4273 , n5575 );
or ( n5578 , n4276 , n5576 , n5577 );
and ( n5579 , n4271 , n5578 );
and ( n5580 , n4269 , n5578 );
or ( n5581 , n4272 , n5579 , n5580 );
and ( n5582 , n4267 , n5581 );
and ( n5583 , n4265 , n5581 );
or ( n5584 , n4268 , n5582 , n5583 );
and ( n5585 , n4263 , n5584 );
and ( n5586 , n4261 , n5584 );
or ( n5587 , n4264 , n5585 , n5586 );
and ( n5588 , n4259 , n5587 );
and ( n5589 , n4257 , n5587 );
or ( n5590 , n4260 , n5588 , n5589 );
and ( n5591 , n4255 , n5590 );
and ( n5592 , n4253 , n5590 );
or ( n5593 , n4256 , n5591 , n5592 );
and ( n5594 , n4251 , n5593 );
and ( n5595 , n4249 , n5593 );
or ( n5596 , n4252 , n5594 , n5595 );
and ( n5597 , n4247 , n5596 );
and ( n5598 , n4245 , n5596 );
or ( n5599 , n4248 , n5597 , n5598 );
and ( n5600 , n4243 , n5599 );
and ( n5601 , n4241 , n5599 );
or ( n5602 , n4244 , n5600 , n5601 );
and ( n5603 , n4239 , n5602 );
and ( n5604 , n4237 , n5602 );
or ( n5605 , n4240 , n5603 , n5604 );
and ( n5606 , n4235 , n5605 );
and ( n5607 , n4233 , n5605 );
or ( n5608 , n4236 , n5606 , n5607 );
and ( n5609 , n4231 , n5608 );
and ( n5610 , n4229 , n5608 );
or ( n5611 , n4232 , n5609 , n5610 );
and ( n5612 , n4227 , n5611 );
and ( n5613 , n4225 , n5611 );
or ( n5614 , n4228 , n5612 , n5613 );
and ( n5615 , n4223 , n5614 );
and ( n5616 , n4221 , n5614 );
or ( n5617 , n4224 , n5615 , n5616 );
and ( n5618 , n4219 , n5617 );
and ( n5619 , n4217 , n5617 );
or ( n5620 , n4220 , n5618 , n5619 );
and ( n5621 , n4215 , n5620 );
and ( n5622 , n4213 , n5620 );
or ( n5623 , n4216 , n5621 , n5622 );
and ( n5624 , n4211 , n5623 );
and ( n5625 , n4209 , n5623 );
or ( n5626 , n4212 , n5624 , n5625 );
and ( n5627 , n4207 , n5626 );
and ( n5628 , n4205 , n5626 );
or ( n5629 , n4208 , n5627 , n5628 );
and ( n5630 , n4203 , n5629 );
and ( n5631 , n4201 , n5629 );
or ( n5632 , n4204 , n5630 , n5631 );
and ( n5633 , n4199 , n5632 );
and ( n5634 , n4197 , n5632 );
or ( n5635 , n4200 , n5633 , n5634 );
and ( n5636 , n4195 , n5635 );
and ( n5637 , n4193 , n5635 );
or ( n5638 , n4196 , n5636 , n5637 );
and ( n5639 , n4191 , n5638 );
and ( n5640 , n4189 , n5638 );
or ( n5641 , n4192 , n5639 , n5640 );
and ( n5642 , n4187 , n5641 );
and ( n5643 , n4185 , n5641 );
or ( n5644 , n4188 , n5642 , n5643 );
and ( n5645 , n4183 , n5644 );
and ( n5646 , n4181 , n5644 );
or ( n5647 , n4184 , n5645 , n5646 );
and ( n5648 , n4179 , n5647 );
and ( n5649 , n4177 , n5647 );
or ( n5650 , n4180 , n5648 , n5649 );
and ( n5651 , n4175 , n5650 );
and ( n5652 , n4173 , n5650 );
or ( n5653 , n4176 , n5651 , n5652 );
and ( n5654 , n4171 , n5653 );
and ( n5655 , n4169 , n5653 );
or ( n5656 , n4172 , n5654 , n5655 );
and ( n5657 , n4167 , n5656 );
and ( n5658 , n4165 , n5656 );
or ( n5659 , n4168 , n5657 , n5658 );
and ( n5660 , n4163 , n5659 );
and ( n5661 , n4161 , n5659 );
or ( n5662 , n4164 , n5660 , n5661 );
and ( n5663 , n4159 , n5662 );
and ( n5664 , n4157 , n5662 );
or ( n5665 , n4160 , n5663 , n5664 );
and ( n5666 , n4155 , n5665 );
and ( n5667 , n4153 , n5665 );
or ( n5668 , n4156 , n5666 , n5667 );
and ( n5669 , n4151 , n5668 );
and ( n5670 , n4149 , n5668 );
or ( n5671 , n4152 , n5669 , n5670 );
and ( n5672 , n4147 , n5671 );
and ( n5673 , n4145 , n5671 );
or ( n5674 , n4148 , n5672 , n5673 );
and ( n5675 , n4143 , n5674 );
and ( n5676 , n4141 , n5674 );
or ( n5677 , n4144 , n5675 , n5676 );
and ( n5678 , n4139 , n5677 );
and ( n5679 , n4137 , n5677 );
or ( n5680 , n4140 , n5678 , n5679 );
and ( n5681 , n4135 , n5680 );
and ( n5682 , n4133 , n5680 );
or ( n5683 , n4136 , n5681 , n5682 );
and ( n5684 , n4131 , n5683 );
and ( n5685 , n4129 , n5683 );
or ( n5686 , n4132 , n5684 , n5685 );
and ( n5687 , n4127 , n5686 );
and ( n5688 , n4125 , n5686 );
or ( n5689 , n4128 , n5687 , n5688 );
and ( n5690 , n4123 , n5689 );
and ( n5691 , n4121 , n5689 );
or ( n5692 , n4124 , n5690 , n5691 );
and ( n5693 , n4119 , n5692 );
and ( n5694 , n4117 , n5692 );
or ( n5695 , n4120 , n5693 , n5694 );
and ( n5696 , n4115 , n5695 );
and ( n5697 , n4113 , n5695 );
or ( n5698 , n4116 , n5696 , n5697 );
and ( n5699 , n4111 , n5698 );
and ( n5700 , n4109 , n5698 );
or ( n5701 , n4112 , n5699 , n5700 );
and ( n5702 , n4107 , n5701 );
and ( n5703 , n4105 , n5701 );
or ( n5704 , n4108 , n5702 , n5703 );
and ( n5705 , n4103 , n5704 );
and ( n5706 , n4101 , n5704 );
or ( n5707 , n4104 , n5705 , n5706 );
and ( n5708 , n4099 , n5707 );
and ( n5709 , n4097 , n5707 );
or ( n5710 , n4100 , n5708 , n5709 );
and ( n5711 , n4095 , n5710 );
and ( n5712 , n4093 , n5710 );
or ( n5713 , n4096 , n5711 , n5712 );
and ( n5714 , n4091 , n5713 );
and ( n5715 , n4089 , n5713 );
or ( n5716 , n4092 , n5714 , n5715 );
and ( n5717 , n4087 , n5716 );
and ( n5718 , n4085 , n5716 );
or ( n5719 , n4088 , n5717 , n5718 );
and ( n5720 , n4083 , n5719 );
and ( n5721 , n4081 , n5719 );
or ( n5722 , n4084 , n5720 , n5721 );
and ( n5723 , n4079 , n5722 );
and ( n5724 , n4077 , n5722 );
or ( n5725 , n4080 , n5723 , n5724 );
and ( n5726 , n4075 , n5725 );
and ( n5727 , n4073 , n5725 );
or ( n5728 , n4076 , n5726 , n5727 );
and ( n5729 , n4071 , n5728 );
and ( n5730 , n4069 , n5728 );
or ( n5731 , n4072 , n5729 , n5730 );
and ( n5732 , n4067 , n5731 );
and ( n5733 , n4065 , n5731 );
or ( n5734 , n4068 , n5732 , n5733 );
and ( n5735 , n4063 , n5734 );
and ( n5736 , n4061 , n5734 );
or ( n5737 , n4064 , n5735 , n5736 );
and ( n5738 , n4059 , n5737 );
and ( n5739 , n4057 , n5737 );
or ( n5740 , n4060 , n5738 , n5739 );
and ( n5741 , n4055 , n5740 );
and ( n5742 , n4053 , n5740 );
or ( n5743 , n4056 , n5741 , n5742 );
and ( n5744 , n4051 , n5743 );
and ( n5745 , n4049 , n5743 );
or ( n5746 , n4052 , n5744 , n5745 );
and ( n5747 , n4047 , n5746 );
and ( n5748 , n4045 , n5746 );
or ( n5749 , n4048 , n5747 , n5748 );
and ( n5750 , n4043 , n5749 );
and ( n5751 , n4041 , n5749 );
or ( n5752 , n4044 , n5750 , n5751 );
and ( n5753 , n4039 , n5752 );
and ( n5754 , n4037 , n5752 );
or ( n5755 , n4040 , n5753 , n5754 );
and ( n5756 , n4035 , n5755 );
and ( n5757 , n4033 , n5755 );
or ( n5758 , n4036 , n5756 , n5757 );
and ( n5759 , n4031 , n5758 );
and ( n5760 , n4029 , n5758 );
or ( n5761 , n4032 , n5759 , n5760 );
and ( n5762 , n4027 , n5761 );
and ( n5763 , n4025 , n5761 );
or ( n5764 , n4028 , n5762 , n5763 );
and ( n5765 , n4023 , n5764 );
and ( n5766 , n4021 , n5764 );
or ( n5767 , n4024 , n5765 , n5766 );
and ( n5768 , n4019 , n5767 );
and ( n5769 , n4017 , n5767 );
or ( n5770 , n4020 , n5768 , n5769 );
and ( n5771 , n4015 , n5770 );
and ( n5772 , n4013 , n5770 );
or ( n5773 , n4016 , n5771 , n5772 );
and ( n5774 , n4011 , n5773 );
and ( n5775 , n4009 , n5773 );
or ( n5776 , n4012 , n5774 , n5775 );
and ( n5777 , n4007 , n5776 );
and ( n5778 , n4005 , n5776 );
or ( n5779 , n4008 , n5777 , n5778 );
and ( n5780 , n4003 , n5779 );
and ( n5781 , n4001 , n5779 );
or ( n5782 , n4004 , n5780 , n5781 );
xor ( n5783 , n4000 , n5782 );
buf ( n5784 , n5783 );
xor ( n5785 , n4001 , n4003 );
xor ( n5786 , n5785 , n5779 );
buf ( n5787 , n5786 );
xor ( n5788 , n5784 , n5787 );
xor ( n5789 , n4005 , n4007 );
xor ( n5790 , n5789 , n5776 );
buf ( n5791 , n5790 );
xor ( n5792 , n4009 , n4011 );
xor ( n5793 , n5792 , n5773 );
buf ( n5794 , n5793 );
xor ( n5795 , n5791 , n5794 );
xor ( n5796 , n5788 , n5795 );
xor ( n5797 , n4013 , n4015 );
xor ( n5798 , n5797 , n5770 );
buf ( n5799 , n5798 );
xor ( n5800 , n4017 , n4019 );
xor ( n5801 , n5800 , n5767 );
buf ( n5802 , n5801 );
xor ( n5803 , n5799 , n5802 );
xor ( n5804 , n4021 , n4023 );
xor ( n5805 , n5804 , n5764 );
buf ( n5806 , n5805 );
xor ( n5807 , n4025 , n4027 );
xor ( n5808 , n5807 , n5761 );
buf ( n5809 , n5808 );
xor ( n5810 , n5806 , n5809 );
xor ( n5811 , n5803 , n5810 );
xor ( n5812 , n5796 , n5811 );
xor ( n5813 , n4029 , n4031 );
xor ( n5814 , n5813 , n5758 );
buf ( n5815 , n5814 );
xor ( n5816 , n4033 , n4035 );
xor ( n5817 , n5816 , n5755 );
buf ( n5818 , n5817 );
xor ( n5819 , n5815 , n5818 );
xor ( n5820 , n4037 , n4039 );
xor ( n5821 , n5820 , n5752 );
buf ( n5822 , n5821 );
xor ( n5823 , n4041 , n4043 );
xor ( n5824 , n5823 , n5749 );
buf ( n5825 , n5824 );
xor ( n5826 , n5822 , n5825 );
xor ( n5827 , n5819 , n5826 );
xor ( n5828 , n4045 , n4047 );
xor ( n5829 , n5828 , n5746 );
buf ( n5830 , n5829 );
xor ( n5831 , n4049 , n4051 );
xor ( n5832 , n5831 , n5743 );
buf ( n5833 , n5832 );
xor ( n5834 , n5830 , n5833 );
xor ( n5835 , n4053 , n4055 );
xor ( n5836 , n5835 , n5740 );
buf ( n5837 , n5836 );
xor ( n5838 , n4057 , n4059 );
xor ( n5839 , n5838 , n5737 );
buf ( n5840 , n5839 );
xor ( n5841 , n5837 , n5840 );
xor ( n5842 , n5834 , n5841 );
xor ( n5843 , n5827 , n5842 );
xor ( n5844 , n5812 , n5843 );
xor ( n5845 , n4061 , n4063 );
xor ( n5846 , n5845 , n5734 );
buf ( n5847 , n5846 );
xor ( n5848 , n4065 , n4067 );
xor ( n5849 , n5848 , n5731 );
buf ( n5850 , n5849 );
xor ( n5851 , n5847 , n5850 );
xor ( n5852 , n4069 , n4071 );
xor ( n5853 , n5852 , n5728 );
buf ( n5854 , n5853 );
xor ( n5855 , n4073 , n4075 );
xor ( n5856 , n5855 , n5725 );
buf ( n5857 , n5856 );
xor ( n5858 , n5854 , n5857 );
xor ( n5859 , n5851 , n5858 );
xor ( n5860 , n4077 , n4079 );
xor ( n5861 , n5860 , n5722 );
buf ( n5862 , n5861 );
xor ( n5863 , n4081 , n4083 );
xor ( n5864 , n5863 , n5719 );
buf ( n5865 , n5864 );
xor ( n5866 , n5862 , n5865 );
xor ( n5867 , n4085 , n4087 );
xor ( n5868 , n5867 , n5716 );
buf ( n5869 , n5868 );
xor ( n5870 , n4089 , n4091 );
xor ( n5871 , n5870 , n5713 );
buf ( n5872 , n5871 );
xor ( n5873 , n5869 , n5872 );
xor ( n5874 , n5866 , n5873 );
xor ( n5875 , n5859 , n5874 );
xor ( n5876 , n4093 , n4095 );
xor ( n5877 , n5876 , n5710 );
buf ( n5878 , n5877 );
xor ( n5879 , n4097 , n4099 );
xor ( n5880 , n5879 , n5707 );
buf ( n5881 , n5880 );
xor ( n5882 , n5878 , n5881 );
xor ( n5883 , n4101 , n4103 );
xor ( n5884 , n5883 , n5704 );
buf ( n5885 , n5884 );
xor ( n5886 , n4105 , n4107 );
xor ( n5887 , n5886 , n5701 );
buf ( n5888 , n5887 );
xor ( n5889 , n5885 , n5888 );
xor ( n5890 , n5882 , n5889 );
xor ( n5891 , n4109 , n4111 );
xor ( n5892 , n5891 , n5698 );
buf ( n5893 , n5892 );
xor ( n5894 , n4113 , n4115 );
xor ( n5895 , n5894 , n5695 );
buf ( n5896 , n5895 );
xor ( n5897 , n5893 , n5896 );
xor ( n5898 , n4117 , n4119 );
xor ( n5899 , n5898 , n5692 );
buf ( n5900 , n5899 );
xor ( n5901 , n4121 , n4123 );
xor ( n5902 , n5901 , n5689 );
buf ( n5903 , n5902 );
xor ( n5904 , n5900 , n5903 );
xor ( n5905 , n5897 , n5904 );
xor ( n5906 , n5890 , n5905 );
xor ( n5907 , n5875 , n5906 );
xor ( n5908 , n5844 , n5907 );
xor ( n5909 , n4125 , n4127 );
xor ( n5910 , n5909 , n5686 );
buf ( n5911 , n5910 );
xor ( n5912 , n4129 , n4131 );
xor ( n5913 , n5912 , n5683 );
buf ( n5914 , n5913 );
xor ( n5915 , n5911 , n5914 );
xor ( n5916 , n4133 , n4135 );
xor ( n5917 , n5916 , n5680 );
buf ( n5918 , n5917 );
xor ( n5919 , n4137 , n4139 );
xor ( n5920 , n5919 , n5677 );
buf ( n5921 , n5920 );
xor ( n5922 , n5918 , n5921 );
xor ( n5923 , n5915 , n5922 );
xor ( n5924 , n4141 , n4143 );
xor ( n5925 , n5924 , n5674 );
buf ( n5926 , n5925 );
xor ( n5927 , n4145 , n4147 );
xor ( n5928 , n5927 , n5671 );
buf ( n5929 , n5928 );
xor ( n5930 , n5926 , n5929 );
xor ( n5931 , n4149 , n4151 );
xor ( n5932 , n5931 , n5668 );
buf ( n5933 , n5932 );
xor ( n5934 , n4153 , n4155 );
xor ( n5935 , n5934 , n5665 );
buf ( n5936 , n5935 );
xor ( n5937 , n5933 , n5936 );
xor ( n5938 , n5930 , n5937 );
xor ( n5939 , n5923 , n5938 );
xor ( n5940 , n4157 , n4159 );
xor ( n5941 , n5940 , n5662 );
buf ( n5942 , n5941 );
xor ( n5943 , n4161 , n4163 );
xor ( n5944 , n5943 , n5659 );
buf ( n5945 , n5944 );
xor ( n5946 , n5942 , n5945 );
xor ( n5947 , n4165 , n4167 );
xor ( n5948 , n5947 , n5656 );
buf ( n5949 , n5948 );
xor ( n5950 , n4169 , n4171 );
xor ( n5951 , n5950 , n5653 );
buf ( n5952 , n5951 );
xor ( n5953 , n5949 , n5952 );
xor ( n5954 , n5946 , n5953 );
xor ( n5955 , n4173 , n4175 );
xor ( n5956 , n5955 , n5650 );
buf ( n5957 , n5956 );
xor ( n5958 , n4177 , n4179 );
xor ( n5959 , n5958 , n5647 );
buf ( n5960 , n5959 );
xor ( n5961 , n5957 , n5960 );
xor ( n5962 , n4181 , n4183 );
xor ( n5963 , n5962 , n5644 );
buf ( n5964 , n5963 );
xor ( n5965 , n4185 , n4187 );
xor ( n5966 , n5965 , n5641 );
buf ( n5967 , n5966 );
xor ( n5968 , n5964 , n5967 );
xor ( n5969 , n5961 , n5968 );
xor ( n5970 , n5954 , n5969 );
xor ( n5971 , n5939 , n5970 );
xor ( n5972 , n4189 , n4191 );
xor ( n5973 , n5972 , n5638 );
buf ( n5974 , n5973 );
xor ( n5975 , n4193 , n4195 );
xor ( n5976 , n5975 , n5635 );
buf ( n5977 , n5976 );
xor ( n5978 , n5974 , n5977 );
xor ( n5979 , n4197 , n4199 );
xor ( n5980 , n5979 , n5632 );
buf ( n5981 , n5980 );
xor ( n5982 , n4201 , n4203 );
xor ( n5983 , n5982 , n5629 );
buf ( n5984 , n5983 );
xor ( n5985 , n5981 , n5984 );
xor ( n5986 , n5978 , n5985 );
xor ( n5987 , n4205 , n4207 );
xor ( n5988 , n5987 , n5626 );
buf ( n5989 , n5988 );
xor ( n5990 , n4209 , n4211 );
xor ( n5991 , n5990 , n5623 );
buf ( n5992 , n5991 );
xor ( n5993 , n5989 , n5992 );
xor ( n5994 , n4213 , n4215 );
xor ( n5995 , n5994 , n5620 );
buf ( n5996 , n5995 );
xor ( n5997 , n4217 , n4219 );
xor ( n5998 , n5997 , n5617 );
buf ( n5999 , n5998 );
xor ( n6000 , n5996 , n5999 );
xor ( n6001 , n5993 , n6000 );
xor ( n6002 , n5986 , n6001 );
xor ( n6003 , n4221 , n4223 );
xor ( n6004 , n6003 , n5614 );
buf ( n6005 , n6004 );
xor ( n6006 , n4225 , n4227 );
xor ( n6007 , n6006 , n5611 );
buf ( n6008 , n6007 );
xor ( n6009 , n6005 , n6008 );
xor ( n6010 , n4229 , n4231 );
xor ( n6011 , n6010 , n5608 );
buf ( n6012 , n6011 );
xor ( n6013 , n4233 , n4235 );
xor ( n6014 , n6013 , n5605 );
buf ( n6015 , n6014 );
xor ( n6016 , n6012 , n6015 );
xor ( n6017 , n6009 , n6016 );
xor ( n6018 , n4237 , n4239 );
xor ( n6019 , n6018 , n5602 );
buf ( n6020 , n6019 );
xor ( n6021 , n4241 , n4243 );
xor ( n6022 , n6021 , n5599 );
buf ( n6023 , n6022 );
xor ( n6024 , n6020 , n6023 );
xor ( n6025 , n4245 , n4247 );
xor ( n6026 , n6025 , n5596 );
buf ( n6027 , n6026 );
xor ( n6028 , n4249 , n4251 );
xor ( n6029 , n6028 , n5593 );
buf ( n6030 , n6029 );
xor ( n6031 , n6027 , n6030 );
xor ( n6032 , n6024 , n6031 );
xor ( n6033 , n6017 , n6032 );
xor ( n6034 , n6002 , n6033 );
xor ( n6035 , n5971 , n6034 );
xor ( n6036 , n5908 , n6035 );
xor ( n6037 , n4253 , n4255 );
xor ( n6038 , n6037 , n5590 );
buf ( n6039 , n6038 );
xor ( n6040 , n4257 , n4259 );
xor ( n6041 , n6040 , n5587 );
buf ( n6042 , n6041 );
xor ( n6043 , n6039 , n6042 );
xor ( n6044 , n4261 , n4263 );
xor ( n6045 , n6044 , n5584 );
buf ( n6046 , n6045 );
xor ( n6047 , n4265 , n4267 );
xor ( n6048 , n6047 , n5581 );
buf ( n6049 , n6048 );
xor ( n6050 , n6046 , n6049 );
xor ( n6051 , n6043 , n6050 );
xor ( n6052 , n4269 , n4271 );
xor ( n6053 , n6052 , n5578 );
buf ( n6054 , n6053 );
xor ( n6055 , n4273 , n4275 );
xor ( n6056 , n6055 , n5575 );
buf ( n6057 , n6056 );
xor ( n6058 , n6054 , n6057 );
xor ( n6059 , n4277 , n4279 );
xor ( n6060 , n6059 , n5572 );
buf ( n6061 , n6060 );
xor ( n6062 , n4281 , n4283 );
xor ( n6063 , n6062 , n5569 );
buf ( n6064 , n6063 );
xor ( n6065 , n6061 , n6064 );
xor ( n6066 , n6058 , n6065 );
xor ( n6067 , n6051 , n6066 );
xor ( n6068 , n4285 , n4287 );
xor ( n6069 , n6068 , n5566 );
buf ( n6070 , n6069 );
xor ( n6071 , n4289 , n4291 );
xor ( n6072 , n6071 , n5563 );
buf ( n6073 , n6072 );
xor ( n6074 , n6070 , n6073 );
xor ( n6075 , n4293 , n4295 );
xor ( n6076 , n6075 , n5560 );
buf ( n6077 , n6076 );
xor ( n6078 , n4297 , n4299 );
xor ( n6079 , n6078 , n5557 );
buf ( n6080 , n6079 );
xor ( n6081 , n6077 , n6080 );
xor ( n6082 , n6074 , n6081 );
xor ( n6083 , n4301 , n4303 );
xor ( n6084 , n6083 , n5554 );
buf ( n6085 , n6084 );
xor ( n6086 , n4305 , n4307 );
xor ( n6087 , n6086 , n5551 );
buf ( n6088 , n6087 );
xor ( n6089 , n6085 , n6088 );
xor ( n6090 , n4309 , n4311 );
xor ( n6091 , n6090 , n5548 );
buf ( n6092 , n6091 );
xor ( n6093 , n4313 , n4315 );
xor ( n6094 , n6093 , n5545 );
buf ( n6095 , n6094 );
xor ( n6096 , n6092 , n6095 );
xor ( n6097 , n6089 , n6096 );
xor ( n6098 , n6082 , n6097 );
xor ( n6099 , n6067 , n6098 );
xor ( n6100 , n4317 , n4319 );
xor ( n6101 , n6100 , n5542 );
buf ( n6102 , n6101 );
xor ( n6103 , n4321 , n4323 );
xor ( n6104 , n6103 , n5539 );
buf ( n6105 , n6104 );
xor ( n6106 , n6102 , n6105 );
xor ( n6107 , n4325 , n4327 );
xor ( n6108 , n6107 , n5536 );
buf ( n6109 , n6108 );
xor ( n6110 , n4329 , n4331 );
xor ( n6111 , n6110 , n5533 );
buf ( n6112 , n6111 );
xor ( n6113 , n6109 , n6112 );
xor ( n6114 , n6106 , n6113 );
xor ( n6115 , n4333 , n4335 );
xor ( n6116 , n6115 , n5530 );
buf ( n6117 , n6116 );
xor ( n6118 , n4337 , n4339 );
xor ( n6119 , n6118 , n5527 );
buf ( n6120 , n6119 );
xor ( n6121 , n6117 , n6120 );
xor ( n6122 , n4341 , n4343 );
xor ( n6123 , n6122 , n5524 );
buf ( n6124 , n6123 );
xor ( n6125 , n4345 , n4347 );
xor ( n6126 , n6125 , n5521 );
buf ( n6127 , n6126 );
xor ( n6128 , n6124 , n6127 );
xor ( n6129 , n6121 , n6128 );
xor ( n6130 , n6114 , n6129 );
xor ( n6131 , n4349 , n4351 );
xor ( n6132 , n6131 , n5518 );
buf ( n6133 , n6132 );
xor ( n6134 , n4353 , n4355 );
xor ( n6135 , n6134 , n5515 );
buf ( n6136 , n6135 );
xor ( n6137 , n6133 , n6136 );
xor ( n6138 , n4357 , n4359 );
xor ( n6139 , n6138 , n5512 );
buf ( n6140 , n6139 );
xor ( n6141 , n4361 , n4363 );
xor ( n6142 , n6141 , n5509 );
buf ( n6143 , n6142 );
xor ( n6144 , n6140 , n6143 );
xor ( n6145 , n6137 , n6144 );
xor ( n6146 , n4365 , n4367 );
xor ( n6147 , n6146 , n5506 );
buf ( n6148 , n6147 );
xor ( n6149 , n4369 , n4371 );
xor ( n6150 , n6149 , n5503 );
buf ( n6151 , n6150 );
xor ( n6152 , n6148 , n6151 );
xor ( n6153 , n4373 , n4375 );
xor ( n6154 , n6153 , n5500 );
buf ( n6155 , n6154 );
xor ( n6156 , n4377 , n4379 );
xor ( n6157 , n6156 , n5497 );
buf ( n6158 , n6157 );
xor ( n6159 , n6155 , n6158 );
xor ( n6160 , n6152 , n6159 );
xor ( n6161 , n6145 , n6160 );
xor ( n6162 , n6130 , n6161 );
xor ( n6163 , n6099 , n6162 );
xor ( n6164 , n4381 , n4383 );
xor ( n6165 , n6164 , n5494 );
buf ( n6166 , n6165 );
xor ( n6167 , n4385 , n4387 );
xor ( n6168 , n6167 , n5491 );
buf ( n6169 , n6168 );
xor ( n6170 , n6166 , n6169 );
xor ( n6171 , n4389 , n4391 );
xor ( n6172 , n6171 , n5488 );
buf ( n6173 , n6172 );
xor ( n6174 , n4393 , n4395 );
xor ( n6175 , n6174 , n5485 );
buf ( n6176 , n6175 );
xor ( n6177 , n6173 , n6176 );
xor ( n6178 , n6170 , n6177 );
xor ( n6179 , n4397 , n4399 );
xor ( n6180 , n6179 , n5482 );
buf ( n6181 , n6180 );
xor ( n6182 , n4401 , n4403 );
xor ( n6183 , n6182 , n5479 );
buf ( n6184 , n6183 );
xor ( n6185 , n6181 , n6184 );
xor ( n6186 , n4405 , n4407 );
xor ( n6187 , n6186 , n5476 );
buf ( n6188 , n6187 );
xor ( n6189 , n4409 , n4411 );
xor ( n6190 , n6189 , n5473 );
buf ( n6191 , n6190 );
xor ( n6192 , n6188 , n6191 );
xor ( n6193 , n6185 , n6192 );
xor ( n6194 , n6178 , n6193 );
xor ( n6195 , n4413 , n4415 );
xor ( n6196 , n6195 , n5470 );
buf ( n6197 , n6196 );
xor ( n6198 , n4417 , n4419 );
xor ( n6199 , n6198 , n5467 );
buf ( n6200 , n6199 );
xor ( n6201 , n6197 , n6200 );
xor ( n6202 , n4421 , n4423 );
xor ( n6203 , n6202 , n5464 );
buf ( n6204 , n6203 );
xor ( n6205 , n4425 , n4427 );
xor ( n6206 , n6205 , n5461 );
buf ( n6207 , n6206 );
xor ( n6208 , n6204 , n6207 );
xor ( n6209 , n6201 , n6208 );
xor ( n6210 , n4429 , n4431 );
xor ( n6211 , n6210 , n5458 );
buf ( n6212 , n6211 );
xor ( n6213 , n4433 , n4435 );
xor ( n6214 , n6213 , n5455 );
buf ( n6215 , n6214 );
xor ( n6216 , n6212 , n6215 );
xor ( n6217 , n4437 , n4439 );
xor ( n6218 , n6217 , n5452 );
buf ( n6219 , n6218 );
xor ( n6220 , n4441 , n4443 );
xor ( n6221 , n6220 , n5449 );
buf ( n6222 , n6221 );
xor ( n6223 , n6219 , n6222 );
xor ( n6224 , n6216 , n6223 );
xor ( n6225 , n6209 , n6224 );
xor ( n6226 , n6194 , n6225 );
xor ( n6227 , n4445 , n4447 );
xor ( n6228 , n6227 , n5446 );
buf ( n6229 , n6228 );
xor ( n6230 , n4449 , n4451 );
xor ( n6231 , n6230 , n5443 );
buf ( n6232 , n6231 );
xor ( n6233 , n6229 , n6232 );
xor ( n6234 , n4453 , n4455 );
xor ( n6235 , n6234 , n5440 );
buf ( n6236 , n6235 );
xor ( n6237 , n4457 , n4459 );
xor ( n6238 , n6237 , n5437 );
buf ( n6239 , n6238 );
xor ( n6240 , n6236 , n6239 );
xor ( n6241 , n6233 , n6240 );
xor ( n6242 , n4461 , n4463 );
xor ( n6243 , n6242 , n5434 );
buf ( n6244 , n6243 );
xor ( n6245 , n4465 , n4467 );
xor ( n6246 , n6245 , n5431 );
buf ( n6247 , n6246 );
xor ( n6248 , n6244 , n6247 );
xor ( n6249 , n4469 , n4471 );
xor ( n6250 , n6249 , n5428 );
buf ( n6251 , n6250 );
xor ( n6252 , n4473 , n4475 );
xor ( n6253 , n6252 , n5425 );
buf ( n6254 , n6253 );
xor ( n6255 , n6251 , n6254 );
xor ( n6256 , n6248 , n6255 );
xor ( n6257 , n6241 , n6256 );
xor ( n6258 , n4477 , n4479 );
xor ( n6259 , n6258 , n5422 );
buf ( n6260 , n6259 );
xor ( n6261 , n4481 , n4483 );
xor ( n6262 , n6261 , n5419 );
buf ( n6263 , n6262 );
xor ( n6264 , n6260 , n6263 );
xor ( n6265 , n4485 , n4487 );
xor ( n6266 , n6265 , n5416 );
buf ( n6267 , n6266 );
xor ( n6268 , n4489 , n4491 );
xor ( n6269 , n6268 , n5413 );
buf ( n6270 , n6269 );
xor ( n6271 , n6267 , n6270 );
xor ( n6272 , n6264 , n6271 );
xor ( n6273 , n4493 , n4495 );
xor ( n6274 , n6273 , n5410 );
buf ( n6275 , n6274 );
xor ( n6276 , n4497 , n4499 );
xor ( n6277 , n6276 , n5407 );
buf ( n6278 , n6277 );
xor ( n6279 , n6275 , n6278 );
xor ( n6280 , n4501 , n4503 );
xor ( n6281 , n6280 , n5404 );
buf ( n6282 , n6281 );
xor ( n6283 , n4505 , n4507 );
xor ( n6284 , n6283 , n5401 );
buf ( n6285 , n6284 );
xor ( n6286 , n6282 , n6285 );
xor ( n6287 , n6279 , n6286 );
xor ( n6288 , n6272 , n6287 );
xor ( n6289 , n6257 , n6288 );
xor ( n6290 , n6226 , n6289 );
xor ( n6291 , n6163 , n6290 );
xor ( n6292 , n6036 , n6291 );
xor ( n6293 , n4509 , n4511 );
xor ( n6294 , n6293 , n5398 );
buf ( n6295 , n6294 );
xor ( n6296 , n4513 , n4515 );
xor ( n6297 , n6296 , n5395 );
buf ( n6298 , n6297 );
xor ( n6299 , n6295 , n6298 );
xor ( n6300 , n4517 , n4519 );
xor ( n6301 , n6300 , n5392 );
buf ( n6302 , n6301 );
xor ( n6303 , n4521 , n4523 );
xor ( n6304 , n6303 , n5389 );
buf ( n6305 , n6304 );
xor ( n6306 , n6302 , n6305 );
xor ( n6307 , n6299 , n6306 );
xor ( n6308 , n4525 , n4527 );
xor ( n6309 , n6308 , n5386 );
buf ( n6310 , n6309 );
xor ( n6311 , n4529 , n4531 );
xor ( n6312 , n6311 , n5383 );
buf ( n6313 , n6312 );
xor ( n6314 , n6310 , n6313 );
xor ( n6315 , n4533 , n4535 );
xor ( n6316 , n6315 , n5380 );
buf ( n6317 , n6316 );
xor ( n6318 , n4537 , n4539 );
xor ( n6319 , n6318 , n5377 );
buf ( n6320 , n6319 );
xor ( n6321 , n6317 , n6320 );
xor ( n6322 , n6314 , n6321 );
xor ( n6323 , n6307 , n6322 );
xor ( n6324 , n4541 , n4543 );
xor ( n6325 , n6324 , n5374 );
buf ( n6326 , n6325 );
xor ( n6327 , n4545 , n4547 );
xor ( n6328 , n6327 , n5371 );
buf ( n6329 , n6328 );
xor ( n6330 , n6326 , n6329 );
xor ( n6331 , n4549 , n4551 );
xor ( n6332 , n6331 , n5368 );
buf ( n6333 , n6332 );
xor ( n6334 , n4553 , n4555 );
xor ( n6335 , n6334 , n5365 );
buf ( n6336 , n6335 );
xor ( n6337 , n6333 , n6336 );
xor ( n6338 , n6330 , n6337 );
xor ( n6339 , n4557 , n4559 );
xor ( n6340 , n6339 , n5362 );
buf ( n6341 , n6340 );
xor ( n6342 , n4561 , n4563 );
xor ( n6343 , n6342 , n5359 );
buf ( n6344 , n6343 );
xor ( n6345 , n6341 , n6344 );
xor ( n6346 , n4565 , n4567 );
xor ( n6347 , n6346 , n5356 );
buf ( n6348 , n6347 );
xor ( n6349 , n4569 , n4571 );
xor ( n6350 , n6349 , n5353 );
buf ( n6351 , n6350 );
xor ( n6352 , n6348 , n6351 );
xor ( n6353 , n6345 , n6352 );
xor ( n6354 , n6338 , n6353 );
xor ( n6355 , n6323 , n6354 );
xor ( n6356 , n4573 , n4575 );
xor ( n6357 , n6356 , n5350 );
buf ( n6358 , n6357 );
xor ( n6359 , n4577 , n4579 );
xor ( n6360 , n6359 , n5347 );
buf ( n6361 , n6360 );
xor ( n6362 , n6358 , n6361 );
xor ( n6363 , n4581 , n4583 );
xor ( n6364 , n6363 , n5344 );
buf ( n6365 , n6364 );
xor ( n6366 , n4585 , n4587 );
xor ( n6367 , n6366 , n5341 );
buf ( n6368 , n6367 );
xor ( n6369 , n6365 , n6368 );
xor ( n6370 , n6362 , n6369 );
xor ( n6371 , n4589 , n4591 );
xor ( n6372 , n6371 , n5338 );
buf ( n6373 , n6372 );
xor ( n6374 , n4593 , n4595 );
xor ( n6375 , n6374 , n5335 );
buf ( n6376 , n6375 );
xor ( n6377 , n6373 , n6376 );
xor ( n6378 , n4597 , n4599 );
xor ( n6379 , n6378 , n5332 );
buf ( n6380 , n6379 );
xor ( n6381 , n4601 , n4603 );
xor ( n6382 , n6381 , n5329 );
buf ( n6383 , n6382 );
xor ( n6384 , n6380 , n6383 );
xor ( n6385 , n6377 , n6384 );
xor ( n6386 , n6370 , n6385 );
xor ( n6387 , n4605 , n4607 );
xor ( n6388 , n6387 , n5326 );
buf ( n6389 , n6388 );
xor ( n6390 , n4609 , n4611 );
xor ( n6391 , n6390 , n5323 );
buf ( n6392 , n6391 );
xor ( n6393 , n6389 , n6392 );
xor ( n6394 , n4613 , n4615 );
xor ( n6395 , n6394 , n5320 );
buf ( n6396 , n6395 );
xor ( n6397 , n4617 , n4619 );
xor ( n6398 , n6397 , n5317 );
buf ( n6399 , n6398 );
xor ( n6400 , n6396 , n6399 );
xor ( n6401 , n6393 , n6400 );
xor ( n6402 , n4621 , n4623 );
xor ( n6403 , n6402 , n5314 );
buf ( n6404 , n6403 );
xor ( n6405 , n4625 , n4627 );
xor ( n6406 , n6405 , n5311 );
buf ( n6407 , n6406 );
xor ( n6408 , n6404 , n6407 );
xor ( n6409 , n4629 , n4631 );
xor ( n6410 , n6409 , n5308 );
buf ( n6411 , n6410 );
xor ( n6412 , n4633 , n4635 );
xor ( n6413 , n6412 , n5305 );
buf ( n6414 , n6413 );
xor ( n6415 , n6411 , n6414 );
xor ( n6416 , n6408 , n6415 );
xor ( n6417 , n6401 , n6416 );
xor ( n6418 , n6386 , n6417 );
xor ( n6419 , n6355 , n6418 );
xor ( n6420 , n4637 , n4639 );
xor ( n6421 , n6420 , n5302 );
buf ( n6422 , n6421 );
xor ( n6423 , n4641 , n4643 );
xor ( n6424 , n6423 , n5299 );
buf ( n6425 , n6424 );
xor ( n6426 , n6422 , n6425 );
xor ( n6427 , n4645 , n4647 );
xor ( n6428 , n6427 , n5296 );
buf ( n6429 , n6428 );
xor ( n6430 , n4649 , n4651 );
xor ( n6431 , n6430 , n5293 );
buf ( n6432 , n6431 );
xor ( n6433 , n6429 , n6432 );
xor ( n6434 , n6426 , n6433 );
xor ( n6435 , n4653 , n4655 );
xor ( n6436 , n6435 , n5290 );
buf ( n6437 , n6436 );
xor ( n6438 , n4657 , n4659 );
xor ( n6439 , n6438 , n5287 );
buf ( n6440 , n6439 );
xor ( n6441 , n6437 , n6440 );
xor ( n6442 , n4661 , n4663 );
xor ( n6443 , n6442 , n5284 );
buf ( n6444 , n6443 );
xor ( n6445 , n4665 , n4667 );
xor ( n6446 , n6445 , n5281 );
buf ( n6447 , n6446 );
xor ( n6448 , n6444 , n6447 );
xor ( n6449 , n6441 , n6448 );
xor ( n6450 , n6434 , n6449 );
xor ( n6451 , n4669 , n4671 );
xor ( n6452 , n6451 , n5278 );
buf ( n6453 , n6452 );
xor ( n6454 , n4673 , n4675 );
xor ( n6455 , n6454 , n5275 );
buf ( n6456 , n6455 );
xor ( n6457 , n6453 , n6456 );
xor ( n6458 , n4677 , n4679 );
xor ( n6459 , n6458 , n5272 );
buf ( n6460 , n6459 );
xor ( n6461 , n4681 , n4683 );
xor ( n6462 , n6461 , n5269 );
buf ( n6463 , n6462 );
xor ( n6464 , n6460 , n6463 );
xor ( n6465 , n6457 , n6464 );
xor ( n6466 , n4685 , n4687 );
xor ( n6467 , n6466 , n5266 );
buf ( n6468 , n6467 );
xor ( n6469 , n4689 , n4691 );
xor ( n6470 , n6469 , n5263 );
buf ( n6471 , n6470 );
xor ( n6472 , n6468 , n6471 );
xor ( n6473 , n4693 , n4695 );
xor ( n6474 , n6473 , n5260 );
buf ( n6475 , n6474 );
xor ( n6476 , n4697 , n4699 );
xor ( n6477 , n6476 , n5257 );
buf ( n6478 , n6477 );
xor ( n6479 , n6475 , n6478 );
xor ( n6480 , n6472 , n6479 );
xor ( n6481 , n6465 , n6480 );
xor ( n6482 , n6450 , n6481 );
xor ( n6483 , n4701 , n4703 );
xor ( n6484 , n6483 , n5254 );
buf ( n6485 , n6484 );
xor ( n6486 , n4705 , n4707 );
xor ( n6487 , n6486 , n5251 );
buf ( n6488 , n6487 );
xor ( n6489 , n6485 , n6488 );
xor ( n6490 , n4709 , n4711 );
xor ( n6491 , n6490 , n5248 );
buf ( n6492 , n6491 );
xor ( n6493 , n4713 , n4715 );
xor ( n6494 , n6493 , n5245 );
buf ( n6495 , n6494 );
xor ( n6496 , n6492 , n6495 );
xor ( n6497 , n6489 , n6496 );
xor ( n6498 , n4717 , n4719 );
xor ( n6499 , n6498 , n5242 );
buf ( n6500 , n6499 );
xor ( n6501 , n4721 , n4723 );
xor ( n6502 , n6501 , n5239 );
buf ( n6503 , n6502 );
xor ( n6504 , n6500 , n6503 );
xor ( n6505 , n4725 , n4727 );
xor ( n6506 , n6505 , n5236 );
buf ( n6507 , n6506 );
xor ( n6508 , n4729 , n4731 );
xor ( n6509 , n6508 , n5233 );
buf ( n6510 , n6509 );
xor ( n6511 , n6507 , n6510 );
xor ( n6512 , n6504 , n6511 );
xor ( n6513 , n6497 , n6512 );
xor ( n6514 , n4733 , n4735 );
xor ( n6515 , n6514 , n5230 );
buf ( n6516 , n6515 );
xor ( n6517 , n4737 , n4739 );
xor ( n6518 , n6517 , n5227 );
buf ( n6519 , n6518 );
xor ( n6520 , n6516 , n6519 );
xor ( n6521 , n4741 , n4743 );
xor ( n6522 , n6521 , n5224 );
buf ( n6523 , n6522 );
xor ( n6524 , n4745 , n4747 );
xor ( n6525 , n6524 , n5221 );
buf ( n6526 , n6525 );
xor ( n6527 , n6523 , n6526 );
xor ( n6528 , n6520 , n6527 );
xor ( n6529 , n4749 , n4751 );
xor ( n6530 , n6529 , n5218 );
buf ( n6531 , n6530 );
xor ( n6532 , n4753 , n4755 );
xor ( n6533 , n6532 , n5215 );
buf ( n6534 , n6533 );
xor ( n6535 , n6531 , n6534 );
xor ( n6536 , n4757 , n4759 );
xor ( n6537 , n6536 , n5212 );
buf ( n6538 , n6537 );
xor ( n6539 , n4761 , n4763 );
xor ( n6540 , n6539 , n5209 );
buf ( n6541 , n6540 );
xor ( n6542 , n6538 , n6541 );
xor ( n6543 , n6535 , n6542 );
xor ( n6544 , n6528 , n6543 );
xor ( n6545 , n6513 , n6544 );
xor ( n6546 , n6482 , n6545 );
xor ( n6547 , n6419 , n6546 );
xor ( n6548 , n4765 , n4767 );
xor ( n6549 , n6548 , n5206 );
buf ( n6550 , n6549 );
xor ( n6551 , n4769 , n4771 );
xor ( n6552 , n6551 , n5203 );
buf ( n6553 , n6552 );
xor ( n6554 , n6550 , n6553 );
xor ( n6555 , n4773 , n4775 );
xor ( n6556 , n6555 , n5200 );
buf ( n6557 , n6556 );
xor ( n6558 , n4777 , n4779 );
xor ( n6559 , n6558 , n5197 );
buf ( n6560 , n6559 );
xor ( n6561 , n6557 , n6560 );
xor ( n6562 , n6554 , n6561 );
xor ( n6563 , n4781 , n4783 );
xor ( n6564 , n6563 , n5194 );
buf ( n6565 , n6564 );
xor ( n6566 , n4785 , n4787 );
xor ( n6567 , n6566 , n5191 );
buf ( n6568 , n6567 );
xor ( n6569 , n6565 , n6568 );
xor ( n6570 , n4789 , n4791 );
xor ( n6571 , n6570 , n5188 );
buf ( n6572 , n6571 );
xor ( n6573 , n4793 , n4795 );
xor ( n6574 , n6573 , n5185 );
buf ( n6575 , n6574 );
xor ( n6576 , n6572 , n6575 );
xor ( n6577 , n6569 , n6576 );
xor ( n6578 , n6562 , n6577 );
xor ( n6579 , n4797 , n4799 );
xor ( n6580 , n6579 , n5182 );
buf ( n6581 , n6580 );
xor ( n6582 , n4801 , n4803 );
xor ( n6583 , n6582 , n5179 );
buf ( n6584 , n6583 );
xor ( n6585 , n6581 , n6584 );
xor ( n6586 , n4805 , n4807 );
xor ( n6587 , n6586 , n5176 );
buf ( n6588 , n6587 );
xor ( n6589 , n4809 , n4811 );
xor ( n6590 , n6589 , n5173 );
buf ( n6591 , n6590 );
xor ( n6592 , n6588 , n6591 );
xor ( n6593 , n6585 , n6592 );
xor ( n6594 , n4813 , n4815 );
xor ( n6595 , n6594 , n5170 );
buf ( n6596 , n6595 );
xor ( n6597 , n4817 , n4819 );
xor ( n6598 , n6597 , n5167 );
buf ( n6599 , n6598 );
xor ( n6600 , n6596 , n6599 );
xor ( n6601 , n4821 , n4823 );
xor ( n6602 , n6601 , n5164 );
buf ( n6603 , n6602 );
xor ( n6604 , n4825 , n4827 );
xor ( n6605 , n6604 , n5161 );
buf ( n6606 , n6605 );
xor ( n6607 , n6603 , n6606 );
xor ( n6608 , n6600 , n6607 );
xor ( n6609 , n6593 , n6608 );
xor ( n6610 , n6578 , n6609 );
xor ( n6611 , n4829 , n4831 );
xor ( n6612 , n6611 , n5158 );
buf ( n6613 , n6612 );
xor ( n6614 , n4833 , n4835 );
xor ( n6615 , n6614 , n5155 );
buf ( n6616 , n6615 );
xor ( n6617 , n6613 , n6616 );
xor ( n6618 , n4837 , n4839 );
xor ( n6619 , n6618 , n5152 );
buf ( n6620 , n6619 );
xor ( n6621 , n4841 , n4843 );
xor ( n6622 , n6621 , n5149 );
buf ( n6623 , n6622 );
xor ( n6624 , n6620 , n6623 );
xor ( n6625 , n6617 , n6624 );
xor ( n6626 , n4845 , n4847 );
xor ( n6627 , n6626 , n5146 );
buf ( n6628 , n6627 );
xor ( n6629 , n4849 , n4851 );
xor ( n6630 , n6629 , n5143 );
buf ( n6631 , n6630 );
xor ( n6632 , n6628 , n6631 );
xor ( n6633 , n4853 , n4855 );
xor ( n6634 , n6633 , n5140 );
buf ( n6635 , n6634 );
xor ( n6636 , n4857 , n4859 );
xor ( n6637 , n6636 , n5137 );
buf ( n6638 , n6637 );
xor ( n6639 , n6635 , n6638 );
xor ( n6640 , n6632 , n6639 );
xor ( n6641 , n6625 , n6640 );
xor ( n6642 , n4861 , n4863 );
xor ( n6643 , n6642 , n5134 );
buf ( n6644 , n6643 );
xor ( n6645 , n4865 , n4867 );
xor ( n6646 , n6645 , n5131 );
buf ( n6647 , n6646 );
xor ( n6648 , n6644 , n6647 );
xor ( n6649 , n4869 , n4871 );
xor ( n6650 , n6649 , n5128 );
buf ( n6651 , n6650 );
xor ( n6652 , n4873 , n4875 );
xor ( n6653 , n6652 , n5125 );
buf ( n6654 , n6653 );
xor ( n6655 , n6651 , n6654 );
xor ( n6656 , n6648 , n6655 );
xor ( n6657 , n4877 , n4879 );
xor ( n6658 , n6657 , n5122 );
buf ( n6659 , n6658 );
xor ( n6660 , n4881 , n4883 );
xor ( n6661 , n6660 , n5119 );
buf ( n6662 , n6661 );
xor ( n6663 , n6659 , n6662 );
xor ( n6664 , n4885 , n4887 );
xor ( n6665 , n6664 , n5116 );
buf ( n6666 , n6665 );
xor ( n6667 , n4889 , n4891 );
xor ( n6668 , n6667 , n5113 );
buf ( n6669 , n6668 );
xor ( n6670 , n6666 , n6669 );
xor ( n6671 , n6663 , n6670 );
xor ( n6672 , n6656 , n6671 );
xor ( n6673 , n6641 , n6672 );
xor ( n6674 , n6610 , n6673 );
xor ( n6675 , n4893 , n4895 );
xor ( n6676 , n6675 , n5110 );
buf ( n6677 , n6676 );
xor ( n6678 , n4897 , n4899 );
xor ( n6679 , n6678 , n5107 );
buf ( n6680 , n6679 );
xor ( n6681 , n6677 , n6680 );
xor ( n6682 , n4901 , n4903 );
xor ( n6683 , n6682 , n5104 );
buf ( n6684 , n6683 );
xor ( n6685 , n4905 , n4907 );
xor ( n6686 , n6685 , n5101 );
buf ( n6687 , n6686 );
xor ( n6688 , n6684 , n6687 );
xor ( n6689 , n6681 , n6688 );
xor ( n6690 , n4909 , n4911 );
xor ( n6691 , n6690 , n5098 );
buf ( n6692 , n6691 );
xor ( n6693 , n4913 , n4915 );
xor ( n6694 , n6693 , n5095 );
buf ( n6695 , n6694 );
xor ( n6696 , n6692 , n6695 );
xor ( n6697 , n4917 , n4919 );
xor ( n6698 , n6697 , n5092 );
buf ( n6699 , n6698 );
xor ( n6700 , n4921 , n4923 );
xor ( n6701 , n6700 , n5089 );
buf ( n6702 , n6701 );
xor ( n6703 , n6699 , n6702 );
xor ( n6704 , n6696 , n6703 );
xor ( n6705 , n6689 , n6704 );
xor ( n6706 , n4925 , n4927 );
xor ( n6707 , n6706 , n5086 );
buf ( n6708 , n6707 );
xor ( n6709 , n4929 , n4931 );
xor ( n6710 , n6709 , n5083 );
buf ( n6711 , n6710 );
xor ( n6712 , n6708 , n6711 );
xor ( n6713 , n4933 , n4935 );
xor ( n6714 , n6713 , n5080 );
buf ( n6715 , n6714 );
xor ( n6716 , n4937 , n4939 );
xor ( n6717 , n6716 , n5077 );
buf ( n6718 , n6717 );
xor ( n6719 , n6715 , n6718 );
xor ( n6720 , n6712 , n6719 );
xor ( n6721 , n4941 , n4943 );
xor ( n6722 , n6721 , n5074 );
buf ( n6723 , n6722 );
xor ( n6724 , n4945 , n4947 );
xor ( n6725 , n6724 , n5071 );
buf ( n6726 , n6725 );
xor ( n6727 , n6723 , n6726 );
xor ( n6728 , n4949 , n4951 );
xor ( n6729 , n6728 , n5068 );
buf ( n6730 , n6729 );
xor ( n6731 , n4953 , n4955 );
xor ( n6732 , n6731 , n5065 );
buf ( n6733 , n6732 );
xor ( n6734 , n6730 , n6733 );
xor ( n6735 , n6727 , n6734 );
xor ( n6736 , n6720 , n6735 );
xor ( n6737 , n6705 , n6736 );
xor ( n6738 , n4957 , n4959 );
xor ( n6739 , n6738 , n5062 );
buf ( n6740 , n6739 );
xor ( n6741 , n4961 , n4963 );
xor ( n6742 , n6741 , n5059 );
buf ( n6743 , n6742 );
xor ( n6744 , n6740 , n6743 );
xor ( n6745 , n4965 , n4967 );
xor ( n6746 , n6745 , n5056 );
buf ( n6747 , n6746 );
xor ( n6748 , n4969 , n4971 );
xor ( n6749 , n6748 , n5053 );
buf ( n6750 , n6749 );
xor ( n6751 , n6747 , n6750 );
xor ( n6752 , n6744 , n6751 );
xor ( n6753 , n4973 , n4975 );
xor ( n6754 , n6753 , n5050 );
buf ( n6755 , n6754 );
xor ( n6756 , n4977 , n4979 );
xor ( n6757 , n6756 , n5047 );
buf ( n6758 , n6757 );
xor ( n6759 , n6755 , n6758 );
xor ( n6760 , n4981 , n4983 );
xor ( n6761 , n6760 , n5044 );
buf ( n6762 , n6761 );
xor ( n6763 , n4985 , n4987 );
xor ( n6764 , n6763 , n5041 );
buf ( n6765 , n6764 );
xor ( n6766 , n6762 , n6765 );
xor ( n6767 , n6759 , n6766 );
xor ( n6768 , n6752 , n6767 );
xor ( n6769 , n4989 , n4991 );
xor ( n6770 , n6769 , n5038 );
buf ( n6771 , n6770 );
xor ( n6772 , n4993 , n4995 );
xor ( n6773 , n6772 , n5035 );
buf ( n6774 , n6773 );
xor ( n6775 , n6771 , n6774 );
xor ( n6776 , n4997 , n4999 );
xor ( n6777 , n6776 , n5032 );
buf ( n6778 , n6777 );
xor ( n6779 , n5001 , n5003 );
xor ( n6780 , n6779 , n5029 );
buf ( n6781 , n6780 );
xor ( n6782 , n6778 , n6781 );
xor ( n6783 , n6775 , n6782 );
xor ( n6784 , n5005 , n5007 );
xor ( n6785 , n6784 , n5026 );
buf ( n6786 , n6785 );
xor ( n6787 , n5009 , n5011 );
xor ( n6788 , n6787 , n5023 );
buf ( n6789 , n6788 );
xor ( n6790 , n6786 , n6789 );
xor ( n6791 , n5013 , n5015 );
xor ( n6792 , n6791 , n5020 );
buf ( n6793 , n6792 );
xor ( n6794 , n5017 , n5018 );
buf ( n6795 , n6794 );
xor ( n6796 , n6793 , n6795 );
xor ( n6797 , n6790 , n6796 );
xor ( n6798 , n6783 , n6797 );
xor ( n6799 , n6768 , n6798 );
xor ( n6800 , n6737 , n6799 );
xor ( n6801 , n6674 , n6800 );
xor ( n6802 , n6547 , n6801 );
xor ( n6803 , n6292 , n6802 );
buf ( n6804 , n6803 );
buf ( n6805 , n6804 );
endmodule

