//
// Conformal-LEC Version 15.20-d227 ( 10-Mar-2016) ( 64 bit executable)
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
output n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 ;

wire n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , 
     n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , 
     n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , 
     n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , 
     n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
     n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
     n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , 
     n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , 
     n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , 
     n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , 
     n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , 
     n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , 
     n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , 
     n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , 
     n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , 
     n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , 
     n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , 
     n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , 
     n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
     n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
     n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
     n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
     n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , 
     n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , 
     n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , 
     n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , 
     n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , 
     n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , 
     n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , 
     n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , 
     n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , 
     n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , 
     n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , 
     n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , 
     n457 , n458 ;
buf ( n47 , n402 );
buf ( n51 , n405 );
buf ( n55 , n408 );
buf ( n49 , n412 );
buf ( n50 , n416 );
buf ( n52 , n420 );
buf ( n46 , n424 );
buf ( n53 , n428 );
buf ( n48 , n432 );
buf ( n57 , n436 );
buf ( n45 , n440 );
buf ( n58 , n444 );
buf ( n56 , n448 );
buf ( n44 , n452 );
buf ( n54 , n455 );
buf ( n43 , n458 );
buf ( n120 , n32 );
buf ( n121 , n27 );
buf ( n122 , n34 );
buf ( n123 , n9 );
buf ( n124 , n37 );
buf ( n125 , n13 );
buf ( n126 , n42 );
buf ( n127 , n12 );
buf ( n128 , n41 );
buf ( n129 , n33 );
buf ( n130 , n15 );
buf ( n131 , n38 );
buf ( n132 , n28 );
buf ( n133 , n1 );
buf ( n134 , n24 );
buf ( n135 , n2 );
buf ( n136 , n23 );
buf ( n137 , n4 );
buf ( n138 , n22 );
buf ( n139 , n11 );
buf ( n140 , n10 );
buf ( n141 , n29 );
buf ( n142 , n3 );
buf ( n143 , n18 );
buf ( n144 , n14 );
buf ( n145 , n36 );
buf ( n146 , n17 );
buf ( n147 , n30 );
buf ( n148 , n35 );
buf ( n149 , n0 );
buf ( n150 , n7 );
buf ( n151 , n31 );
buf ( n152 , n20 );
buf ( n153 , n8 );
buf ( n154 , n21 );
buf ( n155 , n39 );
buf ( n156 , n5 );
buf ( n157 , n19 );
buf ( n158 , n16 );
buf ( n159 , n6 );
buf ( n160 , n25 );
buf ( n161 , n40 );
buf ( n162 , n26 );
buf ( n163 , n120 );
buf ( n164 , n136 );
not ( n165 , n164 );
xor ( n166 , n163 , n165 );
buf ( n167 , n121 );
buf ( n168 , n137 );
not ( n169 , n168 );
and ( n170 , n167 , n169 );
buf ( n171 , n122 );
buf ( n172 , n138 );
not ( n173 , n172 );
and ( n174 , n171 , n173 );
buf ( n175 , n123 );
buf ( n176 , n139 );
not ( n177 , n176 );
and ( n178 , n175 , n177 );
buf ( n179 , n124 );
buf ( n180 , n140 );
not ( n181 , n180 );
and ( n182 , n179 , n181 );
buf ( n183 , n125 );
buf ( n184 , n141 );
not ( n185 , n184 );
and ( n186 , n183 , n185 );
buf ( n187 , n126 );
buf ( n188 , n142 );
not ( n189 , n188 );
and ( n190 , n187 , n189 );
buf ( n191 , n127 );
buf ( n192 , n143 );
not ( n193 , n192 );
and ( n194 , n191 , n193 );
buf ( n195 , n128 );
buf ( n196 , n144 );
not ( n197 , n196 );
and ( n198 , n195 , n197 );
buf ( n199 , n129 );
buf ( n200 , n145 );
not ( n201 , n200 );
and ( n202 , n199 , n201 );
buf ( n203 , n130 );
buf ( n204 , n146 );
not ( n205 , n204 );
and ( n206 , n203 , n205 );
buf ( n207 , n131 );
buf ( n208 , n147 );
not ( n209 , n208 );
and ( n210 , n207 , n209 );
buf ( n211 , n132 );
buf ( n212 , n148 );
not ( n213 , n212 );
and ( n214 , n211 , n213 );
buf ( n215 , n133 );
buf ( n216 , n149 );
not ( n217 , n216 );
and ( n218 , n215 , n217 );
buf ( n219 , n134 );
buf ( n220 , n150 );
not ( n221 , n220 );
and ( n222 , n219 , n221 );
buf ( n223 , n135 );
buf ( n224 , n151 );
not ( n225 , n224 );
or ( n226 , n223 , n225 );
and ( n227 , n221 , n226 );
and ( n228 , n219 , n226 );
or ( n229 , n222 , n227 , n228 );
and ( n230 , n217 , n229 );
and ( n231 , n215 , n229 );
or ( n232 , n218 , n230 , n231 );
and ( n233 , n213 , n232 );
and ( n234 , n211 , n232 );
or ( n235 , n214 , n233 , n234 );
and ( n236 , n209 , n235 );
and ( n237 , n207 , n235 );
or ( n238 , n210 , n236 , n237 );
and ( n239 , n205 , n238 );
and ( n240 , n203 , n238 );
or ( n241 , n206 , n239 , n240 );
and ( n242 , n201 , n241 );
and ( n243 , n199 , n241 );
or ( n244 , n202 , n242 , n243 );
and ( n245 , n197 , n244 );
and ( n246 , n195 , n244 );
or ( n247 , n198 , n245 , n246 );
and ( n248 , n193 , n247 );
and ( n249 , n191 , n247 );
or ( n250 , n194 , n248 , n249 );
and ( n251 , n189 , n250 );
and ( n252 , n187 , n250 );
or ( n253 , n190 , n251 , n252 );
and ( n254 , n185 , n253 );
and ( n255 , n183 , n253 );
or ( n256 , n186 , n254 , n255 );
and ( n257 , n181 , n256 );
and ( n258 , n179 , n256 );
or ( n259 , n182 , n257 , n258 );
and ( n260 , n177 , n259 );
and ( n261 , n175 , n259 );
or ( n262 , n178 , n260 , n261 );
and ( n263 , n173 , n262 );
and ( n264 , n171 , n262 );
or ( n265 , n174 , n263 , n264 );
and ( n266 , n169 , n265 );
and ( n267 , n167 , n265 );
or ( n268 , n170 , n266 , n267 );
xor ( n269 , n166 , n268 );
buf ( n270 , n269 );
buf ( n271 , n270 );
xor ( n272 , n167 , n169 );
xor ( n273 , n272 , n265 );
buf ( n274 , n273 );
buf ( n275 , n274 );
xor ( n276 , n171 , n173 );
xor ( n277 , n276 , n262 );
buf ( n278 , n277 );
buf ( n279 , n278 );
xor ( n280 , n175 , n177 );
xor ( n281 , n280 , n259 );
buf ( n282 , n281 );
buf ( n283 , n282 );
not ( n284 , n152 );
buf ( n285 , n284 );
and ( n286 , n283 , n285 );
xor ( n287 , n179 , n181 );
xor ( n288 , n287 , n256 );
buf ( n289 , n288 );
buf ( n290 , n289 );
not ( n291 , n153 );
buf ( n292 , n291 );
and ( n293 , n290 , n292 );
xor ( n294 , n183 , n185 );
xor ( n295 , n294 , n253 );
buf ( n296 , n295 );
buf ( n297 , n296 );
not ( n298 , n154 );
buf ( n299 , n298 );
and ( n300 , n297 , n299 );
xor ( n301 , n187 , n189 );
xor ( n302 , n301 , n250 );
buf ( n303 , n302 );
buf ( n304 , n303 );
not ( n305 , n155 );
buf ( n306 , n305 );
and ( n307 , n304 , n306 );
xor ( n308 , n191 , n193 );
xor ( n309 , n308 , n247 );
buf ( n310 , n309 );
buf ( n311 , n310 );
not ( n312 , n156 );
buf ( n313 , n312 );
and ( n314 , n311 , n313 );
xor ( n315 , n195 , n197 );
xor ( n316 , n315 , n244 );
buf ( n317 , n316 );
buf ( n318 , n317 );
not ( n319 , n157 );
buf ( n320 , n319 );
and ( n321 , n318 , n320 );
xor ( n322 , n199 , n201 );
xor ( n323 , n322 , n241 );
buf ( n324 , n323 );
buf ( n325 , n324 );
not ( n326 , n158 );
buf ( n327 , n326 );
and ( n328 , n325 , n327 );
xor ( n329 , n203 , n205 );
xor ( n330 , n329 , n238 );
buf ( n331 , n330 );
buf ( n332 , n331 );
not ( n333 , n159 );
buf ( n334 , n333 );
and ( n335 , n332 , n334 );
xor ( n336 , n207 , n209 );
xor ( n337 , n336 , n235 );
buf ( n338 , n337 );
buf ( n339 , n338 );
not ( n340 , n160 );
buf ( n341 , n340 );
and ( n342 , n339 , n341 );
xor ( n343 , n211 , n213 );
xor ( n344 , n343 , n232 );
buf ( n345 , n344 );
buf ( n346 , n345 );
not ( n347 , n161 );
buf ( n348 , n347 );
and ( n349 , n346 , n348 );
xor ( n350 , n215 , n217 );
xor ( n351 , n350 , n229 );
buf ( n352 , n351 );
buf ( n353 , n352 );
not ( n354 , n162 );
buf ( n355 , n354 );
and ( n356 , n353 , n355 );
xor ( n357 , n219 , n221 );
xor ( n358 , n357 , n226 );
buf ( n359 , n358 );
buf ( n360 , n359 );
xor ( n361 , n223 , n224 );
buf ( n362 , n361 );
buf ( n363 , n362 );
or ( n364 , n360 , n363 );
and ( n365 , n355 , n364 );
and ( n366 , n353 , n364 );
or ( n367 , n356 , n365 , n366 );
and ( n368 , n348 , n367 );
and ( n369 , n346 , n367 );
or ( n370 , n349 , n368 , n369 );
and ( n371 , n341 , n370 );
and ( n372 , n339 , n370 );
or ( n373 , n342 , n371 , n372 );
and ( n374 , n334 , n373 );
and ( n375 , n332 , n373 );
or ( n376 , n335 , n374 , n375 );
and ( n377 , n327 , n376 );
and ( n378 , n325 , n376 );
or ( n379 , n328 , n377 , n378 );
and ( n380 , n320 , n379 );
and ( n381 , n318 , n379 );
or ( n382 , n321 , n380 , n381 );
and ( n383 , n313 , n382 );
and ( n384 , n311 , n382 );
or ( n385 , n314 , n383 , n384 );
and ( n386 , n306 , n385 );
and ( n387 , n304 , n385 );
or ( n388 , n307 , n386 , n387 );
and ( n389 , n299 , n388 );
and ( n390 , n297 , n388 );
or ( n391 , n300 , n389 , n390 );
and ( n392 , n292 , n391 );
and ( n393 , n290 , n391 );
or ( n394 , n293 , n392 , n393 );
and ( n395 , n285 , n394 );
and ( n396 , n283 , n394 );
or ( n397 , n286 , n395 , n396 );
and ( n398 , n279 , n397 );
and ( n399 , n275 , n398 );
xor ( n400 , n271 , n399 );
buf ( n401 , n400 );
buf ( n402 , n401 );
xor ( n403 , n275 , n398 );
buf ( n404 , n403 );
buf ( n405 , n404 );
xor ( n406 , n279 , n397 );
buf ( n407 , n406 );
buf ( n408 , n407 );
xor ( n409 , n283 , n285 );
xor ( n410 , n409 , n394 );
buf ( n411 , n410 );
buf ( n412 , n411 );
xor ( n413 , n290 , n292 );
xor ( n414 , n413 , n391 );
buf ( n415 , n414 );
buf ( n416 , n415 );
xor ( n417 , n297 , n299 );
xor ( n418 , n417 , n388 );
buf ( n419 , n418 );
buf ( n420 , n419 );
xor ( n421 , n304 , n306 );
xor ( n422 , n421 , n385 );
buf ( n423 , n422 );
buf ( n424 , n423 );
xor ( n425 , n311 , n313 );
xor ( n426 , n425 , n382 );
buf ( n427 , n426 );
buf ( n428 , n427 );
xor ( n429 , n318 , n320 );
xor ( n430 , n429 , n379 );
buf ( n431 , n430 );
buf ( n432 , n431 );
xor ( n433 , n325 , n327 );
xor ( n434 , n433 , n376 );
buf ( n435 , n434 );
buf ( n436 , n435 );
xor ( n437 , n332 , n334 );
xor ( n438 , n437 , n373 );
buf ( n439 , n438 );
buf ( n440 , n439 );
xor ( n441 , n339 , n341 );
xor ( n442 , n441 , n370 );
buf ( n443 , n442 );
buf ( n444 , n443 );
xor ( n445 , n346 , n348 );
xor ( n446 , n445 , n367 );
buf ( n447 , n446 );
buf ( n448 , n447 );
xor ( n449 , n353 , n355 );
xor ( n450 , n449 , n364 );
buf ( n451 , n450 );
buf ( n452 , n451 );
xnor ( n453 , n360 , n363 );
buf ( n454 , n453 );
buf ( n455 , n454 );
not ( n456 , n363 );
buf ( n457 , n456 );
buf ( n458 , n457 );
endmodule

