//
// Conformal-LEC Version 16.10-d005 ( 21-Apr-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 ;
output n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 ;

wire n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , 
     n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , 
     n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , 
     n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , 
     n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , 
     n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , 
     n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , 
     n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , 
     n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , 
     n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , 
     n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , 
     n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , 
     n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , 
     n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , 
     n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , 
     n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , 
     n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
     n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , 
     n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , 
     n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , 
     n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
     n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , 
     n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , 
     n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , 
     n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , 
     n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , 
     n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , 
     n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , 
     n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , 
     n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , 
     n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , 
     n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , 
     n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , 
     n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , 
     n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , 
     n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , 
     n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , 
     n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , 
     n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , 
     n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , 
     n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , 
     n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , 
     n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , 
     n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , 
     n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , 
     n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , 
     n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , 
     n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , 
     n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , 
     n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , 
     n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , 
     n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , 
     n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , 
     n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , 
     n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , 
     n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , 
     n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , 
     n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , 
     n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , 
     n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , 
     n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , 
     n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , 
     n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , 
     n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , 
     n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , 
     n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , 
     n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , 
     n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , 
     n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , 
     n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , 
     n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , 
     n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , 
     n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , 
     n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , 
     n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , 
     n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , 
     n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , 
     n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , 
     n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , 
     n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , 
     n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , 
     n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , 
     n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , 
     n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , 
     n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , 
     n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , 
     n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , 
     n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , 
     n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , 
     n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , 
     n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , 
     n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , 
     n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , 
     n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , 
     n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , 
     n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , 
     n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , 
     n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , 
     n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , 
     n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , 
     n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , 
     n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , 
     n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , 
     n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , 
     n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , 
     n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , 
     n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , 
     n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , 
     n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , 
     n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , 
     n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , 
     n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , 
     n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , 
     n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , 
     n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , 
     n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , 
     n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , 
     n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , 
     n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , 
     n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , 
     n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , 
     n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , 
     n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , 
     n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , 
     n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , 
     n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , 
     n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , 
     n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , 
     n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , 
     n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , 
     n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , 
     n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , 
     n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , 
     n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , 
     n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , 
     n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , 
     n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , 
     n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , 
     n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , 
     n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , 
     n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , 
     n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , 
     n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , 
     n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , 
     n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , 
     n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , 
     n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , 
     n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , 
     n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , 
     n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , 
     n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , 
     n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , 
     n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , 
     n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , 
     n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , 
     n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , 
     n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , 
     n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , 
     n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , 
     n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , 
     n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , 
     n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , 
     n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , 
     n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , 
     n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , 
     n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , 
     n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , 
     n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , 
     n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , 
     n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , 
     n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , 
     n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , 
     n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , 
     n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , 
     n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , 
     n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , 
     n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , 
     n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , 
     n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , 
     n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , 
     n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , 
     n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , 
     n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , 
     n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , 
     n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , 
     n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , 
     n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , 
     n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , 
     n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , 
     n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , 
     n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , 
     n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , 
     n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , 
     n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , 
     n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , 
     n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , 
     n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , 
     n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , 
     n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , 
     n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , 
     n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , 
     n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , 
     n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , 
     n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , 
     n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , 
     n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , 
     n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , 
     n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , 
     n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , 
     n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , 
     n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , 
     n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , 
     n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , 
     n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , 
     n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , 
     n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , 
     n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , 
     n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , 
     n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , 
     n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , 
     n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , 
     n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , 
     n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , 
     n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , 
     n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , 
     n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , 
     n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , 
     n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , 
     n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , 
     n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , 
     n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , 
     n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , 
     n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , 
     n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , 
     n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , 
     n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , 
     n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , 
     n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , 
     n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , 
     n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , 
     n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , 
     n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , 
     n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , 
     n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , 
     n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , 
     n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , 
     n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , 
     n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , 
     n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , 
     n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , 
     n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , 
     n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , 
     n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , 
     n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , 
     n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , 
     n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , 
     n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , 
     n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , 
     n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , 
     n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , 
     n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , 
     n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , 
     n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , 
     n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , 
     n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , 
     n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , 
     n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , 
     n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , 
     n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , 
     n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , 
     n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , 
     n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , 
     n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , 
     n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , 
     n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , 
     n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , 
     n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , 
     n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , 
     n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , 
     n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , 
     n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , 
     n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , 
     n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , 
     n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , 
     n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , 
     n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , 
     n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , 
     n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , 
     n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , 
     n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , 
     n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , 
     n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , 
     n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , 
     n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , 
     n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , 
     n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , 
     n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , 
     n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , 
     n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , 
     n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , 
     n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , 
     n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , 
     n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , 
     n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , 
     n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , 
     n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , 
     n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , 
     n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , 
     n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , 
     n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , 
     n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , 
     n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , 
     n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , 
     n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , 
     n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , 
     n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , 
     n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , 
     n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , 
     n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , 
     n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , 
     n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , 
     n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , 
     n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , 
     n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , 
     n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , 
     n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , 
     n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , 
     n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , 
     n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , 
     n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , 
     n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , 
     n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , 
     n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , 
     n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , 
     n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , 
     n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , 
     n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , 
     n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , 
     n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , 
     n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , 
     n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , 
     n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , 
     n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , 
     n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , 
     n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , 
     n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , 
     n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , 
     n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , 
     n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , 
     n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , 
     n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , 
     n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , 
     n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , 
     n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , 
     n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , 
     n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , 
     n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , 
     n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , 
     n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , 
     n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , 
     n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , 
     n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , 
     n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , 
     n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , 
     n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , 
     n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , 
     n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , 
     n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , 
     n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , 
     n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , 
     n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , 
     n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , 
     n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 ;
buf ( n197 , n3489 );
buf ( n194 , n3648 );
buf ( n202 , n3705 );
buf ( n195 , n3762 );
buf ( n199 , n3836 );
buf ( n200 , n3897 );
buf ( n201 , n3956 );
buf ( n193 , n4014 );
buf ( n196 , n4072 );
buf ( n198 , n4133 );
buf ( n530 , n104 );
buf ( n531 , n55 );
buf ( n532 , n113 );
buf ( n533 , n145 );
buf ( n534 , n78 );
buf ( n535 , n156 );
buf ( n536 , n191 );
buf ( n537 , n167 );
buf ( n538 , n76 );
buf ( n539 , n107 );
buf ( n540 , n188 );
buf ( n541 , n4 );
buf ( n542 , n27 );
buf ( n543 , n114 );
buf ( n544 , n98 );
buf ( n545 , n95 );
buf ( n546 , n41 );
buf ( n547 , n39 );
buf ( n548 , n152 );
buf ( n549 , n142 );
buf ( n550 , n149 );
buf ( n551 , n179 );
buf ( n552 , n115 );
buf ( n553 , n16 );
buf ( n554 , n155 );
buf ( n555 , n65 );
buf ( n556 , n21 );
buf ( n557 , n86 );
buf ( n558 , n182 );
buf ( n559 , n133 );
buf ( n560 , n157 );
buf ( n561 , n34 );
buf ( n562 , n3 );
buf ( n563 , n105 );
buf ( n564 , n144 );
buf ( n565 , n136 );
buf ( n566 , n14 );
buf ( n567 , n19 );
buf ( n568 , n186 );
buf ( n569 , n54 );
buf ( n570 , n103 );
buf ( n571 , n40 );
buf ( n572 , n141 );
buf ( n573 , n45 );
buf ( n574 , n59 );
buf ( n575 , n46 );
buf ( n576 , n99 );
buf ( n577 , n172 );
buf ( n578 , n69 );
buf ( n579 , n80 );
buf ( n580 , n117 );
buf ( n581 , n2 );
buf ( n582 , n168 );
buf ( n583 , n66 );
buf ( n584 , n92 );
buf ( n585 , n57 );
buf ( n586 , n29 );
buf ( n587 , n79 );
buf ( n588 , n100 );
buf ( n589 , n44 );
buf ( n590 , n154 );
buf ( n591 , n36 );
buf ( n592 , n124 );
buf ( n593 , n120 );
buf ( n594 , n52 );
buf ( n595 , n161 );
buf ( n596 , n68 );
buf ( n597 , n9 );
buf ( n598 , n94 );
buf ( n599 , n175 );
buf ( n600 , n162 );
buf ( n601 , n164 );
buf ( n602 , n5 );
buf ( n603 , n138 );
buf ( n604 , n166 );
buf ( n605 , n181 );
buf ( n606 , n8 );
buf ( n607 , n83 );
buf ( n608 , n75 );
buf ( n609 , n72 );
buf ( n610 , n171 );
buf ( n611 , n170 );
buf ( n612 , n119 );
buf ( n613 , n189 );
buf ( n614 , n118 );
buf ( n615 , n108 );
buf ( n616 , n151 );
buf ( n617 , n126 );
buf ( n618 , n106 );
buf ( n619 , n70 );
buf ( n620 , n146 );
buf ( n621 , n50 );
buf ( n622 , n10 );
buf ( n623 , n89 );
buf ( n624 , n48 );
buf ( n625 , n178 );
buf ( n626 , n143 );
buf ( n627 , n180 );
buf ( n628 , n38 );
buf ( n629 , n122 );
buf ( n630 , n22 );
buf ( n631 , n169 );
buf ( n632 , n43 );
buf ( n633 , n96 );
buf ( n634 , n102 );
buf ( n635 , n91 );
buf ( n636 , n33 );
buf ( n637 , n42 );
buf ( n638 , n123 );
buf ( n639 , n12 );
buf ( n640 , n24 );
buf ( n641 , n163 );
buf ( n642 , n184 );
buf ( n643 , n15 );
buf ( n644 , n147 );
buf ( n645 , n121 );
buf ( n646 , n23 );
buf ( n647 , n63 );
buf ( n648 , n110 );
buf ( n649 , n185 );
buf ( n650 , n187 );
buf ( n651 , n25 );
buf ( n652 , n93 );
buf ( n653 , n7 );
buf ( n654 , n51 );
buf ( n655 , n165 );
buf ( n656 , n190 );
buf ( n657 , n132 );
buf ( n658 , n74 );
buf ( n659 , n160 );
buf ( n660 , n109 );
buf ( n661 , n20 );
buf ( n662 , n64 );
buf ( n663 , n53 );
buf ( n664 , n130 );
buf ( n665 , n11 );
buf ( n666 , n153 );
buf ( n667 , n127 );
buf ( n668 , n31 );
buf ( n669 , n97 );
buf ( n670 , n37 );
buf ( n671 , n0 );
buf ( n672 , n116 );
buf ( n673 , n134 );
buf ( n674 , n61 );
buf ( n675 , n148 );
buf ( n676 , n174 );
buf ( n677 , n137 );
buf ( n678 , n87 );
buf ( n679 , n131 );
buf ( n680 , n140 );
buf ( n681 , n158 );
buf ( n682 , n60 );
buf ( n683 , n85 );
buf ( n684 , n81 );
buf ( n685 , n150 );
buf ( n686 , n71 );
buf ( n687 , n177 );
buf ( n688 , n183 );
buf ( n689 , n84 );
buf ( n690 , n47 );
buf ( n691 , n159 );
buf ( n692 , n17 );
buf ( n693 , n82 );
buf ( n694 , n67 );
buf ( n695 , n139 );
buf ( n696 , n35 );
buf ( n697 , n18 );
buf ( n698 , n173 );
buf ( n699 , n77 );
buf ( n700 , n90 );
buf ( n701 , n111 );
buf ( n702 , n192 );
buf ( n703 , n125 );
buf ( n704 , n30 );
buf ( n705 , n28 );
buf ( n706 , n88 );
buf ( n707 , n13 );
buf ( n708 , n1 );
buf ( n709 , n62 );
buf ( n710 , n135 );
buf ( n711 , n128 );
buf ( n712 , n32 );
buf ( n713 , n58 );
buf ( n714 , n49 );
buf ( n715 , n73 );
buf ( n716 , n6 );
buf ( n717 , n129 );
buf ( n718 , n56 );
buf ( n719 , n26 );
buf ( n720 , n176 );
buf ( n721 , n112 );
not ( n722 , n530 );
not ( n723 , n531 );
not ( n724 , n532 );
not ( n725 , n533 );
not ( n726 , n534 );
not ( n727 , n535 );
not ( n728 , n536 );
not ( n729 , n537 );
not ( n730 , n538 );
not ( n731 , n540 );
not ( n732 , n541 );
not ( n733 , n542 );
not ( n734 , n543 );
not ( n735 , n544 );
not ( n736 , n545 );
not ( n737 , n546 );
not ( n738 , n547 );
not ( n739 , n548 );
not ( n740 , n549 );
not ( n741 , n550 );
not ( n742 , n551 );
not ( n743 , n552 );
not ( n744 , n553 );
not ( n745 , n554 );
not ( n746 , n555 );
not ( n747 , n556 );
not ( n748 , n557 );
not ( n749 , n558 );
not ( n750 , n559 );
not ( n751 , n560 );
not ( n752 , n561 );
and ( n753 , n751 , n752 );
and ( n754 , n750 , n753 );
and ( n755 , n749 , n754 );
and ( n756 , n748 , n755 );
and ( n757 , n747 , n756 );
and ( n758 , n746 , n757 );
and ( n759 , n745 , n758 );
and ( n760 , n744 , n759 );
and ( n761 , n743 , n760 );
and ( n762 , n742 , n761 );
and ( n763 , n741 , n762 );
and ( n764 , n740 , n763 );
and ( n765 , n739 , n764 );
and ( n766 , n738 , n765 );
and ( n767 , n737 , n766 );
and ( n768 , n736 , n767 );
and ( n769 , n735 , n768 );
and ( n770 , n734 , n769 );
and ( n771 , n733 , n770 );
and ( n772 , n732 , n771 );
and ( n773 , n731 , n772 );
buf ( n774 , n773 );
and ( n775 , n730 , n774 );
and ( n776 , n729 , n775 );
and ( n777 , n728 , n776 );
and ( n778 , n727 , n777 );
and ( n779 , n726 , n778 );
and ( n780 , n725 , n779 );
and ( n781 , n724 , n780 );
and ( n782 , n723 , n781 );
xor ( n783 , n722 , n782 );
and ( n784 , n783 , n530 );
not ( n785 , n784 );
and ( n786 , n722 , n538 );
xor ( n787 , n730 , n774 );
and ( n788 , n787 , n530 );
or ( n789 , n786 , n788 );
and ( n790 , n785 , n789 );
not ( n791 , n789 );
and ( n792 , n722 , n539 );
not ( n793 , n773 );
and ( n794 , n793 , n530 );
or ( n795 , n792 , n794 );
not ( n796 , n795 );
and ( n797 , n722 , n540 );
xor ( n798 , n731 , n772 );
and ( n799 , n798 , n530 );
or ( n800 , n797 , n799 );
not ( n801 , n800 );
and ( n802 , n722 , n541 );
xor ( n803 , n732 , n771 );
and ( n804 , n803 , n530 );
or ( n805 , n802 , n804 );
not ( n806 , n805 );
and ( n807 , n722 , n542 );
xor ( n808 , n733 , n770 );
and ( n809 , n808 , n530 );
or ( n810 , n807 , n809 );
not ( n811 , n810 );
and ( n812 , n722 , n543 );
xor ( n813 , n734 , n769 );
and ( n814 , n813 , n530 );
or ( n815 , n812 , n814 );
not ( n816 , n815 );
and ( n817 , n722 , n544 );
xor ( n818 , n735 , n768 );
and ( n819 , n818 , n530 );
or ( n820 , n817 , n819 );
not ( n821 , n820 );
and ( n822 , n722 , n545 );
xor ( n823 , n736 , n767 );
and ( n824 , n823 , n530 );
or ( n825 , n822 , n824 );
not ( n826 , n825 );
and ( n827 , n722 , n546 );
xor ( n828 , n737 , n766 );
and ( n829 , n828 , n530 );
or ( n830 , n827 , n829 );
not ( n831 , n830 );
and ( n832 , n722 , n547 );
xor ( n833 , n738 , n765 );
and ( n834 , n833 , n530 );
or ( n835 , n832 , n834 );
not ( n836 , n835 );
and ( n837 , n722 , n548 );
xor ( n838 , n739 , n764 );
and ( n839 , n838 , n530 );
or ( n840 , n837 , n839 );
not ( n841 , n840 );
and ( n842 , n722 , n549 );
xor ( n843 , n740 , n763 );
and ( n844 , n843 , n530 );
or ( n845 , n842 , n844 );
not ( n846 , n845 );
and ( n847 , n722 , n550 );
xor ( n848 , n741 , n762 );
and ( n849 , n848 , n530 );
or ( n850 , n847 , n849 );
not ( n851 , n850 );
and ( n852 , n722 , n551 );
xor ( n853 , n742 , n761 );
and ( n854 , n853 , n530 );
or ( n855 , n852 , n854 );
not ( n856 , n855 );
and ( n857 , n722 , n552 );
xor ( n858 , n743 , n760 );
and ( n859 , n858 , n530 );
or ( n860 , n857 , n859 );
not ( n861 , n860 );
and ( n862 , n722 , n553 );
xor ( n863 , n744 , n759 );
and ( n864 , n863 , n530 );
or ( n865 , n862 , n864 );
not ( n866 , n865 );
and ( n867 , n722 , n554 );
xor ( n868 , n745 , n758 );
and ( n869 , n868 , n530 );
or ( n870 , n867 , n869 );
not ( n871 , n870 );
and ( n872 , n722 , n555 );
xor ( n873 , n746 , n757 );
and ( n874 , n873 , n530 );
or ( n875 , n872 , n874 );
not ( n876 , n875 );
and ( n877 , n722 , n556 );
xor ( n878 , n747 , n756 );
and ( n879 , n878 , n530 );
or ( n880 , n877 , n879 );
not ( n881 , n880 );
and ( n882 , n722 , n557 );
xor ( n883 , n748 , n755 );
and ( n884 , n883 , n530 );
or ( n885 , n882 , n884 );
not ( n886 , n885 );
and ( n887 , n722 , n558 );
xor ( n888 , n749 , n754 );
and ( n889 , n888 , n530 );
or ( n890 , n887 , n889 );
not ( n891 , n890 );
and ( n892 , n722 , n559 );
xor ( n893 , n750 , n753 );
and ( n894 , n893 , n530 );
or ( n895 , n892 , n894 );
not ( n896 , n895 );
and ( n897 , n722 , n560 );
xor ( n898 , n751 , n752 );
and ( n899 , n898 , n530 );
or ( n900 , n897 , n899 );
not ( n901 , n900 );
and ( n902 , n901 , n752 );
and ( n903 , n896 , n902 );
and ( n904 , n891 , n903 );
and ( n905 , n886 , n904 );
and ( n906 , n881 , n905 );
and ( n907 , n876 , n906 );
and ( n908 , n871 , n907 );
and ( n909 , n866 , n908 );
and ( n910 , n861 , n909 );
and ( n911 , n856 , n910 );
and ( n912 , n851 , n911 );
and ( n913 , n846 , n912 );
and ( n914 , n841 , n913 );
and ( n915 , n836 , n914 );
and ( n916 , n831 , n915 );
and ( n917 , n826 , n916 );
and ( n918 , n821 , n917 );
and ( n919 , n816 , n918 );
and ( n920 , n811 , n919 );
and ( n921 , n806 , n920 );
and ( n922 , n801 , n921 );
and ( n923 , n796 , n922 );
xor ( n924 , n791 , n923 );
and ( n925 , n924 , n784 );
or ( n926 , n790 , n925 );
and ( n927 , n722 , n531 );
xor ( n928 , n723 , n781 );
and ( n929 , n928 , n530 );
or ( n930 , n927 , n929 );
not ( n931 , n930 );
and ( n932 , n722 , n532 );
xor ( n933 , n724 , n780 );
and ( n934 , n933 , n530 );
or ( n935 , n932 , n934 );
not ( n936 , n935 );
and ( n937 , n722 , n533 );
xor ( n938 , n725 , n779 );
and ( n939 , n938 , n530 );
or ( n940 , n937 , n939 );
not ( n941 , n940 );
and ( n942 , n722 , n534 );
xor ( n943 , n726 , n778 );
and ( n944 , n943 , n530 );
or ( n945 , n942 , n944 );
not ( n946 , n945 );
and ( n947 , n722 , n535 );
xor ( n948 , n727 , n777 );
and ( n949 , n948 , n530 );
or ( n950 , n947 , n949 );
not ( n951 , n950 );
and ( n952 , n722 , n536 );
xor ( n953 , n728 , n776 );
and ( n954 , n953 , n530 );
or ( n955 , n952 , n954 );
not ( n956 , n955 );
and ( n957 , n722 , n537 );
xor ( n958 , n729 , n775 );
and ( n959 , n958 , n530 );
or ( n960 , n957 , n959 );
not ( n961 , n960 );
and ( n962 , n791 , n923 );
and ( n963 , n961 , n962 );
and ( n964 , n956 , n963 );
and ( n965 , n951 , n964 );
and ( n966 , n946 , n965 );
and ( n967 , n941 , n966 );
and ( n968 , n936 , n967 );
and ( n969 , n931 , n968 );
xor ( n970 , n785 , n969 );
and ( n971 , n970 , n784 );
not ( n972 , n971 );
and ( n973 , n785 , n930 );
xor ( n974 , n931 , n968 );
and ( n975 , n974 , n784 );
or ( n976 , n973 , n975 );
not ( n977 , n976 );
and ( n978 , n785 , n935 );
xor ( n979 , n936 , n967 );
and ( n980 , n979 , n784 );
or ( n981 , n978 , n980 );
not ( n982 , n981 );
and ( n983 , n785 , n940 );
xor ( n984 , n941 , n966 );
and ( n985 , n984 , n784 );
or ( n986 , n983 , n985 );
not ( n987 , n986 );
and ( n988 , n785 , n945 );
xor ( n989 , n946 , n965 );
and ( n990 , n989 , n784 );
or ( n991 , n988 , n990 );
not ( n992 , n991 );
and ( n993 , n785 , n950 );
xor ( n994 , n951 , n964 );
and ( n995 , n994 , n784 );
or ( n996 , n993 , n995 );
not ( n997 , n996 );
and ( n998 , n785 , n955 );
xor ( n999 , n956 , n963 );
and ( n1000 , n999 , n784 );
or ( n1001 , n998 , n1000 );
not ( n1002 , n1001 );
and ( n1003 , n785 , n960 );
xor ( n1004 , n961 , n962 );
and ( n1005 , n1004 , n784 );
or ( n1006 , n1003 , n1005 );
not ( n1007 , n1006 );
not ( n1008 , n926 );
and ( n1009 , n1007 , n1008 );
and ( n1010 , n1002 , n1009 );
and ( n1011 , n997 , n1010 );
and ( n1012 , n992 , n1011 );
and ( n1013 , n987 , n1012 );
and ( n1014 , n982 , n1013 );
and ( n1015 , n977 , n1014 );
and ( n1016 , n972 , n1015 );
not ( n1017 , n1016 );
and ( n1018 , n1017 , n784 );
and ( n1019 , n926 , n1018 );
not ( n1020 , n1019 );
and ( n1021 , n1020 , n926 );
xor ( n1022 , n926 , n1018 );
xor ( n1023 , n1022 , n1018 );
and ( n1024 , n1023 , n1019 );
or ( n1025 , n1021 , n1024 );
and ( n1026 , n1002 , n1007 );
and ( n1027 , n997 , n1026 );
and ( n1028 , n992 , n1027 );
and ( n1029 , n987 , n1028 );
and ( n1030 , n982 , n1029 );
and ( n1031 , n977 , n1030 );
and ( n1032 , n972 , n1031 );
not ( n1033 , n1032 );
and ( n1034 , n1033 , n784 );
not ( n1035 , n1034 );
and ( n1036 , n785 , n1001 );
xor ( n1037 , n1002 , n1007 );
and ( n1038 , n1037 , n784 );
or ( n1039 , n1036 , n1038 );
and ( n1040 , n1035 , n1039 );
not ( n1041 , n1039 );
xor ( n1042 , n1041 , n1007 );
and ( n1043 , n1042 , n1034 );
or ( n1044 , n1040 , n1043 );
or ( n1045 , n1006 , n1044 );
and ( n1046 , n785 , n996 );
xor ( n1047 , n997 , n1026 );
and ( n1048 , n1047 , n784 );
or ( n1049 , n1046 , n1048 );
and ( n1050 , n1035 , n1049 );
not ( n1051 , n1049 );
and ( n1052 , n1041 , n1007 );
xor ( n1053 , n1051 , n1052 );
and ( n1054 , n1053 , n1034 );
or ( n1055 , n1050 , n1054 );
or ( n1056 , n1045 , n1055 );
and ( n1057 , n1056 , n1034 );
not ( n1058 , n1057 );
and ( n1059 , n1058 , n1006 );
xor ( n1060 , n1006 , n1034 );
xor ( n1061 , n1060 , n1034 );
and ( n1062 , n1061 , n1057 );
or ( n1063 , n1059 , n1062 );
and ( n1064 , n1058 , n1044 );
xor ( n1065 , n1044 , n1034 );
and ( n1066 , n1060 , n1034 );
xor ( n1067 , n1065 , n1066 );
and ( n1068 , n1067 , n1057 );
or ( n1069 , n1064 , n1068 );
and ( n1070 , n1058 , n1055 );
xor ( n1071 , n1055 , n1034 );
and ( n1072 , n1065 , n1066 );
xor ( n1073 , n1071 , n1072 );
and ( n1074 , n1073 , n1057 );
or ( n1075 , n1070 , n1074 );
and ( n1076 , n1063 , n1069 , n1075 );
or ( n1077 , n1025 , n1076 );
not ( n1078 , n1077 );
and ( n1079 , n977 , n982 );
and ( n1080 , n972 , n1079 );
not ( n1081 , n1080 );
and ( n1082 , n1081 , n784 );
not ( n1083 , n1082 );
and ( n1084 , n785 , n976 );
xor ( n1085 , n977 , n982 );
and ( n1086 , n1085 , n784 );
or ( n1087 , n1084 , n1086 );
and ( n1088 , n1083 , n1087 );
not ( n1089 , n1087 );
xor ( n1090 , n1089 , n982 );
and ( n1091 , n1090 , n1082 );
or ( n1092 , n1088 , n1091 );
or ( n1093 , n981 , n1092 );
and ( n1094 , n1093 , n1082 );
not ( n1095 , n1094 );
and ( n1096 , n1095 , n981 );
xor ( n1097 , n981 , n1082 );
xor ( n1098 , n1097 , n1082 );
and ( n1099 , n1098 , n1094 );
or ( n1100 , n1096 , n1099 );
and ( n1101 , n1095 , n1092 );
xor ( n1102 , n1092 , n1082 );
and ( n1103 , n1097 , n1082 );
xor ( n1104 , n1102 , n1103 );
and ( n1105 , n1104 , n1094 );
or ( n1106 , n1101 , n1105 );
and ( n1107 , n1100 , n1106 );
and ( n1108 , n562 , n1107 );
not ( n1109 , n1100 );
and ( n1110 , n1109 , n1106 );
and ( n1111 , n563 , n1110 );
nor ( n1112 , n1109 , n1106 );
and ( n1113 , n564 , n1112 );
nor ( n1114 , n1100 , n1106 );
and ( n1115 , n565 , n1114 );
or ( n1116 , n1108 , n1111 , n1113 , n1115 );
and ( n1117 , n566 , n1110 );
and ( n1118 , n567 , n1112 );
and ( n1119 , n568 , n1114 );
or ( n1120 , 1'b0 , n1117 , n1118 , n1119 );
not ( n1121 , n1120 );
and ( n1122 , n569 , n1107 );
and ( n1123 , n570 , n1110 );
and ( n1124 , n571 , n1112 );
and ( n1125 , n572 , n1114 );
or ( n1126 , n1122 , n1123 , n1124 , n1125 );
and ( n1127 , n1121 , n1126 );
not ( n1128 , n1126 );
not ( n1129 , n1116 );
xor ( n1130 , n1128 , n1129 );
and ( n1131 , n1130 , n1120 );
or ( n1132 , n1127 , n1131 );
or ( n1133 , n1116 , n1132 );
and ( n1134 , n573 , n1107 );
and ( n1135 , n574 , n1110 );
and ( n1136 , n575 , n1112 );
and ( n1137 , n576 , n1114 );
or ( n1138 , n1134 , n1135 , n1136 , n1137 );
and ( n1139 , n1121 , n1138 );
not ( n1140 , n1138 );
and ( n1141 , n1128 , n1129 );
xor ( n1142 , n1140 , n1141 );
and ( n1143 , n1142 , n1120 );
or ( n1144 , n1139 , n1143 );
or ( n1145 , n1133 , n1144 );
not ( n1146 , n577 );
and ( n1147 , n1146 , n1107 );
and ( n1148 , n578 , n1110 );
and ( n1149 , n580 , n1112 );
and ( n1150 , n580 , n1114 );
or ( n1151 , n1147 , n1148 , n1149 , n1150 );
and ( n1152 , n1121 , n1151 );
not ( n1153 , n1151 );
and ( n1154 , n1140 , n1141 );
xor ( n1155 , n1153 , n1154 );
and ( n1156 , n1155 , n1120 );
or ( n1157 , n1152 , n1156 );
or ( n1158 , n1145 , n1157 );
xor ( n1159 , n581 , n577 );
and ( n1160 , n1159 , n1107 );
and ( n1161 , n582 , n1110 );
and ( n1162 , n583 , n1112 );
and ( n1163 , n584 , n1114 );
or ( n1164 , n1160 , n1161 , n1162 , n1163 );
and ( n1165 , n1121 , n1164 );
not ( n1166 , n1164 );
and ( n1167 , n1153 , n1154 );
xor ( n1168 , n1166 , n1167 );
and ( n1169 , n1168 , n1120 );
or ( n1170 , n1165 , n1169 );
or ( n1171 , n1158 , n1170 );
and ( n1172 , n581 , n577 );
xor ( n1173 , n585 , n1172 );
and ( n1174 , n1173 , n1107 );
and ( n1175 , n586 , n1110 );
and ( n1176 , n587 , n1112 );
and ( n1177 , n588 , n1114 );
or ( n1178 , n1174 , n1175 , n1176 , n1177 );
and ( n1179 , n1121 , n1178 );
not ( n1180 , n1178 );
and ( n1181 , n1166 , n1167 );
xor ( n1182 , n1180 , n1181 );
and ( n1183 , n1182 , n1120 );
or ( n1184 , n1179 , n1183 );
or ( n1185 , n1171 , n1184 );
and ( n1186 , n585 , n1172 );
xor ( n1187 , n589 , n1186 );
and ( n1188 , n1187 , n1107 );
and ( n1189 , n590 , n1110 );
and ( n1190 , n591 , n1112 );
and ( n1191 , n592 , n1114 );
or ( n1192 , n1188 , n1189 , n1190 , n1191 );
and ( n1193 , n1121 , n1192 );
not ( n1194 , n1192 );
and ( n1195 , n1180 , n1181 );
xor ( n1196 , n1194 , n1195 );
and ( n1197 , n1196 , n1120 );
or ( n1198 , n1193 , n1197 );
or ( n1199 , n1185 , n1198 );
and ( n1200 , n589 , n1186 );
xor ( n1201 , n593 , n1200 );
and ( n1202 , n1201 , n1107 );
and ( n1203 , n594 , n1110 );
and ( n1204 , n595 , n1112 );
and ( n1205 , n596 , n1114 );
or ( n1206 , n1202 , n1203 , n1204 , n1205 );
and ( n1207 , n1121 , n1206 );
not ( n1208 , n1206 );
and ( n1209 , n1194 , n1195 );
xor ( n1210 , n1208 , n1209 );
and ( n1211 , n1210 , n1120 );
or ( n1212 , n1207 , n1211 );
or ( n1213 , n1199 , n1212 );
and ( n1214 , n593 , n1200 );
xor ( n1215 , n597 , n1214 );
and ( n1216 , n1215 , n1107 );
and ( n1217 , n598 , n1110 );
and ( n1218 , n599 , n1112 );
and ( n1219 , n600 , n1114 );
or ( n1220 , n1216 , n1217 , n1218 , n1219 );
and ( n1221 , n1121 , n1220 );
not ( n1222 , n1220 );
and ( n1223 , n1208 , n1209 );
xor ( n1224 , n1222 , n1223 );
and ( n1225 , n1224 , n1120 );
or ( n1226 , n1221 , n1225 );
or ( n1227 , n1213 , n1226 );
and ( n1228 , n597 , n1214 );
xor ( n1229 , n601 , n1228 );
and ( n1230 , n1229 , n1107 );
and ( n1231 , n602 , n1110 );
and ( n1232 , n603 , n1112 );
and ( n1233 , n604 , n1114 );
or ( n1234 , n1230 , n1231 , n1232 , n1233 );
and ( n1235 , n1121 , n1234 );
not ( n1236 , n1234 );
and ( n1237 , n1222 , n1223 );
xor ( n1238 , n1236 , n1237 );
and ( n1239 , n1238 , n1120 );
or ( n1240 , n1235 , n1239 );
or ( n1241 , n1227 , n1240 );
and ( n1242 , n601 , n1228 );
xor ( n1243 , n605 , n1242 );
and ( n1244 , n1243 , n1107 );
and ( n1245 , n606 , n1110 );
and ( n1246 , n607 , n1112 );
and ( n1247 , n608 , n1114 );
or ( n1248 , n1244 , n1245 , n1246 , n1247 );
and ( n1249 , n1121 , n1248 );
not ( n1250 , n1248 );
and ( n1251 , n1236 , n1237 );
xor ( n1252 , n1250 , n1251 );
and ( n1253 , n1252 , n1120 );
or ( n1254 , n1249 , n1253 );
or ( n1255 , n1241 , n1254 );
and ( n1256 , n605 , n1242 );
xor ( n1257 , n609 , n1256 );
and ( n1258 , n1257 , n1107 );
and ( n1259 , n610 , n1110 );
and ( n1260 , n611 , n1112 );
and ( n1261 , n612 , n1114 );
or ( n1262 , n1258 , n1259 , n1260 , n1261 );
and ( n1263 , n1121 , n1262 );
not ( n1264 , n1262 );
and ( n1265 , n1250 , n1251 );
xor ( n1266 , n1264 , n1265 );
and ( n1267 , n1266 , n1120 );
or ( n1268 , n1263 , n1267 );
or ( n1269 , n1255 , n1268 );
and ( n1270 , n609 , n1256 );
xor ( n1271 , n613 , n1270 );
and ( n1272 , n1271 , n1107 );
and ( n1273 , n614 , n1110 );
and ( n1274 , n615 , n1112 );
and ( n1275 , n616 , n1114 );
or ( n1276 , n1272 , n1273 , n1274 , n1275 );
and ( n1277 , n1121 , n1276 );
not ( n1278 , n1276 );
and ( n1279 , n1264 , n1265 );
xor ( n1280 , n1278 , n1279 );
and ( n1281 , n1280 , n1120 );
or ( n1282 , n1277 , n1281 );
or ( n1283 , n1269 , n1282 );
and ( n1284 , n613 , n1270 );
xor ( n1285 , n617 , n1284 );
and ( n1286 , n1285 , n1107 );
and ( n1287 , n618 , n1110 );
and ( n1288 , n619 , n1112 );
and ( n1289 , n620 , n1114 );
or ( n1290 , n1286 , n1287 , n1288 , n1289 );
and ( n1291 , n1121 , n1290 );
not ( n1292 , n1290 );
and ( n1293 , n1278 , n1279 );
xor ( n1294 , n1292 , n1293 );
and ( n1295 , n1294 , n1120 );
or ( n1296 , n1291 , n1295 );
or ( n1297 , n1283 , n1296 );
and ( n1298 , n617 , n1284 );
xor ( n1299 , n621 , n1298 );
and ( n1300 , n1299 , n1107 );
and ( n1301 , n622 , n1110 );
and ( n1302 , n623 , n1112 );
and ( n1303 , n624 , n1114 );
or ( n1304 , n1300 , n1301 , n1302 , n1303 );
and ( n1305 , n1121 , n1304 );
not ( n1306 , n1304 );
and ( n1307 , n1292 , n1293 );
xor ( n1308 , n1306 , n1307 );
and ( n1309 , n1308 , n1120 );
or ( n1310 , n1305 , n1309 );
or ( n1311 , n1297 , n1310 );
and ( n1312 , n621 , n1298 );
xor ( n1313 , n625 , n1312 );
and ( n1314 , n1313 , n1107 );
and ( n1315 , n626 , n1110 );
and ( n1316 , n627 , n1112 );
and ( n1317 , n628 , n1114 );
or ( n1318 , n1314 , n1315 , n1316 , n1317 );
and ( n1319 , n1121 , n1318 );
not ( n1320 , n1318 );
and ( n1321 , n1306 , n1307 );
xor ( n1322 , n1320 , n1321 );
and ( n1323 , n1322 , n1120 );
or ( n1324 , n1319 , n1323 );
or ( n1325 , n1311 , n1324 );
and ( n1326 , n625 , n1312 );
xor ( n1327 , n629 , n1326 );
and ( n1328 , n1327 , n1107 );
buf ( n1329 , n1110 );
and ( n1330 , n630 , n1112 );
and ( n1331 , n631 , n1114 );
or ( n1332 , n1328 , n1329 , n1330 , n1331 );
and ( n1333 , n1121 , n1332 );
not ( n1334 , n1332 );
and ( n1335 , n1320 , n1321 );
xor ( n1336 , n1334 , n1335 );
and ( n1337 , n1336 , n1120 );
or ( n1338 , n1333 , n1337 );
or ( n1339 , n1325 , n1338 );
and ( n1340 , n629 , n1326 );
xor ( n1341 , n632 , n1340 );
and ( n1342 , n1341 , n1107 );
and ( n1343 , n633 , n1110 );
and ( n1344 , n634 , n1112 );
and ( n1345 , n635 , n1114 );
or ( n1346 , n1342 , n1343 , n1344 , n1345 );
and ( n1347 , n1121 , n1346 );
not ( n1348 , n1346 );
and ( n1349 , n1334 , n1335 );
xor ( n1350 , n1348 , n1349 );
and ( n1351 , n1350 , n1120 );
or ( n1352 , n1347 , n1351 );
or ( n1353 , n1339 , n1352 );
and ( n1354 , n632 , n1340 );
xor ( n1355 , n636 , n1354 );
and ( n1356 , n1355 , n1107 );
and ( n1357 , n637 , n1110 );
and ( n1358 , n638 , n1112 );
and ( n1359 , n639 , n1114 );
or ( n1360 , n1356 , n1357 , n1358 , n1359 );
and ( n1361 , n1121 , n1360 );
not ( n1362 , n1360 );
and ( n1363 , n1348 , n1349 );
xor ( n1364 , n1362 , n1363 );
and ( n1365 , n1364 , n1120 );
or ( n1366 , n1361 , n1365 );
or ( n1367 , n1353 , n1366 );
and ( n1368 , n636 , n1354 );
xor ( n1369 , n640 , n1368 );
and ( n1370 , n1369 , n1107 );
and ( n1371 , n641 , n1110 );
and ( n1372 , n642 , n1112 );
and ( n1373 , n643 , n1114 );
or ( n1374 , n1370 , n1371 , n1372 , n1373 );
and ( n1375 , n1121 , n1374 );
not ( n1376 , n1374 );
and ( n1377 , n1362 , n1363 );
xor ( n1378 , n1376 , n1377 );
and ( n1379 , n1378 , n1120 );
or ( n1380 , n1375 , n1379 );
or ( n1381 , n1367 , n1380 );
and ( n1382 , n640 , n1368 );
xor ( n1383 , n644 , n1382 );
and ( n1384 , n1383 , n1107 );
and ( n1385 , n645 , n1110 );
and ( n1386 , n646 , n1112 );
and ( n1387 , n647 , n1114 );
or ( n1388 , n1384 , n1385 , n1386 , n1387 );
and ( n1389 , n1121 , n1388 );
not ( n1390 , n1388 );
and ( n1391 , n1376 , n1377 );
xor ( n1392 , n1390 , n1391 );
and ( n1393 , n1392 , n1120 );
or ( n1394 , n1389 , n1393 );
or ( n1395 , n1381 , n1394 );
and ( n1396 , n644 , n1382 );
xor ( n1397 , n648 , n1396 );
and ( n1398 , n1397 , n1107 );
and ( n1399 , n649 , n1110 );
and ( n1400 , n650 , n1112 );
and ( n1401 , n651 , n1114 );
or ( n1402 , n1398 , n1399 , n1400 , n1401 );
and ( n1403 , n1121 , n1402 );
not ( n1404 , n1402 );
and ( n1405 , n1390 , n1391 );
xor ( n1406 , n1404 , n1405 );
and ( n1407 , n1406 , n1120 );
or ( n1408 , n1403 , n1407 );
or ( n1409 , n1395 , n1408 );
and ( n1410 , n648 , n1396 );
xor ( n1411 , n652 , n1410 );
and ( n1412 , n1411 , n1107 );
and ( n1413 , n653 , n1110 );
and ( n1414 , n654 , n1112 );
and ( n1415 , n655 , n1114 );
or ( n1416 , n1412 , n1413 , n1414 , n1415 );
and ( n1417 , n1121 , n1416 );
not ( n1418 , n1416 );
and ( n1419 , n1404 , n1405 );
xor ( n1420 , n1418 , n1419 );
and ( n1421 , n1420 , n1120 );
or ( n1422 , n1417 , n1421 );
or ( n1423 , n1409 , n1422 );
and ( n1424 , n652 , n1410 );
xor ( n1425 , n656 , n1424 );
and ( n1426 , n1425 , n1107 );
and ( n1427 , n657 , n1110 );
and ( n1428 , n658 , n1112 );
and ( n1429 , n659 , n1114 );
or ( n1430 , n1426 , n1427 , n1428 , n1429 );
and ( n1431 , n1121 , n1430 );
not ( n1432 , n1430 );
and ( n1433 , n1418 , n1419 );
xor ( n1434 , n1432 , n1433 );
and ( n1435 , n1434 , n1120 );
or ( n1436 , n1431 , n1435 );
or ( n1437 , n1423 , n1436 );
and ( n1438 , n656 , n1424 );
xor ( n1439 , n660 , n1438 );
and ( n1440 , n1439 , n1107 );
and ( n1441 , n661 , n1110 );
and ( n1442 , n662 , n1112 );
and ( n1443 , n663 , n1114 );
or ( n1444 , n1440 , n1441 , n1442 , n1443 );
and ( n1445 , n1121 , n1444 );
not ( n1446 , n1444 );
and ( n1447 , n1432 , n1433 );
xor ( n1448 , n1446 , n1447 );
and ( n1449 , n1448 , n1120 );
or ( n1450 , n1445 , n1449 );
or ( n1451 , n1437 , n1450 );
and ( n1452 , n660 , n1438 );
xor ( n1453 , n664 , n1452 );
and ( n1454 , n1453 , n1107 );
and ( n1455 , n665 , n1110 );
and ( n1456 , n666 , n1112 );
and ( n1457 , n667 , n1114 );
or ( n1458 , n1454 , n1455 , n1456 , n1457 );
and ( n1459 , n1121 , n1458 );
not ( n1460 , n1458 );
and ( n1461 , n1446 , n1447 );
xor ( n1462 , n1460 , n1461 );
and ( n1463 , n1462 , n1120 );
or ( n1464 , n1459 , n1463 );
or ( n1465 , n1451 , n1464 );
and ( n1466 , n664 , n1452 );
xor ( n1467 , n668 , n1466 );
and ( n1468 , n1467 , n1107 );
and ( n1469 , n669 , n1110 );
and ( n1470 , n670 , n1112 );
and ( n1471 , n671 , n1114 );
or ( n1472 , n1468 , n1469 , n1470 , n1471 );
and ( n1473 , n1121 , n1472 );
not ( n1474 , n1472 );
and ( n1475 , n1460 , n1461 );
xor ( n1476 , n1474 , n1475 );
and ( n1477 , n1476 , n1120 );
or ( n1478 , n1473 , n1477 );
or ( n1479 , n1465 , n1478 );
and ( n1480 , n668 , n1466 );
xor ( n1481 , n672 , n1480 );
and ( n1482 , n1481 , n1107 );
and ( n1483 , n673 , n1110 );
and ( n1484 , n674 , n1112 );
and ( n1485 , n675 , n1114 );
or ( n1486 , n1482 , n1483 , n1484 , n1485 );
and ( n1487 , n1121 , n1486 );
not ( n1488 , n1486 );
and ( n1489 , n1474 , n1475 );
xor ( n1490 , n1488 , n1489 );
and ( n1491 , n1490 , n1120 );
or ( n1492 , n1487 , n1491 );
or ( n1493 , n1479 , n1492 );
and ( n1494 , n672 , n1480 );
xor ( n1495 , n676 , n1494 );
and ( n1496 , n1495 , n1107 );
and ( n1497 , n677 , n1110 );
and ( n1498 , n678 , n1112 );
and ( n1499 , n679 , n1114 );
or ( n1500 , n1496 , n1497 , n1498 , n1499 );
and ( n1501 , n1121 , n1500 );
not ( n1502 , n1500 );
and ( n1503 , n1488 , n1489 );
xor ( n1504 , n1502 , n1503 );
and ( n1505 , n1504 , n1120 );
or ( n1506 , n1501 , n1505 );
or ( n1507 , n1493 , n1506 );
and ( n1508 , n1507 , n1120 );
not ( n1509 , n1508 );
and ( n1510 , n1509 , n1310 );
xor ( n1511 , n1310 , n1120 );
xor ( n1512 , n1296 , n1120 );
xor ( n1513 , n1282 , n1120 );
xor ( n1514 , n1268 , n1120 );
xor ( n1515 , n1254 , n1120 );
xor ( n1516 , n1240 , n1120 );
xor ( n1517 , n1226 , n1120 );
xor ( n1518 , n1212 , n1120 );
xor ( n1519 , n1198 , n1120 );
xor ( n1520 , n1184 , n1120 );
xor ( n1521 , n1170 , n1120 );
xor ( n1522 , n1157 , n1120 );
xor ( n1523 , n1144 , n1120 );
xor ( n1524 , n1132 , n1120 );
xor ( n1525 , n1116 , n1120 );
and ( n1526 , n1525 , n1120 );
and ( n1527 , n1524 , n1526 );
and ( n1528 , n1523 , n1527 );
and ( n1529 , n1522 , n1528 );
and ( n1530 , n1521 , n1529 );
and ( n1531 , n1520 , n1530 );
and ( n1532 , n1519 , n1531 );
and ( n1533 , n1518 , n1532 );
and ( n1534 , n1517 , n1533 );
and ( n1535 , n1516 , n1534 );
and ( n1536 , n1515 , n1535 );
and ( n1537 , n1514 , n1536 );
and ( n1538 , n1513 , n1537 );
and ( n1539 , n1512 , n1538 );
xor ( n1540 , n1511 , n1539 );
and ( n1541 , n1540 , n1508 );
or ( n1542 , n1510 , n1541 );
not ( n1543 , n971 );
not ( n1544 , n976 );
not ( n1545 , n981 );
not ( n1546 , n986 );
not ( n1547 , n991 );
and ( n1548 , n1546 , n1547 );
and ( n1549 , n1545 , n1548 );
and ( n1550 , n1544 , n1549 );
and ( n1551 , n1543 , n1550 );
not ( n1552 , n1551 );
and ( n1553 , n1552 , n784 );
not ( n1554 , n1553 );
not ( n1555 , n784 );
and ( n1556 , n1555 , n986 );
xor ( n1557 , n1546 , n1547 );
and ( n1558 , n1557 , n784 );
or ( n1559 , n1556 , n1558 );
and ( n1560 , n1554 , n1559 );
not ( n1561 , n1559 );
xor ( n1562 , n1561 , n1547 );
and ( n1563 , n1562 , n1553 );
or ( n1564 , n1560 , n1563 );
or ( n1565 , n991 , n1564 );
and ( n1566 , n1565 , n1553 );
not ( n1567 , n1566 );
and ( n1568 , n1567 , n991 );
xor ( n1569 , n991 , n1553 );
xor ( n1570 , n1569 , n1553 );
and ( n1571 , n1570 , n1566 );
or ( n1572 , n1568 , n1571 );
and ( n1573 , n1567 , n1564 );
xor ( n1574 , n1564 , n1553 );
and ( n1575 , n1569 , n1553 );
xor ( n1576 , n1574 , n1575 );
and ( n1577 , n1576 , n1566 );
or ( n1578 , n1573 , n1577 );
and ( n1579 , n1572 , n1578 );
and ( n1580 , n1542 , n1579 );
not ( n1581 , n1572 );
and ( n1582 , n1581 , n1578 );
and ( n1583 , n1542 , n1582 );
not ( n1584 , n680 );
not ( n1585 , n1120 );
and ( n1586 , n1585 , n1338 );
not ( n1587 , n1338 );
not ( n1588 , n1324 );
not ( n1589 , n1310 );
not ( n1590 , n1296 );
not ( n1591 , n1282 );
not ( n1592 , n1268 );
not ( n1593 , n1254 );
not ( n1594 , n1240 );
not ( n1595 , n1226 );
not ( n1596 , n1212 );
not ( n1597 , n1198 );
not ( n1598 , n1184 );
not ( n1599 , n1170 );
not ( n1600 , n1157 );
not ( n1601 , n1144 );
not ( n1602 , n1132 );
and ( n1603 , n1601 , n1602 );
and ( n1604 , n1600 , n1603 );
and ( n1605 , n1599 , n1604 );
and ( n1606 , n1598 , n1605 );
and ( n1607 , n1597 , n1606 );
and ( n1608 , n1596 , n1607 );
and ( n1609 , n1595 , n1608 );
and ( n1610 , n1594 , n1609 );
and ( n1611 , n1593 , n1610 );
and ( n1612 , n1592 , n1611 );
and ( n1613 , n1591 , n1612 );
and ( n1614 , n1590 , n1613 );
and ( n1615 , n1589 , n1614 );
and ( n1616 , n1588 , n1615 );
xor ( n1617 , n1587 , n1616 );
and ( n1618 , n1617 , n1120 );
or ( n1619 , n1586 , n1618 );
and ( n1620 , n1584 , n1619 );
not ( n1621 , n1120 );
and ( n1622 , n681 , n1110 );
and ( n1623 , n682 , n1112 );
and ( n1624 , n683 , n1114 );
or ( n1625 , 1'b0 , n1622 , n1623 , n1624 );
not ( n1626 , n1625 );
and ( n1627 , n676 , n1494 );
and ( n1628 , n1627 , n1107 );
and ( n1629 , n684 , n1110 );
and ( n1630 , n685 , n1112 );
and ( n1631 , n686 , n1114 );
or ( n1632 , n1628 , n1629 , n1630 , n1631 );
not ( n1633 , n1632 );
not ( n1634 , n1500 );
and ( n1635 , n1634 , n1503 );
and ( n1636 , n1633 , n1635 );
and ( n1637 , n1626 , n1636 );
xor ( n1638 , n1621 , n1637 );
and ( n1639 , n1638 , n1120 );
not ( n1640 , n1639 );
and ( n1641 , n1121 , n1625 );
xor ( n1642 , n1626 , n1636 );
and ( n1643 , n1642 , n1120 );
or ( n1644 , n1641 , n1643 );
not ( n1645 , n1644 );
and ( n1646 , n1621 , n1632 );
xor ( n1647 , n1633 , n1635 );
and ( n1648 , n1647 , n1120 );
or ( n1649 , n1646 , n1648 );
not ( n1650 , n1649 );
not ( n1651 , n1506 );
not ( n1652 , n1492 );
not ( n1653 , n1478 );
not ( n1654 , n1464 );
not ( n1655 , n1450 );
not ( n1656 , n1436 );
not ( n1657 , n1422 );
not ( n1658 , n1408 );
not ( n1659 , n1394 );
not ( n1660 , n1380 );
not ( n1661 , n1366 );
not ( n1662 , n1352 );
and ( n1663 , n1587 , n1616 );
and ( n1664 , n1662 , n1663 );
and ( n1665 , n1661 , n1664 );
and ( n1666 , n1660 , n1665 );
and ( n1667 , n1659 , n1666 );
and ( n1668 , n1658 , n1667 );
and ( n1669 , n1657 , n1668 );
and ( n1670 , n1656 , n1669 );
and ( n1671 , n1655 , n1670 );
and ( n1672 , n1654 , n1671 );
and ( n1673 , n1653 , n1672 );
and ( n1674 , n1652 , n1673 );
and ( n1675 , n1651 , n1674 );
and ( n1676 , n1650 , n1675 );
and ( n1677 , n1645 , n1676 );
and ( n1678 , n1640 , n1677 );
not ( n1679 , n1678 );
and ( n1680 , n1679 , n1120 );
not ( n1681 , n1680 );
and ( n1682 , n1585 , n1144 );
xor ( n1683 , n1601 , n1602 );
and ( n1684 , n1683 , n1120 );
or ( n1685 , n1682 , n1684 );
and ( n1686 , n1681 , n1685 );
not ( n1687 , n1685 );
xor ( n1688 , n1687 , n1602 );
and ( n1689 , n1688 , n1680 );
or ( n1690 , n1686 , n1689 );
or ( n1691 , n1132 , n1690 );
and ( n1692 , n1585 , n1157 );
xor ( n1693 , n1600 , n1603 );
and ( n1694 , n1693 , n1120 );
or ( n1695 , n1692 , n1694 );
and ( n1696 , n1681 , n1695 );
not ( n1697 , n1695 );
and ( n1698 , n1687 , n1602 );
xor ( n1699 , n1697 , n1698 );
and ( n1700 , n1699 , n1680 );
or ( n1701 , n1696 , n1700 );
or ( n1702 , n1691 , n1701 );
and ( n1703 , n1585 , n1170 );
xor ( n1704 , n1599 , n1604 );
and ( n1705 , n1704 , n1120 );
or ( n1706 , n1703 , n1705 );
and ( n1707 , n1681 , n1706 );
not ( n1708 , n1706 );
and ( n1709 , n1697 , n1698 );
xor ( n1710 , n1708 , n1709 );
and ( n1711 , n1710 , n1680 );
or ( n1712 , n1707 , n1711 );
or ( n1713 , n1702 , n1712 );
and ( n1714 , n1585 , n1184 );
xor ( n1715 , n1598 , n1605 );
and ( n1716 , n1715 , n1120 );
or ( n1717 , n1714 , n1716 );
and ( n1718 , n1681 , n1717 );
not ( n1719 , n1717 );
and ( n1720 , n1708 , n1709 );
xor ( n1721 , n1719 , n1720 );
and ( n1722 , n1721 , n1680 );
or ( n1723 , n1718 , n1722 );
or ( n1724 , n1713 , n1723 );
and ( n1725 , n1585 , n1198 );
xor ( n1726 , n1597 , n1606 );
and ( n1727 , n1726 , n1120 );
or ( n1728 , n1725 , n1727 );
and ( n1729 , n1681 , n1728 );
not ( n1730 , n1728 );
and ( n1731 , n1719 , n1720 );
xor ( n1732 , n1730 , n1731 );
and ( n1733 , n1732 , n1680 );
or ( n1734 , n1729 , n1733 );
or ( n1735 , n1724 , n1734 );
and ( n1736 , n1585 , n1212 );
xor ( n1737 , n1596 , n1607 );
and ( n1738 , n1737 , n1120 );
or ( n1739 , n1736 , n1738 );
and ( n1740 , n1681 , n1739 );
not ( n1741 , n1739 );
and ( n1742 , n1730 , n1731 );
xor ( n1743 , n1741 , n1742 );
and ( n1744 , n1743 , n1680 );
or ( n1745 , n1740 , n1744 );
or ( n1746 , n1735 , n1745 );
and ( n1747 , n1585 , n1226 );
xor ( n1748 , n1595 , n1608 );
and ( n1749 , n1748 , n1120 );
or ( n1750 , n1747 , n1749 );
and ( n1751 , n1681 , n1750 );
not ( n1752 , n1750 );
and ( n1753 , n1741 , n1742 );
xor ( n1754 , n1752 , n1753 );
and ( n1755 , n1754 , n1680 );
or ( n1756 , n1751 , n1755 );
or ( n1757 , n1746 , n1756 );
and ( n1758 , n1585 , n1240 );
xor ( n1759 , n1594 , n1609 );
and ( n1760 , n1759 , n1120 );
or ( n1761 , n1758 , n1760 );
and ( n1762 , n1681 , n1761 );
not ( n1763 , n1761 );
and ( n1764 , n1752 , n1753 );
xor ( n1765 , n1763 , n1764 );
and ( n1766 , n1765 , n1680 );
or ( n1767 , n1762 , n1766 );
or ( n1768 , n1757 , n1767 );
and ( n1769 , n1585 , n1254 );
xor ( n1770 , n1593 , n1610 );
and ( n1771 , n1770 , n1120 );
or ( n1772 , n1769 , n1771 );
and ( n1773 , n1681 , n1772 );
not ( n1774 , n1772 );
and ( n1775 , n1763 , n1764 );
xor ( n1776 , n1774 , n1775 );
and ( n1777 , n1776 , n1680 );
or ( n1778 , n1773 , n1777 );
or ( n1779 , n1768 , n1778 );
and ( n1780 , n1585 , n1268 );
xor ( n1781 , n1592 , n1611 );
and ( n1782 , n1781 , n1120 );
or ( n1783 , n1780 , n1782 );
and ( n1784 , n1681 , n1783 );
not ( n1785 , n1783 );
and ( n1786 , n1774 , n1775 );
xor ( n1787 , n1785 , n1786 );
and ( n1788 , n1787 , n1680 );
or ( n1789 , n1784 , n1788 );
or ( n1790 , n1779 , n1789 );
and ( n1791 , n1585 , n1282 );
xor ( n1792 , n1591 , n1612 );
and ( n1793 , n1792 , n1120 );
or ( n1794 , n1791 , n1793 );
and ( n1795 , n1681 , n1794 );
not ( n1796 , n1794 );
and ( n1797 , n1785 , n1786 );
xor ( n1798 , n1796 , n1797 );
and ( n1799 , n1798 , n1680 );
or ( n1800 , n1795 , n1799 );
or ( n1801 , n1790 , n1800 );
and ( n1802 , n1585 , n1296 );
xor ( n1803 , n1590 , n1613 );
and ( n1804 , n1803 , n1120 );
or ( n1805 , n1802 , n1804 );
and ( n1806 , n1681 , n1805 );
not ( n1807 , n1805 );
and ( n1808 , n1796 , n1797 );
xor ( n1809 , n1807 , n1808 );
and ( n1810 , n1809 , n1680 );
or ( n1811 , n1806 , n1810 );
or ( n1812 , n1801 , n1811 );
and ( n1813 , n1585 , n1310 );
xor ( n1814 , n1589 , n1614 );
and ( n1815 , n1814 , n1120 );
or ( n1816 , n1813 , n1815 );
and ( n1817 , n1681 , n1816 );
not ( n1818 , n1816 );
and ( n1819 , n1807 , n1808 );
xor ( n1820 , n1818 , n1819 );
and ( n1821 , n1820 , n1680 );
or ( n1822 , n1817 , n1821 );
or ( n1823 , n1812 , n1822 );
and ( n1824 , n1585 , n1324 );
xor ( n1825 , n1588 , n1615 );
and ( n1826 , n1825 , n1120 );
or ( n1827 , n1824 , n1826 );
and ( n1828 , n1681 , n1827 );
not ( n1829 , n1827 );
and ( n1830 , n1818 , n1819 );
xor ( n1831 , n1829 , n1830 );
and ( n1832 , n1831 , n1680 );
or ( n1833 , n1828 , n1832 );
or ( n1834 , n1823 , n1833 );
and ( n1835 , n1681 , n1619 );
not ( n1836 , n1619 );
and ( n1837 , n1829 , n1830 );
xor ( n1838 , n1836 , n1837 );
and ( n1839 , n1838 , n1680 );
or ( n1840 , n1835 , n1839 );
or ( n1841 , n1834 , n1840 );
and ( n1842 , n1585 , n1352 );
xor ( n1843 , n1662 , n1663 );
and ( n1844 , n1843 , n1120 );
or ( n1845 , n1842 , n1844 );
and ( n1846 , n1681 , n1845 );
not ( n1847 , n1845 );
and ( n1848 , n1836 , n1837 );
xor ( n1849 , n1847 , n1848 );
and ( n1850 , n1849 , n1680 );
or ( n1851 , n1846 , n1850 );
or ( n1852 , n1841 , n1851 );
and ( n1853 , n1585 , n1366 );
xor ( n1854 , n1661 , n1664 );
and ( n1855 , n1854 , n1120 );
or ( n1856 , n1853 , n1855 );
and ( n1857 , n1681 , n1856 );
not ( n1858 , n1856 );
and ( n1859 , n1847 , n1848 );
xor ( n1860 , n1858 , n1859 );
and ( n1861 , n1860 , n1680 );
or ( n1862 , n1857 , n1861 );
or ( n1863 , n1852 , n1862 );
and ( n1864 , n1585 , n1380 );
xor ( n1865 , n1660 , n1665 );
and ( n1866 , n1865 , n1120 );
or ( n1867 , n1864 , n1866 );
and ( n1868 , n1681 , n1867 );
not ( n1869 , n1867 );
and ( n1870 , n1858 , n1859 );
xor ( n1871 , n1869 , n1870 );
and ( n1872 , n1871 , n1680 );
or ( n1873 , n1868 , n1872 );
or ( n1874 , n1863 , n1873 );
and ( n1875 , n1585 , n1394 );
xor ( n1876 , n1659 , n1666 );
and ( n1877 , n1876 , n1120 );
or ( n1878 , n1875 , n1877 );
and ( n1879 , n1681 , n1878 );
not ( n1880 , n1878 );
and ( n1881 , n1869 , n1870 );
xor ( n1882 , n1880 , n1881 );
and ( n1883 , n1882 , n1680 );
or ( n1884 , n1879 , n1883 );
or ( n1885 , n1874 , n1884 );
and ( n1886 , n1585 , n1408 );
xor ( n1887 , n1658 , n1667 );
and ( n1888 , n1887 , n1120 );
or ( n1889 , n1886 , n1888 );
and ( n1890 , n1681 , n1889 );
not ( n1891 , n1889 );
and ( n1892 , n1880 , n1881 );
xor ( n1893 , n1891 , n1892 );
and ( n1894 , n1893 , n1680 );
or ( n1895 , n1890 , n1894 );
or ( n1896 , n1885 , n1895 );
and ( n1897 , n1585 , n1422 );
xor ( n1898 , n1657 , n1668 );
and ( n1899 , n1898 , n1120 );
or ( n1900 , n1897 , n1899 );
and ( n1901 , n1681 , n1900 );
not ( n1902 , n1900 );
and ( n1903 , n1891 , n1892 );
xor ( n1904 , n1902 , n1903 );
and ( n1905 , n1904 , n1680 );
or ( n1906 , n1901 , n1905 );
or ( n1907 , n1896 , n1906 );
and ( n1908 , n1585 , n1436 );
xor ( n1909 , n1656 , n1669 );
and ( n1910 , n1909 , n1120 );
or ( n1911 , n1908 , n1910 );
and ( n1912 , n1681 , n1911 );
not ( n1913 , n1911 );
and ( n1914 , n1902 , n1903 );
xor ( n1915 , n1913 , n1914 );
and ( n1916 , n1915 , n1680 );
or ( n1917 , n1912 , n1916 );
or ( n1918 , n1907 , n1917 );
and ( n1919 , n1585 , n1450 );
xor ( n1920 , n1655 , n1670 );
and ( n1921 , n1920 , n1120 );
or ( n1922 , n1919 , n1921 );
and ( n1923 , n1681 , n1922 );
not ( n1924 , n1922 );
and ( n1925 , n1913 , n1914 );
xor ( n1926 , n1924 , n1925 );
and ( n1927 , n1926 , n1680 );
or ( n1928 , n1923 , n1927 );
or ( n1929 , n1918 , n1928 );
and ( n1930 , n1585 , n1464 );
xor ( n1931 , n1654 , n1671 );
and ( n1932 , n1931 , n1120 );
or ( n1933 , n1930 , n1932 );
and ( n1934 , n1681 , n1933 );
not ( n1935 , n1933 );
and ( n1936 , n1924 , n1925 );
xor ( n1937 , n1935 , n1936 );
and ( n1938 , n1937 , n1680 );
or ( n1939 , n1934 , n1938 );
or ( n1940 , n1929 , n1939 );
and ( n1941 , n1585 , n1478 );
xor ( n1942 , n1653 , n1672 );
and ( n1943 , n1942 , n1120 );
or ( n1944 , n1941 , n1943 );
and ( n1945 , n1681 , n1944 );
not ( n1946 , n1944 );
and ( n1947 , n1935 , n1936 );
xor ( n1948 , n1946 , n1947 );
and ( n1949 , n1948 , n1680 );
or ( n1950 , n1945 , n1949 );
or ( n1951 , n1940 , n1950 );
and ( n1952 , n1585 , n1492 );
xor ( n1953 , n1652 , n1673 );
and ( n1954 , n1953 , n1120 );
or ( n1955 , n1952 , n1954 );
and ( n1956 , n1681 , n1955 );
not ( n1957 , n1955 );
and ( n1958 , n1946 , n1947 );
xor ( n1959 , n1957 , n1958 );
and ( n1960 , n1959 , n1680 );
or ( n1961 , n1956 , n1960 );
or ( n1962 , n1951 , n1961 );
and ( n1963 , n1585 , n1506 );
xor ( n1964 , n1651 , n1674 );
and ( n1965 , n1964 , n1120 );
or ( n1966 , n1963 , n1965 );
and ( n1967 , n1681 , n1966 );
not ( n1968 , n1966 );
and ( n1969 , n1957 , n1958 );
xor ( n1970 , n1968 , n1969 );
and ( n1971 , n1970 , n1680 );
or ( n1972 , n1967 , n1971 );
or ( n1973 , n1962 , n1972 );
and ( n1974 , n1585 , n1649 );
xor ( n1975 , n1650 , n1675 );
and ( n1976 , n1975 , n1120 );
or ( n1977 , n1974 , n1976 );
and ( n1978 , n1681 , n1977 );
not ( n1979 , n1977 );
and ( n1980 , n1968 , n1969 );
xor ( n1981 , n1979 , n1980 );
and ( n1982 , n1981 , n1680 );
or ( n1983 , n1978 , n1982 );
or ( n1984 , n1973 , n1983 );
and ( n1985 , n1984 , n1680 );
not ( n1986 , n1985 );
and ( n1987 , n1986 , n1840 );
xor ( n1988 , n1840 , n1680 );
xor ( n1989 , n1833 , n1680 );
xor ( n1990 , n1822 , n1680 );
xor ( n1991 , n1811 , n1680 );
xor ( n1992 , n1800 , n1680 );
xor ( n1993 , n1789 , n1680 );
xor ( n1994 , n1778 , n1680 );
xor ( n1995 , n1767 , n1680 );
xor ( n1996 , n1756 , n1680 );
xor ( n1997 , n1745 , n1680 );
xor ( n1998 , n1734 , n1680 );
xor ( n1999 , n1723 , n1680 );
xor ( n2000 , n1712 , n1680 );
xor ( n2001 , n1701 , n1680 );
xor ( n2002 , n1690 , n1680 );
xor ( n2003 , n1132 , n1680 );
and ( n2004 , n2003 , n1680 );
and ( n2005 , n2002 , n2004 );
and ( n2006 , n2001 , n2005 );
and ( n2007 , n2000 , n2006 );
and ( n2008 , n1999 , n2007 );
and ( n2009 , n1998 , n2008 );
and ( n2010 , n1997 , n2009 );
and ( n2011 , n1996 , n2010 );
and ( n2012 , n1995 , n2011 );
and ( n2013 , n1994 , n2012 );
and ( n2014 , n1993 , n2013 );
and ( n2015 , n1992 , n2014 );
and ( n2016 , n1991 , n2015 );
and ( n2017 , n1990 , n2016 );
and ( n2018 , n1989 , n2017 );
xor ( n2019 , n1988 , n2018 );
and ( n2020 , n2019 , n1985 );
or ( n2021 , n1987 , n2020 );
and ( n2022 , n2021 , n680 );
or ( n2023 , n1620 , n2022 );
nor ( n2024 , n1581 , n1578 );
and ( n2025 , n2023 , n2024 );
nor ( n2026 , n1572 , n1578 );
and ( n2027 , n1619 , n2026 );
or ( n2028 , n1580 , n1583 , n2025 , n2027 );
not ( n2029 , n1063 );
not ( n2030 , n1075 );
nor ( n2031 , n2029 , n1069 , n2030 );
not ( n2032 , n2031 );
nor ( n2033 , n1063 , n1069 , n2030 );
not ( n2034 , n2033 );
and ( n2035 , n1063 , n1069 , n2030 );
not ( n2036 , n2035 );
and ( n2037 , n2029 , n1069 , n2030 );
not ( n2038 , n2037 );
nor ( n2039 , n2029 , n1069 , n1075 );
not ( n2040 , n2039 );
nor ( n2041 , n1063 , n1069 , n1075 );
not ( n2042 , n2041 );
and ( n2043 , n2042 , n687 );
and ( n2044 , n2040 , n2043 );
or ( n2045 , n2044 , n2039 );
and ( n2046 , n2038 , n2045 );
and ( n2047 , n2036 , n2046 );
or ( n2048 , n2047 , n2035 );
and ( n2049 , n2034 , n2048 );
not ( n2050 , n680 );
and ( n2051 , n2050 , n687 );
or ( n2052 , n2051 , n680 );
and ( n2053 , n2052 , n2033 );
or ( n2054 , n2049 , n2053 );
and ( n2055 , n2032 , n2054 );
and ( n2056 , n680 , n687 );
or ( n2057 , n2056 , n2050 );
and ( n2058 , n2057 , n2031 );
or ( n2059 , n2055 , n2058 );
not ( n2060 , n2059 );
not ( n2061 , n2031 );
not ( n2062 , n2033 );
not ( n2063 , n2035 );
not ( n2064 , n2037 );
not ( n2065 , n2039 );
not ( n2066 , n2041 );
and ( n2067 , n2066 , n688 );
and ( n2068 , n2065 , n2067 );
and ( n2069 , n2064 , n2068 );
or ( n2070 , n2069 , n2037 );
and ( n2071 , n2063 , n2070 );
or ( n2072 , n2071 , n2035 );
and ( n2073 , n2062 , n2072 );
not ( n2074 , n680 );
and ( n2075 , n2074 , n688 );
or ( n2076 , n2075 , n680 );
and ( n2077 , n2076 , n2033 );
or ( n2078 , n2073 , n2077 );
and ( n2079 , n2061 , n2078 );
and ( n2080 , n680 , n688 );
or ( n2081 , n2080 , n2050 );
and ( n2082 , n2081 , n2031 );
or ( n2083 , n2079 , n2082 );
nor ( n2084 , n2060 , n2083 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
and ( n2085 , n2028 , n2084 );
nor ( n2086 , n2059 , n2083 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
not ( n2087 , n2083 );
nor ( n2088 , n2059 , n2087 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
or ( n2089 , n2086 , n2088 );
nor ( n2090 , n2060 , n2087 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 );
or ( n2091 , n2089 , n2090 );
and ( n2092 , n627 , n2091 );
or ( n2093 , n2085 , n2092 );
and ( n2094 , n1555 , n810 );
not ( n2095 , n810 );
xor ( n2096 , n2095 , n919 );
and ( n2097 , n2096 , n784 );
or ( n2098 , n2094 , n2097 );
not ( n2099 , n996 );
not ( n2100 , n1001 );
not ( n2101 , n1006 );
not ( n2102 , n926 );
and ( n2103 , n1555 , n795 );
not ( n2104 , n795 );
xor ( n2105 , n2104 , n922 );
and ( n2106 , n2105 , n784 );
or ( n2107 , n2103 , n2106 );
not ( n2108 , n2107 );
and ( n2109 , n1555 , n800 );
not ( n2110 , n800 );
xor ( n2111 , n2110 , n921 );
and ( n2112 , n2111 , n784 );
or ( n2113 , n2109 , n2112 );
not ( n2114 , n2113 );
and ( n2115 , n1555 , n805 );
not ( n2116 , n805 );
xor ( n2117 , n2116 , n920 );
and ( n2118 , n2117 , n784 );
or ( n2119 , n2115 , n2118 );
not ( n2120 , n2119 );
not ( n2121 , n2098 );
and ( n2122 , n2120 , n2121 );
and ( n2123 , n2114 , n2122 );
and ( n2124 , n2108 , n2123 );
and ( n2125 , n2102 , n2124 );
and ( n2126 , n2101 , n2125 );
and ( n2127 , n2100 , n2126 );
and ( n2128 , n2099 , n2127 );
and ( n2129 , n1547 , n2128 );
and ( n2130 , n1546 , n2129 );
and ( n2131 , n1545 , n2130 );
and ( n2132 , n1544 , n2131 );
and ( n2133 , n1543 , n2132 );
not ( n2134 , n2133 );
and ( n2135 , n2134 , n784 );
not ( n2136 , n2135 );
and ( n2137 , n1555 , n2119 );
xor ( n2138 , n2120 , n2121 );
and ( n2139 , n2138 , n784 );
or ( n2140 , n2137 , n2139 );
and ( n2141 , n2136 , n2140 );
not ( n2142 , n2140 );
xor ( n2143 , n2142 , n2121 );
and ( n2144 , n2143 , n2135 );
or ( n2145 , n2141 , n2144 );
or ( n2146 , n2098 , n2145 );
and ( n2147 , n1555 , n2113 );
xor ( n2148 , n2114 , n2122 );
and ( n2149 , n2148 , n784 );
or ( n2150 , n2147 , n2149 );
and ( n2151 , n2136 , n2150 );
not ( n2152 , n2150 );
and ( n2153 , n2142 , n2121 );
xor ( n2154 , n2152 , n2153 );
and ( n2155 , n2154 , n2135 );
or ( n2156 , n2151 , n2155 );
or ( n2157 , n2146 , n2156 );
and ( n2158 , n1555 , n2107 );
xor ( n2159 , n2108 , n2123 );
and ( n2160 , n2159 , n784 );
or ( n2161 , n2158 , n2160 );
and ( n2162 , n2136 , n2161 );
not ( n2163 , n2161 );
and ( n2164 , n2152 , n2153 );
xor ( n2165 , n2163 , n2164 );
and ( n2166 , n2165 , n2135 );
or ( n2167 , n2162 , n2166 );
or ( n2168 , n2157 , n2167 );
and ( n2169 , n2168 , n2135 );
not ( n2170 , n2169 );
and ( n2171 , n2170 , n2098 );
xor ( n2172 , n2098 , n2135 );
xor ( n2173 , n2172 , n2135 );
and ( n2174 , n2173 , n2169 );
or ( n2175 , n2171 , n2174 );
not ( n2176 , n2175 );
and ( n2177 , n2170 , n2145 );
xor ( n2178 , n2145 , n2135 );
and ( n2179 , n2172 , n2135 );
xor ( n2180 , n2178 , n2179 );
and ( n2181 , n2180 , n2169 );
or ( n2182 , n2177 , n2181 );
not ( n2183 , n2182 );
and ( n2184 , n2170 , n2156 );
xor ( n2185 , n2156 , n2135 );
and ( n2186 , n2178 , n2179 );
xor ( n2187 , n2185 , n2186 );
and ( n2188 , n2187 , n2169 );
or ( n2189 , n2184 , n2188 );
and ( n2190 , n2170 , n2167 );
xor ( n2191 , n2167 , n2135 );
and ( n2192 , n2185 , n2186 );
xor ( n2193 , n2191 , n2192 );
and ( n2194 , n2193 , n2169 );
or ( n2195 , n2190 , n2194 );
and ( n2196 , n2176 , n2183 , n2189 , n2195 );
and ( n2197 , n2093 , n2196 );
or ( n2198 , n2024 , n1582 );
or ( n2199 , n2198 , n1579 );
and ( n2200 , n689 , n2199 );
not ( n2201 , n784 );
and ( n2202 , n2201 , n900 );
not ( n2203 , n900 );
not ( n2204 , n561 );
xor ( n2205 , n2203 , n2204 );
and ( n2206 , n2205 , n784 );
or ( n2207 , n2202 , n2206 );
or ( n2208 , n561 , n2207 );
and ( n2209 , n2201 , n895 );
not ( n2210 , n895 );
xor ( n2211 , n2210 , n902 );
and ( n2212 , n2211 , n784 );
or ( n2213 , n2209 , n2212 );
or ( n2214 , n2208 , n2213 );
and ( n2215 , n2201 , n890 );
not ( n2216 , n890 );
xor ( n2217 , n2216 , n903 );
and ( n2218 , n2217 , n784 );
or ( n2219 , n2215 , n2218 );
or ( n2220 , n2214 , n2219 );
and ( n2221 , n2201 , n885 );
not ( n2222 , n885 );
xor ( n2223 , n2222 , n904 );
and ( n2224 , n2223 , n784 );
or ( n2225 , n2221 , n2224 );
or ( n2226 , n2220 , n2225 );
and ( n2227 , n2201 , n880 );
not ( n2228 , n880 );
xor ( n2229 , n2228 , n905 );
and ( n2230 , n2229 , n784 );
or ( n2231 , n2227 , n2230 );
or ( n2232 , n2226 , n2231 );
and ( n2233 , n2201 , n875 );
not ( n2234 , n875 );
xor ( n2235 , n2234 , n906 );
and ( n2236 , n2235 , n784 );
or ( n2237 , n2233 , n2236 );
or ( n2238 , n2232 , n2237 );
and ( n2239 , n2201 , n870 );
not ( n2240 , n870 );
xor ( n2241 , n2240 , n907 );
and ( n2242 , n2241 , n784 );
or ( n2243 , n2239 , n2242 );
or ( n2244 , n2238 , n2243 );
and ( n2245 , n2201 , n865 );
not ( n2246 , n865 );
xor ( n2247 , n2246 , n908 );
and ( n2248 , n2247 , n784 );
or ( n2249 , n2245 , n2248 );
or ( n2250 , n2244 , n2249 );
and ( n2251 , n2201 , n860 );
not ( n2252 , n860 );
xor ( n2253 , n2252 , n909 );
and ( n2254 , n2253 , n784 );
or ( n2255 , n2251 , n2254 );
or ( n2256 , n2250 , n2255 );
and ( n2257 , n2201 , n855 );
not ( n2258 , n855 );
xor ( n2259 , n2258 , n910 );
and ( n2260 , n2259 , n784 );
or ( n2261 , n2257 , n2260 );
or ( n2262 , n2256 , n2261 );
and ( n2263 , n2201 , n850 );
not ( n2264 , n850 );
xor ( n2265 , n2264 , n911 );
and ( n2266 , n2265 , n784 );
or ( n2267 , n2263 , n2266 );
or ( n2268 , n2262 , n2267 );
and ( n2269 , n2201 , n845 );
not ( n2270 , n845 );
xor ( n2271 , n2270 , n912 );
and ( n2272 , n2271 , n784 );
or ( n2273 , n2269 , n2272 );
or ( n2274 , n2268 , n2273 );
and ( n2275 , n2201 , n840 );
not ( n2276 , n840 );
xor ( n2277 , n2276 , n913 );
and ( n2278 , n2277 , n784 );
or ( n2279 , n2275 , n2278 );
or ( n2280 , n2274 , n2279 );
and ( n2281 , n2201 , n835 );
not ( n2282 , n835 );
xor ( n2283 , n2282 , n914 );
and ( n2284 , n2283 , n784 );
or ( n2285 , n2281 , n2284 );
or ( n2286 , n2280 , n2285 );
and ( n2287 , n2201 , n830 );
not ( n2288 , n830 );
xor ( n2289 , n2288 , n915 );
and ( n2290 , n2289 , n784 );
or ( n2291 , n2287 , n2290 );
or ( n2292 , n2286 , n2291 );
and ( n2293 , n2201 , n825 );
not ( n2294 , n825 );
xor ( n2295 , n2294 , n916 );
and ( n2296 , n2295 , n784 );
or ( n2297 , n2293 , n2296 );
or ( n2298 , n2292 , n2297 );
and ( n2299 , n2201 , n820 );
not ( n2300 , n820 );
xor ( n2301 , n2300 , n917 );
and ( n2302 , n2301 , n784 );
or ( n2303 , n2299 , n2302 );
or ( n2304 , n2298 , n2303 );
and ( n2305 , n2201 , n815 );
not ( n2306 , n815 );
xor ( n2307 , n2306 , n918 );
and ( n2308 , n2307 , n784 );
or ( n2309 , n2305 , n2308 );
or ( n2310 , n2304 , n2309 );
or ( n2311 , n2310 , n2098 );
and ( n2312 , n2311 , n784 );
not ( n2313 , n2312 );
and ( n2314 , n2313 , n561 );
xor ( n2315 , n561 , n784 );
xor ( n2316 , n2315 , n784 );
and ( n2317 , n2316 , n2312 );
or ( n2318 , n2314 , n2317 );
and ( n2319 , n2318 , n2026 );
or ( n2320 , n2200 , n2319 );
xor ( n2321 , n1116 , n2320 );
and ( n2322 , n690 , n2199 );
not ( n2323 , n2322 );
xor ( n2324 , n1120 , n2323 );
and ( n2325 , n691 , n2199 );
not ( n2326 , n2325 );
and ( n2327 , n2326 , n1625 );
not ( n2328 , n2325 );
and ( n2329 , n692 , n2199 );
not ( n2330 , n2329 );
and ( n2331 , n2330 , n1632 );
not ( n2332 , n2329 );
and ( n2333 , n693 , n2199 );
not ( n2334 , n2333 );
and ( n2335 , n2334 , n1500 );
not ( n2336 , n2333 );
and ( n2337 , n694 , n2199 );
not ( n2338 , n2337 );
and ( n2339 , n2338 , n1486 );
not ( n2340 , n2337 );
and ( n2341 , n695 , n2199 );
not ( n2342 , n2341 );
and ( n2343 , n2342 , n1472 );
not ( n2344 , n2341 );
and ( n2345 , n696 , n2199 );
not ( n2346 , n2345 );
and ( n2347 , n2346 , n1458 );
not ( n2348 , n2345 );
and ( n2349 , n697 , n2199 );
not ( n2350 , n2349 );
and ( n2351 , n2350 , n1444 );
not ( n2352 , n2349 );
and ( n2353 , n698 , n2199 );
not ( n2354 , n2353 );
and ( n2355 , n2354 , n1430 );
not ( n2356 , n2353 );
and ( n2357 , n699 , n2199 );
not ( n2358 , n2357 );
and ( n2359 , n2358 , n1416 );
not ( n2360 , n2357 );
and ( n2361 , n700 , n2199 );
not ( n2362 , n2361 );
and ( n2363 , n2362 , n1402 );
not ( n2364 , n2361 );
and ( n2365 , n701 , n2199 );
not ( n2366 , n2365 );
and ( n2367 , n2366 , n1388 );
not ( n2368 , n2365 );
and ( n2369 , n702 , n2199 );
and ( n2370 , n2313 , n2098 );
xor ( n2371 , n2098 , n784 );
xor ( n2372 , n2309 , n784 );
xor ( n2373 , n2303 , n784 );
xor ( n2374 , n2297 , n784 );
xor ( n2375 , n2291 , n784 );
xor ( n2376 , n2285 , n784 );
xor ( n2377 , n2279 , n784 );
xor ( n2378 , n2273 , n784 );
xor ( n2379 , n2267 , n784 );
xor ( n2380 , n2261 , n784 );
xor ( n2381 , n2255 , n784 );
xor ( n2382 , n2249 , n784 );
xor ( n2383 , n2243 , n784 );
xor ( n2384 , n2237 , n784 );
xor ( n2385 , n2231 , n784 );
xor ( n2386 , n2225 , n784 );
xor ( n2387 , n2219 , n784 );
xor ( n2388 , n2213 , n784 );
xor ( n2389 , n2207 , n784 );
and ( n2390 , n2315 , n784 );
and ( n2391 , n2389 , n2390 );
and ( n2392 , n2388 , n2391 );
and ( n2393 , n2387 , n2392 );
and ( n2394 , n2386 , n2393 );
and ( n2395 , n2385 , n2394 );
and ( n2396 , n2384 , n2395 );
and ( n2397 , n2383 , n2396 );
and ( n2398 , n2382 , n2397 );
and ( n2399 , n2381 , n2398 );
and ( n2400 , n2380 , n2399 );
and ( n2401 , n2379 , n2400 );
and ( n2402 , n2378 , n2401 );
and ( n2403 , n2377 , n2402 );
and ( n2404 , n2376 , n2403 );
and ( n2405 , n2375 , n2404 );
and ( n2406 , n2374 , n2405 );
and ( n2407 , n2373 , n2406 );
and ( n2408 , n2372 , n2407 );
xor ( n2409 , n2371 , n2408 );
and ( n2410 , n2409 , n2312 );
or ( n2411 , n2370 , n2410 );
and ( n2412 , n2411 , n2026 );
or ( n2413 , n2369 , n2412 );
not ( n2414 , n2413 );
and ( n2415 , n2414 , n1374 );
not ( n2416 , n2413 );
and ( n2417 , n703 , n2199 );
and ( n2418 , n2313 , n2309 );
xor ( n2419 , n2372 , n2407 );
and ( n2420 , n2419 , n2312 );
or ( n2421 , n2418 , n2420 );
and ( n2422 , n2421 , n2026 );
or ( n2423 , n2417 , n2422 );
not ( n2424 , n2423 );
and ( n2425 , n2424 , n1360 );
not ( n2426 , n2423 );
and ( n2427 , n704 , n2199 );
and ( n2428 , n2313 , n2303 );
xor ( n2429 , n2373 , n2406 );
and ( n2430 , n2429 , n2312 );
or ( n2431 , n2428 , n2430 );
and ( n2432 , n2431 , n2026 );
or ( n2433 , n2427 , n2432 );
not ( n2434 , n2433 );
and ( n2435 , n2434 , n1346 );
not ( n2436 , n2433 );
and ( n2437 , n705 , n2199 );
and ( n2438 , n2313 , n2297 );
xor ( n2439 , n2374 , n2405 );
and ( n2440 , n2439 , n2312 );
or ( n2441 , n2438 , n2440 );
and ( n2442 , n2441 , n2026 );
or ( n2443 , n2437 , n2442 );
not ( n2444 , n2443 );
and ( n2445 , n2444 , n1332 );
not ( n2446 , n2443 );
and ( n2447 , n706 , n2199 );
and ( n2448 , n2313 , n2291 );
xor ( n2449 , n2375 , n2404 );
and ( n2450 , n2449 , n2312 );
or ( n2451 , n2448 , n2450 );
and ( n2452 , n2451 , n2026 );
or ( n2453 , n2447 , n2452 );
not ( n2454 , n2453 );
and ( n2455 , n2454 , n1318 );
not ( n2456 , n2453 );
and ( n2457 , n707 , n2199 );
and ( n2458 , n2313 , n2285 );
xor ( n2459 , n2376 , n2403 );
and ( n2460 , n2459 , n2312 );
or ( n2461 , n2458 , n2460 );
and ( n2462 , n2461 , n2026 );
or ( n2463 , n2457 , n2462 );
not ( n2464 , n2463 );
and ( n2465 , n2464 , n1304 );
not ( n2466 , n2463 );
and ( n2467 , n708 , n2199 );
and ( n2468 , n2313 , n2279 );
xor ( n2469 , n2377 , n2402 );
and ( n2470 , n2469 , n2312 );
or ( n2471 , n2468 , n2470 );
and ( n2472 , n2471 , n2026 );
or ( n2473 , n2467 , n2472 );
not ( n2474 , n2473 );
and ( n2475 , n2474 , n1290 );
not ( n2476 , n2473 );
and ( n2477 , n709 , n2199 );
and ( n2478 , n2313 , n2273 );
xor ( n2479 , n2378 , n2401 );
and ( n2480 , n2479 , n2312 );
or ( n2481 , n2478 , n2480 );
and ( n2482 , n2481 , n2026 );
or ( n2483 , n2477 , n2482 );
not ( n2484 , n2483 );
and ( n2485 , n2484 , n1276 );
not ( n2486 , n2483 );
and ( n2487 , n710 , n2199 );
and ( n2488 , n2313 , n2267 );
xor ( n2489 , n2379 , n2400 );
and ( n2490 , n2489 , n2312 );
or ( n2491 , n2488 , n2490 );
and ( n2492 , n2491 , n2026 );
or ( n2493 , n2487 , n2492 );
not ( n2494 , n2493 );
and ( n2495 , n2494 , n1262 );
not ( n2496 , n2493 );
and ( n2497 , n711 , n2199 );
and ( n2498 , n2313 , n2261 );
xor ( n2499 , n2380 , n2399 );
and ( n2500 , n2499 , n2312 );
or ( n2501 , n2498 , n2500 );
and ( n2502 , n2501 , n2026 );
or ( n2503 , n2497 , n2502 );
not ( n2504 , n2503 );
and ( n2505 , n2504 , n1248 );
not ( n2506 , n2503 );
and ( n2507 , n712 , n2199 );
and ( n2508 , n2313 , n2255 );
xor ( n2509 , n2381 , n2398 );
and ( n2510 , n2509 , n2312 );
or ( n2511 , n2508 , n2510 );
and ( n2512 , n2511 , n2026 );
or ( n2513 , n2507 , n2512 );
not ( n2514 , n2513 );
and ( n2515 , n2514 , n1234 );
not ( n2516 , n2513 );
and ( n2517 , n713 , n2199 );
and ( n2518 , n2313 , n2249 );
xor ( n2519 , n2382 , n2397 );
and ( n2520 , n2519 , n2312 );
or ( n2521 , n2518 , n2520 );
and ( n2522 , n2521 , n2026 );
or ( n2523 , n2517 , n2522 );
not ( n2524 , n2523 );
and ( n2525 , n2524 , n1220 );
not ( n2526 , n2523 );
and ( n2527 , n714 , n2199 );
and ( n2528 , n2313 , n2243 );
xor ( n2529 , n2383 , n2396 );
and ( n2530 , n2529 , n2312 );
or ( n2531 , n2528 , n2530 );
and ( n2532 , n2531 , n2026 );
or ( n2533 , n2527 , n2532 );
not ( n2534 , n2533 );
and ( n2535 , n2534 , n1206 );
not ( n2536 , n2533 );
and ( n2537 , n715 , n2199 );
and ( n2538 , n2313 , n2237 );
xor ( n2539 , n2384 , n2395 );
and ( n2540 , n2539 , n2312 );
or ( n2541 , n2538 , n2540 );
and ( n2542 , n2541 , n2026 );
or ( n2543 , n2537 , n2542 );
not ( n2544 , n2543 );
and ( n2545 , n2544 , n1192 );
not ( n2546 , n2543 );
and ( n2547 , n716 , n2199 );
and ( n2548 , n2313 , n2231 );
xor ( n2549 , n2385 , n2394 );
and ( n2550 , n2549 , n2312 );
or ( n2551 , n2548 , n2550 );
and ( n2552 , n2551 , n2026 );
or ( n2553 , n2547 , n2552 );
not ( n2554 , n2553 );
and ( n2555 , n2554 , n1178 );
not ( n2556 , n2553 );
and ( n2557 , n717 , n2199 );
and ( n2558 , n2313 , n2225 );
xor ( n2559 , n2386 , n2393 );
and ( n2560 , n2559 , n2312 );
or ( n2561 , n2558 , n2560 );
and ( n2562 , n2561 , n2026 );
or ( n2563 , n2557 , n2562 );
not ( n2564 , n2563 );
and ( n2565 , n2564 , n1164 );
not ( n2566 , n2563 );
and ( n2567 , n718 , n2199 );
and ( n2568 , n2313 , n2219 );
xor ( n2569 , n2387 , n2392 );
and ( n2570 , n2569 , n2312 );
or ( n2571 , n2568 , n2570 );
and ( n2572 , n2571 , n2026 );
or ( n2573 , n2567 , n2572 );
not ( n2574 , n2573 );
and ( n2575 , n2574 , n1151 );
not ( n2576 , n2573 );
and ( n2577 , n719 , n2199 );
and ( n2578 , n2313 , n2213 );
xor ( n2579 , n2388 , n2391 );
and ( n2580 , n2579 , n2312 );
or ( n2581 , n2578 , n2580 );
and ( n2582 , n2581 , n2026 );
or ( n2583 , n2577 , n2582 );
not ( n2584 , n2583 );
and ( n2585 , n2584 , n1138 );
not ( n2586 , n2583 );
and ( n2587 , n720 , n2199 );
and ( n2588 , n2313 , n2207 );
xor ( n2589 , n2389 , n2390 );
and ( n2590 , n2589 , n2312 );
or ( n2591 , n2588 , n2590 );
and ( n2592 , n2591 , n2026 );
or ( n2593 , n2587 , n2592 );
not ( n2594 , n2593 );
and ( n2595 , n2594 , n1126 );
not ( n2596 , n2593 );
not ( n2597 , n2320 );
or ( n2598 , n1116 , n2597 );
and ( n2599 , n2596 , n2598 );
and ( n2600 , n1126 , n2598 );
or ( n2601 , n2595 , n2599 , n2600 );
and ( n2602 , n2586 , n2601 );
and ( n2603 , n1138 , n2601 );
or ( n2604 , n2585 , n2602 , n2603 );
and ( n2605 , n2576 , n2604 );
and ( n2606 , n1151 , n2604 );
or ( n2607 , n2575 , n2605 , n2606 );
and ( n2608 , n2566 , n2607 );
and ( n2609 , n1164 , n2607 );
or ( n2610 , n2565 , n2608 , n2609 );
and ( n2611 , n2556 , n2610 );
and ( n2612 , n1178 , n2610 );
or ( n2613 , n2555 , n2611 , n2612 );
and ( n2614 , n2546 , n2613 );
and ( n2615 , n1192 , n2613 );
or ( n2616 , n2545 , n2614 , n2615 );
and ( n2617 , n2536 , n2616 );
and ( n2618 , n1206 , n2616 );
or ( n2619 , n2535 , n2617 , n2618 );
and ( n2620 , n2526 , n2619 );
and ( n2621 , n1220 , n2619 );
or ( n2622 , n2525 , n2620 , n2621 );
and ( n2623 , n2516 , n2622 );
and ( n2624 , n1234 , n2622 );
or ( n2625 , n2515 , n2623 , n2624 );
and ( n2626 , n2506 , n2625 );
and ( n2627 , n1248 , n2625 );
or ( n2628 , n2505 , n2626 , n2627 );
and ( n2629 , n2496 , n2628 );
and ( n2630 , n1262 , n2628 );
or ( n2631 , n2495 , n2629 , n2630 );
and ( n2632 , n2486 , n2631 );
and ( n2633 , n1276 , n2631 );
or ( n2634 , n2485 , n2632 , n2633 );
and ( n2635 , n2476 , n2634 );
and ( n2636 , n1290 , n2634 );
or ( n2637 , n2475 , n2635 , n2636 );
and ( n2638 , n2466 , n2637 );
and ( n2639 , n1304 , n2637 );
or ( n2640 , n2465 , n2638 , n2639 );
and ( n2641 , n2456 , n2640 );
and ( n2642 , n1318 , n2640 );
or ( n2643 , n2455 , n2641 , n2642 );
and ( n2644 , n2446 , n2643 );
and ( n2645 , n1332 , n2643 );
or ( n2646 , n2445 , n2644 , n2645 );
and ( n2647 , n2436 , n2646 );
and ( n2648 , n1346 , n2646 );
or ( n2649 , n2435 , n2647 , n2648 );
and ( n2650 , n2426 , n2649 );
and ( n2651 , n1360 , n2649 );
or ( n2652 , n2425 , n2650 , n2651 );
and ( n2653 , n2416 , n2652 );
and ( n2654 , n1374 , n2652 );
or ( n2655 , n2415 , n2653 , n2654 );
and ( n2656 , n2368 , n2655 );
and ( n2657 , n1388 , n2655 );
or ( n2658 , n2367 , n2656 , n2657 );
and ( n2659 , n2364 , n2658 );
and ( n2660 , n1402 , n2658 );
or ( n2661 , n2363 , n2659 , n2660 );
and ( n2662 , n2360 , n2661 );
and ( n2663 , n1416 , n2661 );
or ( n2664 , n2359 , n2662 , n2663 );
and ( n2665 , n2356 , n2664 );
and ( n2666 , n1430 , n2664 );
or ( n2667 , n2355 , n2665 , n2666 );
and ( n2668 , n2352 , n2667 );
and ( n2669 , n1444 , n2667 );
or ( n2670 , n2351 , n2668 , n2669 );
and ( n2671 , n2348 , n2670 );
and ( n2672 , n1458 , n2670 );
or ( n2673 , n2347 , n2671 , n2672 );
and ( n2674 , n2344 , n2673 );
and ( n2675 , n1472 , n2673 );
or ( n2676 , n2343 , n2674 , n2675 );
and ( n2677 , n2340 , n2676 );
and ( n2678 , n1486 , n2676 );
or ( n2679 , n2339 , n2677 , n2678 );
and ( n2680 , n2336 , n2679 );
and ( n2681 , n1500 , n2679 );
or ( n2682 , n2335 , n2680 , n2681 );
and ( n2683 , n2332 , n2682 );
and ( n2684 , n1632 , n2682 );
or ( n2685 , n2331 , n2683 , n2684 );
and ( n2686 , n2328 , n2685 );
and ( n2687 , n1625 , n2685 );
or ( n2688 , n2327 , n2686 , n2687 );
xor ( n2689 , n2324 , n2688 );
not ( n2690 , n2689 );
xor ( n2691 , n1126 , n2596 );
xor ( n2692 , n2691 , n2598 );
and ( n2693 , n2690 , n2692 );
not ( n2694 , n2692 );
not ( n2695 , n2321 );
xor ( n2696 , n2694 , n2695 );
and ( n2697 , n2696 , n2689 );
or ( n2698 , n2693 , n2697 );
or ( n2699 , n2321 , n2698 );
xor ( n2700 , n1138 , n2586 );
xor ( n2701 , n2700 , n2601 );
and ( n2702 , n2690 , n2701 );
not ( n2703 , n2701 );
and ( n2704 , n2694 , n2695 );
xor ( n2705 , n2703 , n2704 );
and ( n2706 , n2705 , n2689 );
or ( n2707 , n2702 , n2706 );
or ( n2708 , n2699 , n2707 );
xor ( n2709 , n1151 , n2576 );
xor ( n2710 , n2709 , n2604 );
and ( n2711 , n2690 , n2710 );
not ( n2712 , n2710 );
and ( n2713 , n2703 , n2704 );
xor ( n2714 , n2712 , n2713 );
and ( n2715 , n2714 , n2689 );
or ( n2716 , n2711 , n2715 );
or ( n2717 , n2708 , n2716 );
xor ( n2718 , n1164 , n2566 );
xor ( n2719 , n2718 , n2607 );
and ( n2720 , n2690 , n2719 );
not ( n2721 , n2719 );
and ( n2722 , n2712 , n2713 );
xor ( n2723 , n2721 , n2722 );
and ( n2724 , n2723 , n2689 );
or ( n2725 , n2720 , n2724 );
or ( n2726 , n2717 , n2725 );
xor ( n2727 , n1178 , n2556 );
xor ( n2728 , n2727 , n2610 );
and ( n2729 , n2690 , n2728 );
not ( n2730 , n2728 );
and ( n2731 , n2721 , n2722 );
xor ( n2732 , n2730 , n2731 );
and ( n2733 , n2732 , n2689 );
or ( n2734 , n2729 , n2733 );
or ( n2735 , n2726 , n2734 );
xor ( n2736 , n1192 , n2546 );
xor ( n2737 , n2736 , n2613 );
and ( n2738 , n2690 , n2737 );
not ( n2739 , n2737 );
and ( n2740 , n2730 , n2731 );
xor ( n2741 , n2739 , n2740 );
and ( n2742 , n2741 , n2689 );
or ( n2743 , n2738 , n2742 );
or ( n2744 , n2735 , n2743 );
xor ( n2745 , n1206 , n2536 );
xor ( n2746 , n2745 , n2616 );
and ( n2747 , n2690 , n2746 );
not ( n2748 , n2746 );
and ( n2749 , n2739 , n2740 );
xor ( n2750 , n2748 , n2749 );
and ( n2751 , n2750 , n2689 );
or ( n2752 , n2747 , n2751 );
or ( n2753 , n2744 , n2752 );
xor ( n2754 , n1220 , n2526 );
xor ( n2755 , n2754 , n2619 );
and ( n2756 , n2690 , n2755 );
not ( n2757 , n2755 );
and ( n2758 , n2748 , n2749 );
xor ( n2759 , n2757 , n2758 );
and ( n2760 , n2759 , n2689 );
or ( n2761 , n2756 , n2760 );
or ( n2762 , n2753 , n2761 );
xor ( n2763 , n1234 , n2516 );
xor ( n2764 , n2763 , n2622 );
and ( n2765 , n2690 , n2764 );
not ( n2766 , n2764 );
and ( n2767 , n2757 , n2758 );
xor ( n2768 , n2766 , n2767 );
and ( n2769 , n2768 , n2689 );
or ( n2770 , n2765 , n2769 );
or ( n2771 , n2762 , n2770 );
xor ( n2772 , n1248 , n2506 );
xor ( n2773 , n2772 , n2625 );
and ( n2774 , n2690 , n2773 );
not ( n2775 , n2773 );
and ( n2776 , n2766 , n2767 );
xor ( n2777 , n2775 , n2776 );
and ( n2778 , n2777 , n2689 );
or ( n2779 , n2774 , n2778 );
or ( n2780 , n2771 , n2779 );
xor ( n2781 , n1262 , n2496 );
xor ( n2782 , n2781 , n2628 );
and ( n2783 , n2690 , n2782 );
not ( n2784 , n2782 );
and ( n2785 , n2775 , n2776 );
xor ( n2786 , n2784 , n2785 );
and ( n2787 , n2786 , n2689 );
or ( n2788 , n2783 , n2787 );
or ( n2789 , n2780 , n2788 );
xor ( n2790 , n1276 , n2486 );
xor ( n2791 , n2790 , n2631 );
and ( n2792 , n2690 , n2791 );
not ( n2793 , n2791 );
and ( n2794 , n2784 , n2785 );
xor ( n2795 , n2793 , n2794 );
and ( n2796 , n2795 , n2689 );
or ( n2797 , n2792 , n2796 );
or ( n2798 , n2789 , n2797 );
xor ( n2799 , n1290 , n2476 );
xor ( n2800 , n2799 , n2634 );
and ( n2801 , n2690 , n2800 );
not ( n2802 , n2800 );
and ( n2803 , n2793 , n2794 );
xor ( n2804 , n2802 , n2803 );
and ( n2805 , n2804 , n2689 );
or ( n2806 , n2801 , n2805 );
or ( n2807 , n2798 , n2806 );
xor ( n2808 , n1304 , n2466 );
xor ( n2809 , n2808 , n2637 );
and ( n2810 , n2690 , n2809 );
not ( n2811 , n2809 );
and ( n2812 , n2802 , n2803 );
xor ( n2813 , n2811 , n2812 );
and ( n2814 , n2813 , n2689 );
or ( n2815 , n2810 , n2814 );
or ( n2816 , n2807 , n2815 );
xor ( n2817 , n1318 , n2456 );
xor ( n2818 , n2817 , n2640 );
and ( n2819 , n2690 , n2818 );
not ( n2820 , n2818 );
and ( n2821 , n2811 , n2812 );
xor ( n2822 , n2820 , n2821 );
and ( n2823 , n2822 , n2689 );
or ( n2824 , n2819 , n2823 );
or ( n2825 , n2816 , n2824 );
xor ( n2826 , n1332 , n2446 );
xor ( n2827 , n2826 , n2643 );
and ( n2828 , n2690 , n2827 );
not ( n2829 , n2827 );
and ( n2830 , n2820 , n2821 );
xor ( n2831 , n2829 , n2830 );
and ( n2832 , n2831 , n2689 );
or ( n2833 , n2828 , n2832 );
or ( n2834 , n2825 , n2833 );
xor ( n2835 , n1346 , n2436 );
xor ( n2836 , n2835 , n2646 );
and ( n2837 , n2690 , n2836 );
not ( n2838 , n2836 );
and ( n2839 , n2829 , n2830 );
xor ( n2840 , n2838 , n2839 );
and ( n2841 , n2840 , n2689 );
or ( n2842 , n2837 , n2841 );
or ( n2843 , n2834 , n2842 );
xor ( n2844 , n1360 , n2426 );
xor ( n2845 , n2844 , n2649 );
and ( n2846 , n2690 , n2845 );
not ( n2847 , n2845 );
and ( n2848 , n2838 , n2839 );
xor ( n2849 , n2847 , n2848 );
and ( n2850 , n2849 , n2689 );
or ( n2851 , n2846 , n2850 );
or ( n2852 , n2843 , n2851 );
xor ( n2853 , n1374 , n2416 );
xor ( n2854 , n2853 , n2652 );
and ( n2855 , n2690 , n2854 );
not ( n2856 , n2854 );
and ( n2857 , n2847 , n2848 );
xor ( n2858 , n2856 , n2857 );
and ( n2859 , n2858 , n2689 );
or ( n2860 , n2855 , n2859 );
or ( n2861 , n2852 , n2860 );
xor ( n2862 , n1388 , n2368 );
xor ( n2863 , n2862 , n2655 );
and ( n2864 , n2690 , n2863 );
not ( n2865 , n2863 );
and ( n2866 , n2856 , n2857 );
xor ( n2867 , n2865 , n2866 );
and ( n2868 , n2867 , n2689 );
or ( n2869 , n2864 , n2868 );
or ( n2870 , n2861 , n2869 );
xor ( n2871 , n1402 , n2364 );
xor ( n2872 , n2871 , n2658 );
and ( n2873 , n2690 , n2872 );
not ( n2874 , n2872 );
and ( n2875 , n2865 , n2866 );
xor ( n2876 , n2874 , n2875 );
and ( n2877 , n2876 , n2689 );
or ( n2878 , n2873 , n2877 );
or ( n2879 , n2870 , n2878 );
xor ( n2880 , n1416 , n2360 );
xor ( n2881 , n2880 , n2661 );
and ( n2882 , n2690 , n2881 );
not ( n2883 , n2881 );
and ( n2884 , n2874 , n2875 );
xor ( n2885 , n2883 , n2884 );
and ( n2886 , n2885 , n2689 );
or ( n2887 , n2882 , n2886 );
or ( n2888 , n2879 , n2887 );
xor ( n2889 , n1430 , n2356 );
xor ( n2890 , n2889 , n2664 );
and ( n2891 , n2690 , n2890 );
not ( n2892 , n2890 );
and ( n2893 , n2883 , n2884 );
xor ( n2894 , n2892 , n2893 );
and ( n2895 , n2894 , n2689 );
or ( n2896 , n2891 , n2895 );
or ( n2897 , n2888 , n2896 );
xor ( n2898 , n1444 , n2352 );
xor ( n2899 , n2898 , n2667 );
and ( n2900 , n2690 , n2899 );
not ( n2901 , n2899 );
and ( n2902 , n2892 , n2893 );
xor ( n2903 , n2901 , n2902 );
and ( n2904 , n2903 , n2689 );
or ( n2905 , n2900 , n2904 );
or ( n2906 , n2897 , n2905 );
xor ( n2907 , n1458 , n2348 );
xor ( n2908 , n2907 , n2670 );
and ( n2909 , n2690 , n2908 );
not ( n2910 , n2908 );
and ( n2911 , n2901 , n2902 );
xor ( n2912 , n2910 , n2911 );
and ( n2913 , n2912 , n2689 );
or ( n2914 , n2909 , n2913 );
or ( n2915 , n2906 , n2914 );
xor ( n2916 , n1472 , n2344 );
xor ( n2917 , n2916 , n2673 );
and ( n2918 , n2690 , n2917 );
not ( n2919 , n2917 );
and ( n2920 , n2910 , n2911 );
xor ( n2921 , n2919 , n2920 );
and ( n2922 , n2921 , n2689 );
or ( n2923 , n2918 , n2922 );
or ( n2924 , n2915 , n2923 );
xor ( n2925 , n1486 , n2340 );
xor ( n2926 , n2925 , n2676 );
and ( n2927 , n2690 , n2926 );
not ( n2928 , n2926 );
and ( n2929 , n2919 , n2920 );
xor ( n2930 , n2928 , n2929 );
and ( n2931 , n2930 , n2689 );
or ( n2932 , n2927 , n2931 );
or ( n2933 , n2924 , n2932 );
xor ( n2934 , n1500 , n2336 );
xor ( n2935 , n2934 , n2679 );
and ( n2936 , n2690 , n2935 );
not ( n2937 , n2935 );
and ( n2938 , n2928 , n2929 );
xor ( n2939 , n2937 , n2938 );
and ( n2940 , n2939 , n2689 );
or ( n2941 , n2936 , n2940 );
or ( n2942 , n2933 , n2941 );
xor ( n2943 , n1632 , n2332 );
xor ( n2944 , n2943 , n2682 );
and ( n2945 , n2690 , n2944 );
not ( n2946 , n2944 );
and ( n2947 , n2937 , n2938 );
xor ( n2948 , n2946 , n2947 );
and ( n2949 , n2948 , n2689 );
or ( n2950 , n2945 , n2949 );
or ( n2951 , n2942 , n2950 );
and ( n2952 , n2951 , n2689 );
not ( n2953 , n2952 );
and ( n2954 , n2953 , n2824 );
xor ( n2955 , n2824 , n2689 );
xor ( n2956 , n2815 , n2689 );
xor ( n2957 , n2806 , n2689 );
xor ( n2958 , n2797 , n2689 );
xor ( n2959 , n2788 , n2689 );
xor ( n2960 , n2779 , n2689 );
xor ( n2961 , n2770 , n2689 );
xor ( n2962 , n2761 , n2689 );
xor ( n2963 , n2752 , n2689 );
xor ( n2964 , n2743 , n2689 );
xor ( n2965 , n2734 , n2689 );
xor ( n2966 , n2725 , n2689 );
xor ( n2967 , n2716 , n2689 );
xor ( n2968 , n2707 , n2689 );
xor ( n2969 , n2698 , n2689 );
xor ( n2970 , n2321 , n2689 );
and ( n2971 , n2970 , n2689 );
and ( n2972 , n2969 , n2971 );
and ( n2973 , n2968 , n2972 );
and ( n2974 , n2967 , n2973 );
and ( n2975 , n2966 , n2974 );
and ( n2976 , n2965 , n2975 );
and ( n2977 , n2964 , n2976 );
and ( n2978 , n2963 , n2977 );
and ( n2979 , n2962 , n2978 );
and ( n2980 , n2961 , n2979 );
and ( n2981 , n2960 , n2980 );
and ( n2982 , n2959 , n2981 );
and ( n2983 , n2958 , n2982 );
and ( n2984 , n2957 , n2983 );
and ( n2985 , n2956 , n2984 );
xor ( n2986 , n2955 , n2985 );
and ( n2987 , n2986 , n2952 );
or ( n2988 , n2954 , n2987 );
and ( n2989 , n2988 , n2084 );
or ( n2990 , n2989 , n2092 );
not ( n2991 , n2195 );
and ( n2992 , n2176 , n2182 , n2189 , n2991 );
and ( n2993 , n2175 , n2182 , n2189 , n2991 );
or ( n2994 , n2992 , n2993 );
nor ( n2995 , n2176 , n2182 , n2189 , n2991 );
or ( n2996 , n2994 , n2995 );
nor ( n2997 , n2176 , n2183 , n2189 , n2991 );
or ( n2998 , n2996 , n2997 );
and ( n2999 , n2990 , n2998 );
xor ( n3000 , n1120 , n2322 );
and ( n3001 , n1625 , n2325 );
and ( n3002 , n1632 , n2329 );
and ( n3003 , n1500 , n2333 );
and ( n3004 , n1486 , n2337 );
and ( n3005 , n1472 , n2341 );
and ( n3006 , n1458 , n2345 );
and ( n3007 , n1444 , n2349 );
and ( n3008 , n1430 , n2353 );
and ( n3009 , n1416 , n2357 );
and ( n3010 , n1402 , n2361 );
and ( n3011 , n1388 , n2365 );
and ( n3012 , n1374 , n2413 );
and ( n3013 , n1360 , n2423 );
and ( n3014 , n1346 , n2433 );
and ( n3015 , n1332 , n2443 );
and ( n3016 , n1318 , n2453 );
and ( n3017 , n1304 , n2463 );
and ( n3018 , n1290 , n2473 );
and ( n3019 , n1276 , n2483 );
and ( n3020 , n1262 , n2493 );
and ( n3021 , n1248 , n2503 );
and ( n3022 , n1234 , n2513 );
and ( n3023 , n1220 , n2523 );
and ( n3024 , n1206 , n2533 );
and ( n3025 , n1192 , n2543 );
and ( n3026 , n1178 , n2553 );
and ( n3027 , n1164 , n2563 );
and ( n3028 , n1151 , n2573 );
and ( n3029 , n1138 , n2583 );
and ( n3030 , n1126 , n2593 );
and ( n3031 , n1116 , n2320 );
and ( n3032 , n2593 , n3031 );
and ( n3033 , n1126 , n3031 );
or ( n3034 , n3030 , n3032 , n3033 );
and ( n3035 , n2583 , n3034 );
and ( n3036 , n1138 , n3034 );
or ( n3037 , n3029 , n3035 , n3036 );
and ( n3038 , n2573 , n3037 );
and ( n3039 , n1151 , n3037 );
or ( n3040 , n3028 , n3038 , n3039 );
and ( n3041 , n2563 , n3040 );
and ( n3042 , n1164 , n3040 );
or ( n3043 , n3027 , n3041 , n3042 );
and ( n3044 , n2553 , n3043 );
and ( n3045 , n1178 , n3043 );
or ( n3046 , n3026 , n3044 , n3045 );
and ( n3047 , n2543 , n3046 );
and ( n3048 , n1192 , n3046 );
or ( n3049 , n3025 , n3047 , n3048 );
and ( n3050 , n2533 , n3049 );
and ( n3051 , n1206 , n3049 );
or ( n3052 , n3024 , n3050 , n3051 );
and ( n3053 , n2523 , n3052 );
and ( n3054 , n1220 , n3052 );
or ( n3055 , n3023 , n3053 , n3054 );
and ( n3056 , n2513 , n3055 );
and ( n3057 , n1234 , n3055 );
or ( n3058 , n3022 , n3056 , n3057 );
and ( n3059 , n2503 , n3058 );
and ( n3060 , n1248 , n3058 );
or ( n3061 , n3021 , n3059 , n3060 );
and ( n3062 , n2493 , n3061 );
and ( n3063 , n1262 , n3061 );
or ( n3064 , n3020 , n3062 , n3063 );
and ( n3065 , n2483 , n3064 );
and ( n3066 , n1276 , n3064 );
or ( n3067 , n3019 , n3065 , n3066 );
and ( n3068 , n2473 , n3067 );
and ( n3069 , n1290 , n3067 );
or ( n3070 , n3018 , n3068 , n3069 );
and ( n3071 , n2463 , n3070 );
and ( n3072 , n1304 , n3070 );
or ( n3073 , n3017 , n3071 , n3072 );
and ( n3074 , n2453 , n3073 );
and ( n3075 , n1318 , n3073 );
or ( n3076 , n3016 , n3074 , n3075 );
and ( n3077 , n2443 , n3076 );
and ( n3078 , n1332 , n3076 );
or ( n3079 , n3015 , n3077 , n3078 );
and ( n3080 , n2433 , n3079 );
and ( n3081 , n1346 , n3079 );
or ( n3082 , n3014 , n3080 , n3081 );
and ( n3083 , n2423 , n3082 );
and ( n3084 , n1360 , n3082 );
or ( n3085 , n3013 , n3083 , n3084 );
and ( n3086 , n2413 , n3085 );
and ( n3087 , n1374 , n3085 );
or ( n3088 , n3012 , n3086 , n3087 );
and ( n3089 , n2365 , n3088 );
and ( n3090 , n1388 , n3088 );
or ( n3091 , n3011 , n3089 , n3090 );
and ( n3092 , n2361 , n3091 );
and ( n3093 , n1402 , n3091 );
or ( n3094 , n3010 , n3092 , n3093 );
and ( n3095 , n2357 , n3094 );
and ( n3096 , n1416 , n3094 );
or ( n3097 , n3009 , n3095 , n3096 );
and ( n3098 , n2353 , n3097 );
and ( n3099 , n1430 , n3097 );
or ( n3100 , n3008 , n3098 , n3099 );
and ( n3101 , n2349 , n3100 );
and ( n3102 , n1444 , n3100 );
or ( n3103 , n3007 , n3101 , n3102 );
and ( n3104 , n2345 , n3103 );
and ( n3105 , n1458 , n3103 );
or ( n3106 , n3006 , n3104 , n3105 );
and ( n3107 , n2341 , n3106 );
and ( n3108 , n1472 , n3106 );
or ( n3109 , n3005 , n3107 , n3108 );
and ( n3110 , n2337 , n3109 );
and ( n3111 , n1486 , n3109 );
or ( n3112 , n3004 , n3110 , n3111 );
and ( n3113 , n2333 , n3112 );
and ( n3114 , n1500 , n3112 );
or ( n3115 , n3003 , n3113 , n3114 );
and ( n3116 , n2329 , n3115 );
and ( n3117 , n1632 , n3115 );
or ( n3118 , n3002 , n3116 , n3117 );
and ( n3119 , n2325 , n3118 );
and ( n3120 , n1625 , n3118 );
or ( n3121 , n3001 , n3119 , n3120 );
xor ( n3122 , n3000 , n3121 );
not ( n3123 , n3122 );
xor ( n3124 , n1126 , n2593 );
xor ( n3125 , n3124 , n3031 );
and ( n3126 , n3123 , n3125 );
not ( n3127 , n3125 );
xor ( n3128 , n3127 , n2695 );
and ( n3129 , n3128 , n3122 );
or ( n3130 , n3126 , n3129 );
or ( n3131 , n2321 , n3130 );
xor ( n3132 , n1138 , n2583 );
xor ( n3133 , n3132 , n3034 );
and ( n3134 , n3123 , n3133 );
not ( n3135 , n3133 );
and ( n3136 , n3127 , n2695 );
xor ( n3137 , n3135 , n3136 );
and ( n3138 , n3137 , n3122 );
or ( n3139 , n3134 , n3138 );
or ( n3140 , n3131 , n3139 );
xor ( n3141 , n1151 , n2573 );
xor ( n3142 , n3141 , n3037 );
and ( n3143 , n3123 , n3142 );
not ( n3144 , n3142 );
and ( n3145 , n3135 , n3136 );
xor ( n3146 , n3144 , n3145 );
and ( n3147 , n3146 , n3122 );
or ( n3148 , n3143 , n3147 );
or ( n3149 , n3140 , n3148 );
xor ( n3150 , n1164 , n2563 );
xor ( n3151 , n3150 , n3040 );
and ( n3152 , n3123 , n3151 );
not ( n3153 , n3151 );
and ( n3154 , n3144 , n3145 );
xor ( n3155 , n3153 , n3154 );
and ( n3156 , n3155 , n3122 );
or ( n3157 , n3152 , n3156 );
or ( n3158 , n3149 , n3157 );
xor ( n3159 , n1178 , n2553 );
xor ( n3160 , n3159 , n3043 );
and ( n3161 , n3123 , n3160 );
not ( n3162 , n3160 );
and ( n3163 , n3153 , n3154 );
xor ( n3164 , n3162 , n3163 );
and ( n3165 , n3164 , n3122 );
or ( n3166 , n3161 , n3165 );
or ( n3167 , n3158 , n3166 );
xor ( n3168 , n1192 , n2543 );
xor ( n3169 , n3168 , n3046 );
and ( n3170 , n3123 , n3169 );
not ( n3171 , n3169 );
and ( n3172 , n3162 , n3163 );
xor ( n3173 , n3171 , n3172 );
and ( n3174 , n3173 , n3122 );
or ( n3175 , n3170 , n3174 );
or ( n3176 , n3167 , n3175 );
xor ( n3177 , n1206 , n2533 );
xor ( n3178 , n3177 , n3049 );
and ( n3179 , n3123 , n3178 );
not ( n3180 , n3178 );
and ( n3181 , n3171 , n3172 );
xor ( n3182 , n3180 , n3181 );
and ( n3183 , n3182 , n3122 );
or ( n3184 , n3179 , n3183 );
or ( n3185 , n3176 , n3184 );
xor ( n3186 , n1220 , n2523 );
xor ( n3187 , n3186 , n3052 );
and ( n3188 , n3123 , n3187 );
not ( n3189 , n3187 );
and ( n3190 , n3180 , n3181 );
xor ( n3191 , n3189 , n3190 );
and ( n3192 , n3191 , n3122 );
or ( n3193 , n3188 , n3192 );
or ( n3194 , n3185 , n3193 );
xor ( n3195 , n1234 , n2513 );
xor ( n3196 , n3195 , n3055 );
and ( n3197 , n3123 , n3196 );
not ( n3198 , n3196 );
and ( n3199 , n3189 , n3190 );
xor ( n3200 , n3198 , n3199 );
and ( n3201 , n3200 , n3122 );
or ( n3202 , n3197 , n3201 );
or ( n3203 , n3194 , n3202 );
xor ( n3204 , n1248 , n2503 );
xor ( n3205 , n3204 , n3058 );
and ( n3206 , n3123 , n3205 );
not ( n3207 , n3205 );
and ( n3208 , n3198 , n3199 );
xor ( n3209 , n3207 , n3208 );
and ( n3210 , n3209 , n3122 );
or ( n3211 , n3206 , n3210 );
or ( n3212 , n3203 , n3211 );
xor ( n3213 , n1262 , n2493 );
xor ( n3214 , n3213 , n3061 );
and ( n3215 , n3123 , n3214 );
not ( n3216 , n3214 );
and ( n3217 , n3207 , n3208 );
xor ( n3218 , n3216 , n3217 );
and ( n3219 , n3218 , n3122 );
or ( n3220 , n3215 , n3219 );
or ( n3221 , n3212 , n3220 );
xor ( n3222 , n1276 , n2483 );
xor ( n3223 , n3222 , n3064 );
and ( n3224 , n3123 , n3223 );
not ( n3225 , n3223 );
and ( n3226 , n3216 , n3217 );
xor ( n3227 , n3225 , n3226 );
and ( n3228 , n3227 , n3122 );
or ( n3229 , n3224 , n3228 );
or ( n3230 , n3221 , n3229 );
xor ( n3231 , n1290 , n2473 );
xor ( n3232 , n3231 , n3067 );
and ( n3233 , n3123 , n3232 );
not ( n3234 , n3232 );
and ( n3235 , n3225 , n3226 );
xor ( n3236 , n3234 , n3235 );
and ( n3237 , n3236 , n3122 );
or ( n3238 , n3233 , n3237 );
or ( n3239 , n3230 , n3238 );
xor ( n3240 , n1304 , n2463 );
xor ( n3241 , n3240 , n3070 );
and ( n3242 , n3123 , n3241 );
not ( n3243 , n3241 );
and ( n3244 , n3234 , n3235 );
xor ( n3245 , n3243 , n3244 );
and ( n3246 , n3245 , n3122 );
or ( n3247 , n3242 , n3246 );
or ( n3248 , n3239 , n3247 );
xor ( n3249 , n1318 , n2453 );
xor ( n3250 , n3249 , n3073 );
and ( n3251 , n3123 , n3250 );
not ( n3252 , n3250 );
and ( n3253 , n3243 , n3244 );
xor ( n3254 , n3252 , n3253 );
and ( n3255 , n3254 , n3122 );
or ( n3256 , n3251 , n3255 );
or ( n3257 , n3248 , n3256 );
xor ( n3258 , n1332 , n2443 );
xor ( n3259 , n3258 , n3076 );
and ( n3260 , n3123 , n3259 );
not ( n3261 , n3259 );
and ( n3262 , n3252 , n3253 );
xor ( n3263 , n3261 , n3262 );
and ( n3264 , n3263 , n3122 );
or ( n3265 , n3260 , n3264 );
or ( n3266 , n3257 , n3265 );
xor ( n3267 , n1346 , n2433 );
xor ( n3268 , n3267 , n3079 );
and ( n3269 , n3123 , n3268 );
not ( n3270 , n3268 );
and ( n3271 , n3261 , n3262 );
xor ( n3272 , n3270 , n3271 );
and ( n3273 , n3272 , n3122 );
or ( n3274 , n3269 , n3273 );
or ( n3275 , n3266 , n3274 );
xor ( n3276 , n1360 , n2423 );
xor ( n3277 , n3276 , n3082 );
and ( n3278 , n3123 , n3277 );
not ( n3279 , n3277 );
and ( n3280 , n3270 , n3271 );
xor ( n3281 , n3279 , n3280 );
and ( n3282 , n3281 , n3122 );
or ( n3283 , n3278 , n3282 );
or ( n3284 , n3275 , n3283 );
xor ( n3285 , n1374 , n2413 );
xor ( n3286 , n3285 , n3085 );
and ( n3287 , n3123 , n3286 );
not ( n3288 , n3286 );
and ( n3289 , n3279 , n3280 );
xor ( n3290 , n3288 , n3289 );
and ( n3291 , n3290 , n3122 );
or ( n3292 , n3287 , n3291 );
or ( n3293 , n3284 , n3292 );
xor ( n3294 , n1388 , n2365 );
xor ( n3295 , n3294 , n3088 );
and ( n3296 , n3123 , n3295 );
not ( n3297 , n3295 );
and ( n3298 , n3288 , n3289 );
xor ( n3299 , n3297 , n3298 );
and ( n3300 , n3299 , n3122 );
or ( n3301 , n3296 , n3300 );
or ( n3302 , n3293 , n3301 );
xor ( n3303 , n1402 , n2361 );
xor ( n3304 , n3303 , n3091 );
and ( n3305 , n3123 , n3304 );
not ( n3306 , n3304 );
and ( n3307 , n3297 , n3298 );
xor ( n3308 , n3306 , n3307 );
and ( n3309 , n3308 , n3122 );
or ( n3310 , n3305 , n3309 );
or ( n3311 , n3302 , n3310 );
xor ( n3312 , n1416 , n2357 );
xor ( n3313 , n3312 , n3094 );
and ( n3314 , n3123 , n3313 );
not ( n3315 , n3313 );
and ( n3316 , n3306 , n3307 );
xor ( n3317 , n3315 , n3316 );
and ( n3318 , n3317 , n3122 );
or ( n3319 , n3314 , n3318 );
or ( n3320 , n3311 , n3319 );
xor ( n3321 , n1430 , n2353 );
xor ( n3322 , n3321 , n3097 );
and ( n3323 , n3123 , n3322 );
not ( n3324 , n3322 );
and ( n3325 , n3315 , n3316 );
xor ( n3326 , n3324 , n3325 );
and ( n3327 , n3326 , n3122 );
or ( n3328 , n3323 , n3327 );
or ( n3329 , n3320 , n3328 );
xor ( n3330 , n1444 , n2349 );
xor ( n3331 , n3330 , n3100 );
and ( n3332 , n3123 , n3331 );
not ( n3333 , n3331 );
and ( n3334 , n3324 , n3325 );
xor ( n3335 , n3333 , n3334 );
and ( n3336 , n3335 , n3122 );
or ( n3337 , n3332 , n3336 );
or ( n3338 , n3329 , n3337 );
xor ( n3339 , n1458 , n2345 );
xor ( n3340 , n3339 , n3103 );
and ( n3341 , n3123 , n3340 );
not ( n3342 , n3340 );
and ( n3343 , n3333 , n3334 );
xor ( n3344 , n3342 , n3343 );
and ( n3345 , n3344 , n3122 );
or ( n3346 , n3341 , n3345 );
or ( n3347 , n3338 , n3346 );
xor ( n3348 , n1472 , n2341 );
xor ( n3349 , n3348 , n3106 );
and ( n3350 , n3123 , n3349 );
not ( n3351 , n3349 );
and ( n3352 , n3342 , n3343 );
xor ( n3353 , n3351 , n3352 );
and ( n3354 , n3353 , n3122 );
or ( n3355 , n3350 , n3354 );
or ( n3356 , n3347 , n3355 );
xor ( n3357 , n1486 , n2337 );
xor ( n3358 , n3357 , n3109 );
and ( n3359 , n3123 , n3358 );
not ( n3360 , n3358 );
and ( n3361 , n3351 , n3352 );
xor ( n3362 , n3360 , n3361 );
and ( n3363 , n3362 , n3122 );
or ( n3364 , n3359 , n3363 );
or ( n3365 , n3356 , n3364 );
xor ( n3366 , n1500 , n2333 );
xor ( n3367 , n3366 , n3112 );
and ( n3368 , n3123 , n3367 );
not ( n3369 , n3367 );
and ( n3370 , n3360 , n3361 );
xor ( n3371 , n3369 , n3370 );
and ( n3372 , n3371 , n3122 );
or ( n3373 , n3368 , n3372 );
or ( n3374 , n3365 , n3373 );
xor ( n3375 , n1632 , n2329 );
xor ( n3376 , n3375 , n3115 );
and ( n3377 , n3123 , n3376 );
not ( n3378 , n3376 );
and ( n3379 , n3369 , n3370 );
xor ( n3380 , n3378 , n3379 );
and ( n3381 , n3380 , n3122 );
or ( n3382 , n3377 , n3381 );
or ( n3383 , n3374 , n3382 );
and ( n3384 , n3383 , n3122 );
not ( n3385 , n3384 );
and ( n3386 , n3385 , n3256 );
xor ( n3387 , n3256 , n3122 );
xor ( n3388 , n3247 , n3122 );
xor ( n3389 , n3238 , n3122 );
xor ( n3390 , n3229 , n3122 );
xor ( n3391 , n3220 , n3122 );
xor ( n3392 , n3211 , n3122 );
xor ( n3393 , n3202 , n3122 );
xor ( n3394 , n3193 , n3122 );
xor ( n3395 , n3184 , n3122 );
xor ( n3396 , n3175 , n3122 );
xor ( n3397 , n3166 , n3122 );
xor ( n3398 , n3157 , n3122 );
xor ( n3399 , n3148 , n3122 );
xor ( n3400 , n3139 , n3122 );
xor ( n3401 , n3130 , n3122 );
xor ( n3402 , n2321 , n3122 );
and ( n3403 , n3402 , n3122 );
and ( n3404 , n3401 , n3403 );
and ( n3405 , n3400 , n3404 );
and ( n3406 , n3399 , n3405 );
and ( n3407 , n3398 , n3406 );
and ( n3408 , n3397 , n3407 );
and ( n3409 , n3396 , n3408 );
and ( n3410 , n3395 , n3409 );
and ( n3411 , n3394 , n3410 );
and ( n3412 , n3393 , n3411 );
and ( n3413 , n3392 , n3412 );
and ( n3414 , n3391 , n3413 );
and ( n3415 , n3390 , n3414 );
and ( n3416 , n3389 , n3415 );
and ( n3417 , n3388 , n3416 );
xor ( n3418 , n3387 , n3417 );
and ( n3419 , n3418 , n3384 );
or ( n3420 , n3386 , n3419 );
and ( n3421 , n3420 , n2084 );
or ( n3422 , n3421 , n2092 );
and ( n3423 , n2176 , n2183 , n2189 , n2991 );
and ( n3424 , n2175 , n2183 , n2189 , n2991 );
or ( n3425 , n3423 , n3424 );
nor ( n3426 , n2175 , n2182 , n2189 , n2991 );
or ( n3427 , n3425 , n3426 );
nor ( n3428 , n2175 , n2183 , n2189 , n2991 );
or ( n3429 , n3427 , n3428 );
and ( n3430 , n3422 , n3429 );
and ( n3431 , n2453 , n2084 );
or ( n3432 , n3431 , n2092 );
nor ( n3433 , n2175 , n2183 , n2189 , n2195 );
nor ( n3434 , n2176 , n2183 , n2189 , n2195 );
or ( n3435 , n3433 , n3434 );
and ( n3436 , n3432 , n3435 );
not ( n3437 , n2453 );
not ( n3438 , n2463 );
not ( n3439 , n2473 );
not ( n3440 , n2483 );
not ( n3441 , n2493 );
not ( n3442 , n2503 );
not ( n3443 , n2513 );
not ( n3444 , n2523 );
not ( n3445 , n2533 );
not ( n3446 , n2543 );
not ( n3447 , n2553 );
not ( n3448 , n2563 );
not ( n3449 , n2573 );
not ( n3450 , n2583 );
not ( n3451 , n2593 );
not ( n3452 , n2320 );
and ( n3453 , n3451 , n3452 );
and ( n3454 , n3450 , n3453 );
and ( n3455 , n3449 , n3454 );
and ( n3456 , n3448 , n3455 );
and ( n3457 , n3447 , n3456 );
and ( n3458 , n3446 , n3457 );
and ( n3459 , n3445 , n3458 );
and ( n3460 , n3444 , n3459 );
and ( n3461 , n3443 , n3460 );
and ( n3462 , n3442 , n3461 );
and ( n3463 , n3441 , n3462 );
and ( n3464 , n3440 , n3463 );
and ( n3465 , n3439 , n3464 );
and ( n3466 , n3438 , n3465 );
xor ( n3467 , n3437 , n3466 );
and ( n3468 , n3467 , n2084 );
or ( n3469 , n3468 , n2092 );
nor ( n3470 , n2175 , n2182 , n2189 , n2195 );
and ( n3471 , n3469 , n3470 );
nor ( n3472 , n2176 , n2182 , n2189 , n2195 );
and ( n3473 , n2175 , n2183 , n2189 , n2195 );
and ( n3474 , n2176 , n2182 , n2189 , n2195 );
or ( n3475 , n3473 , n3474 );
and ( n3476 , n2175 , n2182 , n2189 , n2195 );
or ( n3477 , n3475 , n3476 );
or ( n3478 , n3472 , n3477 );
and ( n3479 , n627 , n3478 );
or ( n3480 , n2197 , n2999 , n3430 , n3436 , n3471 , n3479 );
and ( n3481 , n1078 , n3480 );
and ( n3482 , n627 , n1077 );
or ( n3483 , n3481 , n3482 );
and ( n3484 , n3483 , n721 );
not ( n3485 , n721 );
and ( n3486 , n627 , n3485 );
or ( n3487 , n3484 , n3486 );
buf ( n3488 , n3487 );
buf ( n3489 , n3488 );
not ( n3490 , n1077 );
xor ( n3491 , n1506 , n1120 );
xor ( n3492 , n1492 , n1120 );
xor ( n3493 , n1478 , n1120 );
xor ( n3494 , n1464 , n1120 );
xor ( n3495 , n1450 , n1120 );
xor ( n3496 , n1436 , n1120 );
xor ( n3497 , n1422 , n1120 );
xor ( n3498 , n1408 , n1120 );
xor ( n3499 , n1394 , n1120 );
xor ( n3500 , n1380 , n1120 );
xor ( n3501 , n1366 , n1120 );
xor ( n3502 , n1352 , n1120 );
xor ( n3503 , n1338 , n1120 );
xor ( n3504 , n1324 , n1120 );
and ( n3505 , n1511 , n1539 );
and ( n3506 , n3504 , n3505 );
and ( n3507 , n3503 , n3506 );
and ( n3508 , n3502 , n3507 );
and ( n3509 , n3501 , n3508 );
and ( n3510 , n3500 , n3509 );
and ( n3511 , n3499 , n3510 );
and ( n3512 , n3498 , n3511 );
and ( n3513 , n3497 , n3512 );
and ( n3514 , n3496 , n3513 );
and ( n3515 , n3495 , n3514 );
and ( n3516 , n3494 , n3515 );
and ( n3517 , n3493 , n3516 );
and ( n3518 , n3492 , n3517 );
and ( n3519 , n3491 , n3518 );
and ( n3520 , n3519 , n1508 );
and ( n3521 , n3520 , n1579 );
and ( n3522 , n3520 , n1582 );
not ( n3523 , n680 );
xor ( n3524 , n1640 , n1677 );
and ( n3525 , n3524 , n1120 );
and ( n3526 , n3523 , n3525 );
and ( n3527 , n3526 , n2024 );
and ( n3528 , n3525 , n2026 );
or ( n3529 , n3521 , n3522 , n3527 , n3528 );
and ( n3530 , n3529 , n2086 );
or ( n3531 , n2084 , n2088 );
or ( n3532 , n3531 , n2090 );
and ( n3533 , n683 , n3532 );
or ( n3534 , n3530 , n3533 );
and ( n3535 , n3534 , n2196 );
xor ( n3536 , n2950 , n2689 );
xor ( n3537 , n2941 , n2689 );
xor ( n3538 , n2932 , n2689 );
xor ( n3539 , n2923 , n2689 );
xor ( n3540 , n2914 , n2689 );
xor ( n3541 , n2905 , n2689 );
xor ( n3542 , n2896 , n2689 );
xor ( n3543 , n2887 , n2689 );
xor ( n3544 , n2878 , n2689 );
xor ( n3545 , n2869 , n2689 );
xor ( n3546 , n2860 , n2689 );
xor ( n3547 , n2851 , n2689 );
xor ( n3548 , n2842 , n2689 );
xor ( n3549 , n2833 , n2689 );
and ( n3550 , n2955 , n2985 );
and ( n3551 , n3549 , n3550 );
and ( n3552 , n3548 , n3551 );
and ( n3553 , n3547 , n3552 );
and ( n3554 , n3546 , n3553 );
and ( n3555 , n3545 , n3554 );
and ( n3556 , n3544 , n3555 );
and ( n3557 , n3543 , n3556 );
and ( n3558 , n3542 , n3557 );
and ( n3559 , n3541 , n3558 );
and ( n3560 , n3540 , n3559 );
and ( n3561 , n3539 , n3560 );
and ( n3562 , n3538 , n3561 );
and ( n3563 , n3537 , n3562 );
and ( n3564 , n3536 , n3563 );
and ( n3565 , n3564 , n2952 );
and ( n3566 , n3565 , n2086 );
or ( n3567 , n3566 , n3533 );
and ( n3568 , n3567 , n2998 );
xor ( n3569 , n3382 , n3122 );
xor ( n3570 , n3373 , n3122 );
xor ( n3571 , n3364 , n3122 );
xor ( n3572 , n3355 , n3122 );
xor ( n3573 , n3346 , n3122 );
xor ( n3574 , n3337 , n3122 );
xor ( n3575 , n3328 , n3122 );
xor ( n3576 , n3319 , n3122 );
xor ( n3577 , n3310 , n3122 );
xor ( n3578 , n3301 , n3122 );
xor ( n3579 , n3292 , n3122 );
xor ( n3580 , n3283 , n3122 );
xor ( n3581 , n3274 , n3122 );
xor ( n3582 , n3265 , n3122 );
and ( n3583 , n3387 , n3417 );
and ( n3584 , n3582 , n3583 );
and ( n3585 , n3581 , n3584 );
and ( n3586 , n3580 , n3585 );
and ( n3587 , n3579 , n3586 );
and ( n3588 , n3578 , n3587 );
and ( n3589 , n3577 , n3588 );
and ( n3590 , n3576 , n3589 );
and ( n3591 , n3575 , n3590 );
and ( n3592 , n3574 , n3591 );
and ( n3593 , n3573 , n3592 );
and ( n3594 , n3572 , n3593 );
and ( n3595 , n3571 , n3594 );
and ( n3596 , n3570 , n3595 );
and ( n3597 , n3569 , n3596 );
and ( n3598 , n3597 , n3384 );
and ( n3599 , n3598 , n2086 );
or ( n3600 , n3599 , n3533 );
and ( n3601 , n3600 , n3429 );
and ( n3602 , n2325 , n2086 );
or ( n3603 , n3602 , n3533 );
and ( n3604 , n3603 , n3435 );
not ( n3605 , n2325 );
not ( n3606 , n2329 );
not ( n3607 , n2333 );
not ( n3608 , n2337 );
not ( n3609 , n2341 );
not ( n3610 , n2345 );
not ( n3611 , n2349 );
not ( n3612 , n2353 );
not ( n3613 , n2357 );
not ( n3614 , n2361 );
not ( n3615 , n2365 );
not ( n3616 , n2413 );
not ( n3617 , n2423 );
not ( n3618 , n2433 );
not ( n3619 , n2443 );
and ( n3620 , n3437 , n3466 );
and ( n3621 , n3619 , n3620 );
and ( n3622 , n3618 , n3621 );
and ( n3623 , n3617 , n3622 );
and ( n3624 , n3616 , n3623 );
and ( n3625 , n3615 , n3624 );
and ( n3626 , n3614 , n3625 );
and ( n3627 , n3613 , n3626 );
and ( n3628 , n3612 , n3627 );
and ( n3629 , n3611 , n3628 );
and ( n3630 , n3610 , n3629 );
and ( n3631 , n3609 , n3630 );
and ( n3632 , n3608 , n3631 );
and ( n3633 , n3607 , n3632 );
and ( n3634 , n3606 , n3633 );
xor ( n3635 , n3605 , n3634 );
and ( n3636 , n3635 , n2086 );
or ( n3637 , n3636 , n3533 );
and ( n3638 , n3637 , n3470 );
and ( n3639 , n683 , n3478 );
or ( n3640 , n3535 , n3568 , n3601 , n3604 , n3638 , n3639 );
and ( n3641 , n3490 , n3640 );
and ( n3642 , n683 , n1077 );
or ( n3643 , n3641 , n3642 );
and ( n3644 , n3643 , n721 );
and ( n3645 , n683 , n3485 );
or ( n3646 , n3644 , n3645 );
buf ( n3647 , n3646 );
buf ( n3648 , n3647 );
not ( n3649 , n1077 );
not ( n3650 , n1508 );
and ( n3651 , n3650 , n1144 );
xor ( n3652 , n1523 , n1527 );
and ( n3653 , n3652 , n1508 );
or ( n3654 , n3651 , n3653 );
and ( n3655 , n3654 , n1579 );
and ( n3656 , n3654 , n1582 );
not ( n3657 , n680 );
and ( n3658 , n3657 , n1706 );
not ( n3659 , n1985 );
and ( n3660 , n3659 , n1712 );
xor ( n3661 , n2000 , n2006 );
and ( n3662 , n3661 , n1985 );
or ( n3663 , n3660 , n3662 );
and ( n3664 , n3663 , n680 );
or ( n3665 , n3658 , n3664 );
and ( n3666 , n3665 , n2024 );
and ( n3667 , n1706 , n2026 );
or ( n3668 , n3655 , n3656 , n3666 , n3667 );
and ( n3669 , n3668 , n2084 );
and ( n3670 , n579 , n2091 );
or ( n3671 , n3669 , n3670 );
and ( n3672 , n3671 , n2196 );
not ( n3673 , n2952 );
and ( n3674 , n3673 , n2716 );
xor ( n3675 , n2967 , n2973 );
and ( n3676 , n3675 , n2952 );
or ( n3677 , n3674 , n3676 );
and ( n3678 , n3677 , n2084 );
or ( n3679 , n3678 , n3670 );
and ( n3680 , n3679 , n2998 );
not ( n3681 , n3384 );
and ( n3682 , n3681 , n3148 );
xor ( n3683 , n3399 , n3405 );
and ( n3684 , n3683 , n3384 );
or ( n3685 , n3682 , n3684 );
and ( n3686 , n3685 , n2084 );
or ( n3687 , n3686 , n3670 );
and ( n3688 , n3687 , n3429 );
and ( n3689 , n2573 , n2084 );
or ( n3690 , n3689 , n3670 );
and ( n3691 , n3690 , n3435 );
xor ( n3692 , n3449 , n3454 );
and ( n3693 , n3692 , n2084 );
or ( n3694 , n3693 , n3670 );
and ( n3695 , n3694 , n3470 );
and ( n3696 , n579 , n3478 );
or ( n3697 , n3672 , n3680 , n3688 , n3691 , n3695 , n3696 );
and ( n3698 , n3649 , n3697 );
and ( n3699 , n579 , n1077 );
or ( n3700 , n3698 , n3699 );
and ( n3701 , n3700 , n721 );
and ( n3702 , n579 , n3485 );
or ( n3703 , n3701 , n3702 );
buf ( n3704 , n3703 );
buf ( n3705 , n3704 );
not ( n3706 , n1077 );
not ( n3707 , n1508 );
and ( n3708 , n3707 , n1132 );
xor ( n3709 , n1524 , n1526 );
and ( n3710 , n3709 , n1508 );
or ( n3711 , n3708 , n3710 );
and ( n3712 , n3711 , n1579 );
and ( n3713 , n3711 , n1582 );
not ( n3714 , n680 );
and ( n3715 , n3714 , n1695 );
not ( n3716 , n1985 );
and ( n3717 , n3716 , n1701 );
xor ( n3718 , n2001 , n2005 );
and ( n3719 , n3718 , n1985 );
or ( n3720 , n3717 , n3719 );
and ( n3721 , n3720 , n680 );
or ( n3722 , n3715 , n3721 );
and ( n3723 , n3722 , n2024 );
and ( n3724 , n1695 , n2026 );
or ( n3725 , n3712 , n3713 , n3723 , n3724 );
and ( n3726 , n3725 , n2086 );
and ( n3727 , n576 , n3532 );
or ( n3728 , n3726 , n3727 );
and ( n3729 , n3728 , n2196 );
not ( n3730 , n2952 );
and ( n3731 , n3730 , n2707 );
xor ( n3732 , n2968 , n2972 );
and ( n3733 , n3732 , n2952 );
or ( n3734 , n3731 , n3733 );
and ( n3735 , n3734 , n2086 );
or ( n3736 , n3735 , n3727 );
and ( n3737 , n3736 , n2998 );
not ( n3738 , n3384 );
and ( n3739 , n3738 , n3139 );
xor ( n3740 , n3400 , n3404 );
and ( n3741 , n3740 , n3384 );
or ( n3742 , n3739 , n3741 );
and ( n3743 , n3742 , n2086 );
or ( n3744 , n3743 , n3727 );
and ( n3745 , n3744 , n3429 );
and ( n3746 , n2583 , n2086 );
or ( n3747 , n3746 , n3727 );
and ( n3748 , n3747 , n3435 );
xor ( n3749 , n3450 , n3453 );
and ( n3750 , n3749 , n2086 );
or ( n3751 , n3750 , n3727 );
and ( n3752 , n3751 , n3470 );
and ( n3753 , n576 , n3478 );
or ( n3754 , n3729 , n3737 , n3745 , n3748 , n3752 , n3753 );
and ( n3755 , n3706 , n3754 );
and ( n3756 , n576 , n1077 );
or ( n3757 , n3755 , n3756 );
and ( n3758 , n3757 , n721 );
and ( n3759 , n576 , n3485 );
or ( n3760 , n3758 , n3759 );
buf ( n3761 , n3760 );
buf ( n3762 , n3761 );
not ( n3763 , n1077 );
and ( n3764 , n1411 , n3477 );
not ( n3765 , n1508 );
and ( n3766 , n3765 , n1408 );
xor ( n3767 , n3498 , n3511 );
and ( n3768 , n3767 , n1508 );
or ( n3769 , n3766 , n3768 );
and ( n3770 , n3769 , n1579 );
and ( n3771 , n3769 , n1582 );
not ( n3772 , n680 );
and ( n3773 , n3772 , n1911 );
not ( n3774 , n1985 );
and ( n3775 , n3774 , n1917 );
xor ( n3776 , n1917 , n1680 );
xor ( n3777 , n1906 , n1680 );
xor ( n3778 , n1895 , n1680 );
xor ( n3779 , n1884 , n1680 );
xor ( n3780 , n1873 , n1680 );
xor ( n3781 , n1862 , n1680 );
xor ( n3782 , n1851 , n1680 );
and ( n3783 , n1988 , n2018 );
and ( n3784 , n3782 , n3783 );
and ( n3785 , n3781 , n3784 );
and ( n3786 , n3780 , n3785 );
and ( n3787 , n3779 , n3786 );
and ( n3788 , n3778 , n3787 );
and ( n3789 , n3777 , n3788 );
xor ( n3790 , n3776 , n3789 );
and ( n3791 , n3790 , n1985 );
or ( n3792 , n3775 , n3791 );
and ( n3793 , n3792 , n680 );
or ( n3794 , n3773 , n3793 );
and ( n3795 , n3794 , n2024 );
and ( n3796 , n1911 , n2026 );
or ( n3797 , n3770 , n3771 , n3795 , n3796 );
and ( n3798 , n3797 , n2090 );
or ( n3799 , n2084 , n2086 );
or ( n3800 , n3799 , n2088 );
and ( n3801 , n1411 , n3800 );
or ( n3802 , n3798 , n3801 );
and ( n3803 , n3802 , n2196 );
not ( n3804 , n2952 );
and ( n3805 , n3804 , n2887 );
xor ( n3806 , n3543 , n3556 );
and ( n3807 , n3806 , n2952 );
or ( n3808 , n3805 , n3807 );
and ( n3809 , n3808 , n2090 );
or ( n3810 , n3809 , n3801 );
and ( n3811 , n3810 , n2998 );
not ( n3812 , n3384 );
and ( n3813 , n3812 , n3319 );
xor ( n3814 , n3576 , n3589 );
and ( n3815 , n3814 , n3384 );
or ( n3816 , n3813 , n3815 );
and ( n3817 , n3816 , n2090 );
or ( n3818 , n3817 , n3801 );
and ( n3819 , n3818 , n3429 );
and ( n3820 , n2357 , n2090 );
or ( n3821 , n3820 , n3801 );
and ( n3822 , n3821 , n3435 );
and ( n3823 , n2357 , n3472 );
xor ( n3824 , n3613 , n3626 );
and ( n3825 , n3824 , n2090 );
or ( n3826 , n3825 , n3801 );
and ( n3827 , n3826 , n3470 );
or ( n3828 , n3764 , n3803 , n3811 , n3819 , n3822 , n3823 , n3827 );
and ( n3829 , n3763 , n3828 );
and ( n3830 , n1411 , n1077 );
or ( n3831 , n3829 , n3830 );
and ( n3832 , n3831 , n721 );
and ( n3833 , n652 , n3485 );
or ( n3834 , n3832 , n3833 );
buf ( n3835 , n3834 );
buf ( n3836 , n3835 );
not ( n3837 , n1077 );
not ( n3838 , n1508 );
and ( n3839 , n3838 , n1436 );
xor ( n3840 , n3496 , n3513 );
and ( n3841 , n3840 , n1508 );
or ( n3842 , n3839 , n3841 );
and ( n3843 , n3842 , n1579 );
and ( n3844 , n3842 , n1582 );
not ( n3845 , n680 );
and ( n3846 , n3845 , n1933 );
not ( n3847 , n1985 );
and ( n3848 , n3847 , n1939 );
xor ( n3849 , n1939 , n1680 );
xor ( n3850 , n1928 , n1680 );
and ( n3851 , n3776 , n3789 );
and ( n3852 , n3850 , n3851 );
xor ( n3853 , n3849 , n3852 );
and ( n3854 , n3853 , n1985 );
or ( n3855 , n3848 , n3854 );
and ( n3856 , n3855 , n680 );
or ( n3857 , n3846 , n3856 );
and ( n3858 , n3857 , n2024 );
and ( n3859 , n1933 , n2026 );
or ( n3860 , n3843 , n3844 , n3858 , n3859 );
and ( n3861 , n3860 , n2086 );
and ( n3862 , n663 , n3532 );
or ( n3863 , n3861 , n3862 );
and ( n3864 , n3863 , n2196 );
not ( n3865 , n2952 );
and ( n3866 , n3865 , n2905 );
xor ( n3867 , n3541 , n3558 );
and ( n3868 , n3867 , n2952 );
or ( n3869 , n3866 , n3868 );
and ( n3870 , n3869 , n2086 );
or ( n3871 , n3870 , n3862 );
and ( n3872 , n3871 , n2998 );
not ( n3873 , n3384 );
and ( n3874 , n3873 , n3337 );
xor ( n3875 , n3574 , n3591 );
and ( n3876 , n3875 , n3384 );
or ( n3877 , n3874 , n3876 );
and ( n3878 , n3877 , n2086 );
or ( n3879 , n3878 , n3862 );
and ( n3880 , n3879 , n3429 );
and ( n3881 , n2349 , n2086 );
or ( n3882 , n3881 , n3862 );
and ( n3883 , n3882 , n3435 );
xor ( n3884 , n3611 , n3628 );
and ( n3885 , n3884 , n2086 );
or ( n3886 , n3885 , n3862 );
and ( n3887 , n3886 , n3470 );
and ( n3888 , n663 , n3478 );
or ( n3889 , n3864 , n3872 , n3880 , n3883 , n3887 , n3888 );
and ( n3890 , n3837 , n3889 );
and ( n3891 , n663 , n1077 );
or ( n3892 , n3890 , n3891 );
and ( n3893 , n3892 , n721 );
and ( n3894 , n663 , n3485 );
or ( n3895 , n3893 , n3894 );
buf ( n3896 , n3895 );
buf ( n3897 , n3896 );
not ( n3898 , n1077 );
and ( n3899 , n633 , n3477 );
not ( n3900 , n1508 );
and ( n3901 , n3900 , n1338 );
xor ( n3902 , n3503 , n3506 );
and ( n3903 , n3902 , n1508 );
or ( n3904 , n3901 , n3903 );
and ( n3905 , n3904 , n1579 );
and ( n3906 , n3904 , n1582 );
not ( n3907 , n680 );
and ( n3908 , n3907 , n1856 );
not ( n3909 , n1985 );
and ( n3910 , n3909 , n1862 );
xor ( n3911 , n3781 , n3784 );
and ( n3912 , n3911 , n1985 );
or ( n3913 , n3910 , n3912 );
and ( n3914 , n3913 , n680 );
or ( n3915 , n3908 , n3914 );
and ( n3916 , n3915 , n2024 );
and ( n3917 , n1856 , n2026 );
or ( n3918 , n3905 , n3906 , n3916 , n3917 );
and ( n3919 , n3918 , n2088 );
or ( n3920 , n3799 , n2090 );
and ( n3921 , n633 , n3920 );
or ( n3922 , n3919 , n3921 );
and ( n3923 , n3922 , n2196 );
not ( n3924 , n2952 );
and ( n3925 , n3924 , n2842 );
xor ( n3926 , n3548 , n3551 );
and ( n3927 , n3926 , n2952 );
or ( n3928 , n3925 , n3927 );
and ( n3929 , n3928 , n2088 );
or ( n3930 , n3929 , n3921 );
and ( n3931 , n3930 , n2998 );
not ( n3932 , n3384 );
and ( n3933 , n3932 , n3274 );
xor ( n3934 , n3581 , n3584 );
and ( n3935 , n3934 , n3384 );
or ( n3936 , n3933 , n3935 );
and ( n3937 , n3936 , n2088 );
or ( n3938 , n3937 , n3921 );
and ( n3939 , n3938 , n3429 );
and ( n3940 , n2433 , n2088 );
or ( n3941 , n3940 , n3921 );
and ( n3942 , n3941 , n3435 );
and ( n3943 , n1341 , n3472 );
xor ( n3944 , n3618 , n3621 );
and ( n3945 , n3944 , n2088 );
or ( n3946 , n3945 , n3921 );
and ( n3947 , n3946 , n3470 );
or ( n3948 , n3899 , n3923 , n3931 , n3939 , n3942 , n3943 , n3947 );
and ( n3949 , n3898 , n3948 );
and ( n3950 , n633 , n1077 );
or ( n3951 , n3949 , n3950 );
and ( n3952 , n3951 , n721 );
and ( n3953 , n633 , n3485 );
or ( n3954 , n3952 , n3953 );
buf ( n3955 , n3954 );
buf ( n3956 , n3955 );
not ( n3957 , n1077 );
and ( n3958 , n637 , n3477 );
not ( n3959 , n1508 );
and ( n3960 , n3959 , n1352 );
xor ( n3961 , n3502 , n3507 );
and ( n3962 , n3961 , n1508 );
or ( n3963 , n3960 , n3962 );
and ( n3964 , n3963 , n1579 );
and ( n3965 , n3963 , n1582 );
not ( n3966 , n680 );
and ( n3967 , n3966 , n1867 );
not ( n3968 , n1985 );
and ( n3969 , n3968 , n1873 );
xor ( n3970 , n3780 , n3785 );
and ( n3971 , n3970 , n1985 );
or ( n3972 , n3969 , n3971 );
and ( n3973 , n3972 , n680 );
or ( n3974 , n3967 , n3973 );
and ( n3975 , n3974 , n2024 );
and ( n3976 , n1867 , n2026 );
or ( n3977 , n3964 , n3965 , n3975 , n3976 );
and ( n3978 , n3977 , n2088 );
and ( n3979 , n637 , n3920 );
or ( n3980 , n3978 , n3979 );
and ( n3981 , n3980 , n2196 );
not ( n3982 , n2952 );
and ( n3983 , n3982 , n2851 );
xor ( n3984 , n3547 , n3552 );
and ( n3985 , n3984 , n2952 );
or ( n3986 , n3983 , n3985 );
and ( n3987 , n3986 , n2088 );
or ( n3988 , n3987 , n3979 );
and ( n3989 , n3988 , n2998 );
not ( n3990 , n3384 );
and ( n3991 , n3990 , n3283 );
xor ( n3992 , n3580 , n3585 );
and ( n3993 , n3992 , n3384 );
or ( n3994 , n3991 , n3993 );
and ( n3995 , n3994 , n2088 );
or ( n3996 , n3995 , n3979 );
and ( n3997 , n3996 , n3429 );
and ( n3998 , n2423 , n2088 );
or ( n3999 , n3998 , n3979 );
and ( n4000 , n3999 , n3435 );
and ( n4001 , n1355 , n3472 );
xor ( n4002 , n3617 , n3622 );
and ( n4003 , n4002 , n2088 );
or ( n4004 , n4003 , n3979 );
and ( n4005 , n4004 , n3470 );
or ( n4006 , n3958 , n3981 , n3989 , n3997 , n4000 , n4001 , n4005 );
and ( n4007 , n3957 , n4006 );
and ( n4008 , n637 , n1077 );
or ( n4009 , n4007 , n4008 );
and ( n4010 , n4009 , n721 );
and ( n4011 , n637 , n3485 );
or ( n4012 , n4010 , n4011 );
buf ( n4013 , n4012 );
buf ( n4014 , n4013 );
not ( n4015 , n1077 );
and ( n4016 , n1173 , n3477 );
not ( n4017 , n1508 );
and ( n4018 , n4017 , n1170 );
xor ( n4019 , n1521 , n1529 );
and ( n4020 , n4019 , n1508 );
or ( n4021 , n4018 , n4020 );
and ( n4022 , n4021 , n1579 );
and ( n4023 , n4021 , n1582 );
not ( n4024 , n680 );
and ( n4025 , n4024 , n1728 );
not ( n4026 , n1985 );
and ( n4027 , n4026 , n1734 );
xor ( n4028 , n1998 , n2008 );
and ( n4029 , n4028 , n1985 );
or ( n4030 , n4027 , n4029 );
and ( n4031 , n4030 , n680 );
or ( n4032 , n4025 , n4031 );
and ( n4033 , n4032 , n2024 );
and ( n4034 , n1728 , n2026 );
or ( n4035 , n4022 , n4023 , n4033 , n4034 );
and ( n4036 , n4035 , n2090 );
and ( n4037 , n1173 , n3800 );
or ( n4038 , n4036 , n4037 );
and ( n4039 , n4038 , n2196 );
not ( n4040 , n2952 );
and ( n4041 , n4040 , n2734 );
xor ( n4042 , n2965 , n2975 );
and ( n4043 , n4042 , n2952 );
or ( n4044 , n4041 , n4043 );
and ( n4045 , n4044 , n2090 );
or ( n4046 , n4045 , n4037 );
and ( n4047 , n4046 , n2998 );
not ( n4048 , n3384 );
and ( n4049 , n4048 , n3166 );
xor ( n4050 , n3397 , n3407 );
and ( n4051 , n4050 , n3384 );
or ( n4052 , n4049 , n4051 );
and ( n4053 , n4052 , n2090 );
or ( n4054 , n4053 , n4037 );
and ( n4055 , n4054 , n3429 );
and ( n4056 , n2553 , n2090 );
or ( n4057 , n4056 , n4037 );
and ( n4058 , n4057 , n3435 );
and ( n4059 , n2553 , n3472 );
xor ( n4060 , n3447 , n3456 );
and ( n4061 , n4060 , n2090 );
or ( n4062 , n4061 , n4037 );
and ( n4063 , n4062 , n3470 );
or ( n4064 , n4016 , n4039 , n4047 , n4055 , n4058 , n4059 , n4063 );
and ( n4065 , n4015 , n4064 );
and ( n4066 , n1173 , n1077 );
or ( n4067 , n4065 , n4066 );
and ( n4068 , n4067 , n721 );
and ( n4069 , n585 , n3485 );
or ( n4070 , n4068 , n4069 );
buf ( n4071 , n4070 );
buf ( n4072 , n4071 );
not ( n4073 , n1077 );
not ( n4074 , n1508 );
and ( n4075 , n4074 , n1464 );
xor ( n4076 , n3494 , n3515 );
and ( n4077 , n4076 , n1508 );
or ( n4078 , n4075 , n4077 );
and ( n4079 , n4078 , n1579 );
and ( n4080 , n4078 , n1582 );
not ( n4081 , n680 );
and ( n4082 , n4081 , n1955 );
not ( n4083 , n1985 );
and ( n4084 , n4083 , n1961 );
xor ( n4085 , n1961 , n1680 );
xor ( n4086 , n1950 , n1680 );
and ( n4087 , n3849 , n3852 );
and ( n4088 , n4086 , n4087 );
xor ( n4089 , n4085 , n4088 );
and ( n4090 , n4089 , n1985 );
or ( n4091 , n4084 , n4090 );
and ( n4092 , n4091 , n680 );
or ( n4093 , n4082 , n4092 );
and ( n4094 , n4093 , n2024 );
and ( n4095 , n1955 , n2026 );
or ( n4096 , n4079 , n4080 , n4094 , n4095 );
and ( n4097 , n4096 , n2084 );
and ( n4098 , n670 , n2091 );
or ( n4099 , n4097 , n4098 );
and ( n4100 , n4099 , n2196 );
not ( n4101 , n2952 );
and ( n4102 , n4101 , n2923 );
xor ( n4103 , n3539 , n3560 );
and ( n4104 , n4103 , n2952 );
or ( n4105 , n4102 , n4104 );
and ( n4106 , n4105 , n2084 );
or ( n4107 , n4106 , n4098 );
and ( n4108 , n4107 , n2998 );
not ( n4109 , n3384 );
and ( n4110 , n4109 , n3355 );
xor ( n4111 , n3572 , n3593 );
and ( n4112 , n4111 , n3384 );
or ( n4113 , n4110 , n4112 );
and ( n4114 , n4113 , n2084 );
or ( n4115 , n4114 , n4098 );
and ( n4116 , n4115 , n3429 );
and ( n4117 , n2341 , n2084 );
or ( n4118 , n4117 , n4098 );
and ( n4119 , n4118 , n3435 );
xor ( n4120 , n3609 , n3630 );
and ( n4121 , n4120 , n2084 );
or ( n4122 , n4121 , n4098 );
and ( n4123 , n4122 , n3470 );
and ( n4124 , n670 , n3478 );
or ( n4125 , n4100 , n4108 , n4116 , n4119 , n4123 , n4124 );
and ( n4126 , n4073 , n4125 );
and ( n4127 , n670 , n1077 );
or ( n4128 , n4126 , n4127 );
and ( n4129 , n4128 , n721 );
and ( n4130 , n670 , n3485 );
or ( n4131 , n4129 , n4130 );
buf ( n4132 , n4131 );
buf ( n4133 , n4132 );
endmodule

