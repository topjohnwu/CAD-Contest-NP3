//
// Conformal-LEC Version 15.20-d227 ( 10-Mar-2016) ( 64 bit executable)
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n8 , n9 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 );
input n0 , n1 , n2 , n3 , n4 , n5 , n8 , n9 , n11 , n12 , n13 , n14 , n15 ;
output n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;

wire n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , 
     n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , 
     n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , 
     n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , 
     n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , 
     n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , 
     n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , 
     n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , 
     n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , 
     n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , 
     n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , 
     n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , 
     n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , 
     n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , 
     n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , 
     n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , 
     n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , 
     n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , 
     n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , 
     n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , 
     n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , 
     n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , 
     n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , 
     n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , 
     n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , 
     n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , 
     n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , 
     n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , 
     n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , 
     n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , 
     n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , 
     n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , 
     n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , 
     n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , 
     n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , 
     n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , 
     n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , 
     n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , 
     n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , 
     n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , 
     n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , 
     n473 , n474 , n475 ;
buf ( n23 , n432 );
buf ( n26 , n435 );
buf ( n31 , n438 );
buf ( n28 , n441 );
buf ( n29 , n444 );
buf ( n21 , n447 );
buf ( n27 , n450 );
buf ( n30 , n453 );
buf ( n19 , n456 );
buf ( n18 , n459 );
buf ( n16 , n462 );
buf ( n22 , n466 );
buf ( n20 , n470 );
buf ( n24 , n474 );
buf ( n25 , n475 );
buf ( n17 , 1'b0 );
buf ( n70 , n15 );
buf ( n71 , n4 );
buf ( n72 , n1 );
buf ( n73 , n2 );
buf ( n74 , n9 );
buf ( n75 , n5 );
buf ( n76 , n12 );
buf ( n77 , n0 );
buf ( n78 , n14 );
buf ( n79 , n13 );
buf ( n80 , n11 );
buf ( n81 , n8 );
buf ( n82 , n3 );
buf ( n83 , n70 );
buf ( n84 , n75 );
and ( n85 , n83 , n84 );
buf ( n86 , n73 );
not ( n87 , n86 );
not ( n88 , n84 );
and ( n89 , n88 , n86 );
nor ( n90 , n87 , n89 );
buf ( n91 , n72 );
buf ( n92 , n76 );
and ( n93 , n91 , n92 );
and ( n94 , n90 , n93 );
buf ( n95 , n71 );
buf ( n96 , n77 );
and ( n97 , n95 , n96 );
and ( n98 , n93 , n97 );
and ( n99 , n90 , n97 );
or ( n100 , n94 , n98 , n99 );
not ( n101 , n91 );
and ( n102 , n88 , n91 );
nor ( n103 , n101 , n102 );
and ( n104 , n100 , n103 );
and ( n105 , n95 , n92 );
and ( n106 , n103 , n105 );
and ( n107 , n100 , n105 );
or ( n108 , n104 , n106 , n107 );
not ( n109 , n95 );
and ( n110 , n88 , n95 );
nor ( n111 , n109 , n110 );
and ( n112 , n108 , n111 );
not ( n113 , n83 );
and ( n114 , n113 , n92 );
not ( n115 , n92 );
nor ( n116 , n114 , n115 );
and ( n117 , n111 , n116 );
and ( n118 , n108 , n116 );
or ( n119 , n112 , n117 , n118 );
and ( n120 , n85 , n119 );
xor ( n121 , n85 , n119 );
xor ( n122 , n108 , n111 );
xor ( n123 , n122 , n116 );
buf ( n124 , n74 );
not ( n125 , n124 );
and ( n126 , n88 , n124 );
nor ( n127 , n125 , n126 );
and ( n128 , n86 , n92 );
and ( n129 , n127 , n128 );
buf ( n130 , n79 );
and ( n131 , n113 , n130 );
not ( n132 , n130 );
nor ( n133 , n131 , n132 );
and ( n134 , n128 , n133 );
and ( n135 , n127 , n133 );
or ( n136 , n129 , n134 , n135 );
and ( n137 , n86 , n96 );
buf ( n138 , n78 );
and ( n139 , n91 , n138 );
and ( n140 , n137 , n139 );
and ( n141 , n95 , n130 );
and ( n142 , n139 , n141 );
and ( n143 , n137 , n141 );
or ( n144 , n140 , n142 , n143 );
and ( n145 , n91 , n96 );
and ( n146 , n144 , n145 );
and ( n147 , n95 , n138 );
and ( n148 , n145 , n147 );
and ( n149 , n144 , n147 );
or ( n150 , n146 , n148 , n149 );
and ( n151 , n136 , n150 );
xor ( n152 , n90 , n93 );
xor ( n153 , n152 , n97 );
and ( n154 , n150 , n153 );
and ( n155 , n136 , n153 );
or ( n156 , n151 , n154 , n155 );
and ( n157 , n113 , n96 );
not ( n158 , n96 );
nor ( n159 , n157 , n158 );
and ( n160 , n156 , n159 );
xor ( n161 , n100 , n103 );
xor ( n162 , n161 , n105 );
and ( n163 , n159 , n162 );
and ( n164 , n156 , n162 );
or ( n165 , n160 , n163 , n164 );
and ( n166 , n123 , n165 );
xor ( n167 , n123 , n165 );
xor ( n168 , n156 , n159 );
xor ( n169 , n168 , n162 );
and ( n170 , n86 , n138 );
and ( n171 , n91 , n130 );
and ( n172 , n170 , n171 );
buf ( n173 , n80 );
and ( n174 , n95 , n173 );
and ( n175 , n171 , n174 );
and ( n176 , n170 , n174 );
or ( n177 , n172 , n175 , n176 );
buf ( n178 , n92 );
and ( n179 , n124 , n96 );
and ( n180 , n178 , n179 );
and ( n181 , n177 , n180 );
xor ( n182 , n137 , n139 );
xor ( n183 , n182 , n141 );
and ( n184 , n180 , n183 );
and ( n185 , n177 , n183 );
or ( n186 , n181 , n184 , n185 );
xor ( n187 , n127 , n128 );
xor ( n188 , n187 , n133 );
and ( n189 , n186 , n188 );
xor ( n190 , n144 , n145 );
xor ( n191 , n190 , n147 );
and ( n192 , n188 , n191 );
and ( n193 , n186 , n191 );
or ( n194 , n189 , n192 , n193 );
and ( n195 , n113 , n138 );
not ( n196 , n138 );
nor ( n197 , n195 , n196 );
and ( n198 , n194 , n197 );
xor ( n199 , n136 , n150 );
xor ( n200 , n199 , n153 );
and ( n201 , n197 , n200 );
and ( n202 , n194 , n200 );
or ( n203 , n198 , n201 , n202 );
and ( n204 , n169 , n203 );
xor ( n205 , n169 , n203 );
xor ( n206 , n194 , n197 );
xor ( n207 , n206 , n200 );
buf ( n208 , n88 );
not ( n209 , n208 );
and ( n210 , n124 , n92 );
and ( n211 , n209 , n210 );
and ( n212 , n113 , n173 );
not ( n213 , n173 );
nor ( n214 , n212 , n213 );
and ( n215 , n210 , n214 );
and ( n216 , n209 , n214 );
or ( n217 , n211 , n215 , n216 );
and ( n218 , n86 , n130 );
and ( n219 , n91 , n173 );
and ( n220 , n218 , n219 );
buf ( n221 , n81 );
and ( n222 , n95 , n221 );
and ( n223 , n219 , n222 );
and ( n224 , n218 , n222 );
or ( n225 , n220 , n223 , n224 );
xor ( n226 , n170 , n171 );
xor ( n227 , n226 , n174 );
and ( n228 , n225 , n227 );
xor ( n229 , n178 , n179 );
and ( n230 , n227 , n229 );
and ( n231 , n225 , n229 );
or ( n232 , n228 , n230 , n231 );
xor ( n233 , n209 , n210 );
xor ( n234 , n233 , n214 );
and ( n235 , n232 , n234 );
xor ( n236 , n177 , n180 );
xor ( n237 , n236 , n183 );
and ( n238 , n234 , n237 );
and ( n239 , n232 , n237 );
or ( n240 , n235 , n238 , n239 );
and ( n241 , n217 , n240 );
xor ( n242 , n186 , n188 );
xor ( n243 , n242 , n191 );
and ( n244 , n240 , n243 );
and ( n245 , n217 , n243 );
or ( n246 , n241 , n244 , n245 );
and ( n247 , n207 , n246 );
xor ( n248 , n207 , n246 );
xor ( n249 , n217 , n240 );
xor ( n250 , n249 , n243 );
buf ( n251 , n92 );
buf ( n252 , n96 );
and ( n253 , n251 , n252 );
and ( n254 , n124 , n138 );
and ( n255 , n252 , n254 );
and ( n256 , n251 , n254 );
or ( n257 , n253 , n255 , n256 );
buf ( n258 , n88 );
not ( n259 , n258 );
and ( n260 , n257 , n259 );
and ( n261 , n113 , n221 );
not ( n262 , n221 );
nor ( n263 , n261 , n262 );
and ( n264 , n259 , n263 );
and ( n265 , n257 , n263 );
or ( n266 , n260 , n264 , n265 );
and ( n267 , n86 , n173 );
and ( n268 , n91 , n221 );
and ( n269 , n267 , n268 );
buf ( n270 , n82 );
and ( n271 , n95 , n270 );
and ( n272 , n268 , n271 );
and ( n273 , n267 , n271 );
or ( n274 , n269 , n272 , n273 );
xor ( n275 , n251 , n252 );
xor ( n276 , n275 , n254 );
and ( n277 , n274 , n276 );
xor ( n278 , n218 , n219 );
xor ( n279 , n278 , n222 );
and ( n280 , n276 , n279 );
and ( n281 , n274 , n279 );
or ( n282 , n277 , n280 , n281 );
xor ( n283 , n257 , n259 );
xor ( n284 , n283 , n263 );
and ( n285 , n282 , n284 );
xor ( n286 , n225 , n227 );
xor ( n287 , n286 , n229 );
and ( n288 , n284 , n287 );
and ( n289 , n282 , n287 );
or ( n290 , n285 , n288 , n289 );
and ( n291 , n266 , n290 );
xor ( n292 , n232 , n234 );
xor ( n293 , n292 , n237 );
and ( n294 , n290 , n293 );
and ( n295 , n266 , n293 );
or ( n296 , n291 , n294 , n295 );
and ( n297 , n250 , n296 );
xor ( n298 , n250 , n296 );
xor ( n299 , n266 , n290 );
xor ( n300 , n299 , n293 );
and ( n301 , n86 , n221 );
and ( n302 , n91 , n270 );
and ( n303 , n301 , n302 );
and ( n304 , n124 , n130 );
and ( n305 , n303 , n304 );
xor ( n306 , n267 , n268 );
xor ( n307 , n306 , n271 );
and ( n308 , n304 , n307 );
and ( n309 , n303 , n307 );
or ( n310 , n305 , n308 , n309 );
xor ( n311 , n274 , n276 );
xor ( n312 , n311 , n279 );
and ( n313 , n310 , n312 );
and ( n314 , n113 , n270 );
not ( n315 , n270 );
nor ( n316 , n314 , n315 );
buf ( n317 , n316 );
and ( n318 , n312 , n317 );
and ( n319 , n310 , n317 );
or ( n320 , n313 , n318 , n319 );
xor ( n321 , n282 , n284 );
xor ( n322 , n321 , n287 );
and ( n323 , n320 , n322 );
buf ( n324 , n323 );
and ( n325 , n300 , n324 );
xor ( n326 , n300 , n324 );
buf ( n327 , n320 );
xor ( n328 , n327 , n322 );
buf ( n329 , n96 );
buf ( n330 , n138 );
and ( n331 , n329 , n330 );
buf ( n332 , n331 );
buf ( n333 , n173 );
and ( n334 , n124 , n221 );
and ( n335 , n333 , n334 );
and ( n336 , n86 , n270 );
and ( n337 , n334 , n336 );
and ( n338 , n333 , n336 );
or ( n339 , n335 , n337 , n338 );
and ( n340 , n124 , n173 );
and ( n341 , n339 , n340 );
xor ( n342 , n301 , n302 );
and ( n343 , n340 , n342 );
and ( n344 , n339 , n342 );
or ( n345 , n341 , n343 , n344 );
buf ( n346 , n329 );
xor ( n347 , n346 , n330 );
and ( n348 , n345 , n347 );
xor ( n349 , n303 , n304 );
xor ( n350 , n349 , n307 );
and ( n351 , n347 , n350 );
and ( n352 , n345 , n350 );
or ( n353 , n348 , n351 , n352 );
and ( n354 , n332 , n353 );
xor ( n355 , n310 , n312 );
xor ( n356 , n355 , n317 );
and ( n357 , n353 , n356 );
and ( n358 , n332 , n356 );
or ( n359 , n354 , n357 , n358 );
and ( n360 , n328 , n359 );
xor ( n361 , n328 , n359 );
xor ( n362 , n332 , n353 );
xor ( n363 , n362 , n356 );
buf ( n364 , n138 );
buf ( n365 , n130 );
and ( n366 , n364 , n365 );
buf ( n367 , n173 );
buf ( n368 , n221 );
and ( n369 , n367 , n368 );
and ( n370 , n124 , n270 );
and ( n371 , n368 , n370 );
and ( n372 , n367 , n370 );
or ( n373 , n369 , n371 , n372 );
buf ( n374 , n130 );
and ( n375 , n373 , n374 );
xor ( n376 , n333 , n334 );
xor ( n377 , n376 , n336 );
and ( n378 , n374 , n377 );
and ( n379 , n373 , n377 );
or ( n380 , n375 , n378 , n379 );
xor ( n381 , n364 , n365 );
and ( n382 , n380 , n381 );
xor ( n383 , n339 , n340 );
xor ( n384 , n383 , n342 );
and ( n385 , n381 , n384 );
and ( n386 , n380 , n384 );
or ( n387 , n382 , n385 , n386 );
and ( n388 , n366 , n387 );
xor ( n389 , n345 , n347 );
xor ( n390 , n389 , n350 );
and ( n391 , n387 , n390 );
and ( n392 , n366 , n390 );
or ( n393 , n388 , n391 , n392 );
and ( n394 , n363 , n393 );
xor ( n395 , n363 , n393 );
xor ( n396 , n366 , n387 );
xor ( n397 , n396 , n390 );
buf ( n398 , n221 );
buf ( n399 , n270 );
and ( n400 , n398 , n399 );
buf ( n401 , n400 );
xor ( n402 , n367 , n368 );
xor ( n403 , n402 , n370 );
and ( n404 , n401 , n403 );
buf ( n405 , n404 );
xor ( n406 , n373 , n374 );
xor ( n407 , n406 , n377 );
and ( n408 , n405 , n407 );
buf ( n409 , n408 );
xor ( n410 , n380 , n381 );
xor ( n411 , n410 , n384 );
and ( n412 , n409 , n411 );
and ( n413 , n397 , n412 );
buf ( n414 , n413 );
and ( n415 , n395 , n414 );
or ( n416 , n394 , n415 );
and ( n417 , n361 , n416 );
or ( n418 , n360 , n417 );
and ( n419 , n326 , n418 );
or ( n420 , n325 , n419 );
and ( n421 , n298 , n420 );
or ( n422 , n297 , n421 );
and ( n423 , n248 , n422 );
or ( n424 , n247 , n423 );
and ( n425 , n205 , n424 );
or ( n426 , n204 , n425 );
and ( n427 , n167 , n426 );
or ( n428 , n166 , n427 );
and ( n429 , n121 , n428 );
or ( n430 , n120 , n429 );
buf ( n431 , n430 );
buf ( n432 , n431 );
xor ( n433 , n121 , n428 );
buf ( n434 , n433 );
buf ( n435 , n434 );
xor ( n436 , n167 , n426 );
buf ( n437 , n436 );
buf ( n438 , n437 );
xor ( n439 , n205 , n424 );
buf ( n440 , n439 );
buf ( n441 , n440 );
xor ( n442 , n248 , n422 );
buf ( n443 , n442 );
buf ( n444 , n443 );
xor ( n445 , n298 , n420 );
buf ( n446 , n445 );
buf ( n447 , n446 );
xor ( n448 , n326 , n418 );
buf ( n449 , n448 );
buf ( n450 , n449 );
xor ( n451 , n361 , n416 );
buf ( n452 , n451 );
buf ( n453 , n452 );
xor ( n454 , n395 , n414 );
buf ( n455 , n454 );
buf ( n456 , n455 );
xor ( n457 , n397 , n412 );
buf ( n458 , n457 );
buf ( n459 , n458 );
xor ( n460 , n409 , n411 );
buf ( n461 , n460 );
buf ( n462 , n461 );
buf ( n463 , n405 );
xor ( n464 , n463 , n407 );
buf ( n465 , n464 );
buf ( n466 , n465 );
buf ( n467 , n401 );
xor ( n468 , n467 , n403 );
buf ( n469 , n468 );
buf ( n470 , n469 );
buf ( n471 , n398 );
xor ( n472 , n471 , n399 );
buf ( n473 , n472 );
buf ( n474 , n473 );
buf ( n475 , n270 );
endmodule

