//
// Conformal-LEC Version 16.10-d005 ( 21-Apr-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 ;
output n512 , n513 , n514 , n515 , n516 ;

wire n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , 
     n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , 
     n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , 
     n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , 
     n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , 
     n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , 
     n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , 
     n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , 
     n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , 
     n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , 
     n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , 
     n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , 
     n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , 
     n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , 
     n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , 
     n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , 
     n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , 
     n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , 
     n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , 
     n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , 
     n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , 
     n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , 
     n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , 
     n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , 
     n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , 
     n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , 
     n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , 
     n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , 
     n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , 
     n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , 
     n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , 
     n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , 
     n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , 
     n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , 
     n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , 
     n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , 
     n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , 
     n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , 
     n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , 
     n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , 
     n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , 
     n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , 
     n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , 
     n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , 
     n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , 
     n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , 
     n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , 
     n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , 
     n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , 
     n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , 
     n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , 
     n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , 
     n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , 
     n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , 
     n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , 
     n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , 
     n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , 
     n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , 
     n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , 
     n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , 
     n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , 
     n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , 
     n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , 
     n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , 
     n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , 
     n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , 
     n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , 
     n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , 
     n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , 
     n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , 
     n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , 
     n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , 
     n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , 
     n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , 
     n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , 
     n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , 
     n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , 
     n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , 
     n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , 
     n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , 
     n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , 
     n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , 
     n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , 
     n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , 
     n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , 
     n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , 
     n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , 
     n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , 
     n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , 
     n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , 
     n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , 
     n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , 
     n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , 
     n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , 
     n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , 
     n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , 
     n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , 
     n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , 
     n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , 
     n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , 
     n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , 
     n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , 
     n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , 
     n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , 
     n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , 
     n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , 
     n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , 
     n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , 
     n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , 
     n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , 
     n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , 
     n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , 
     n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , 
     n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , 
     n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , 
     n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , 
     n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , 
     n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , 
     n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , 
     n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , 
     n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , 
     n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , 
     n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , 
     n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , 
     n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , 
     n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , 
     n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , 
     n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , 
     n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , 
     n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , 
     n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , 
     n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , 
     n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , 
     n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , 
     n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , 
     n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , 
     n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , 
     n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , 
     n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , 
     n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , 
     n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , 
     n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , 
     n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , 
     n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , 
     n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , 
     n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , 
     n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , 
     n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , 
     n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , 
     n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , 
     n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , 
     n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , 
     n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , 
     n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , 
     n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , 
     n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , 
     n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , 
     n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , 
     n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , 
     n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , 
     n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , 
     n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , 
     n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , 
     n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , 
     n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , 
     n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , 
     n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , 
     n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , 
     n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , 
     n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , 
     n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , 
     n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , 
     n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , 
     n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , 
     n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , 
     n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , 
     n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , 
     n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , 
     n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , 
     n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , 
     n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , 
     n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , 
     n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , 
     n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , 
     n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , 
     n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , 
     n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , 
     n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , 
     n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , 
     n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , 
     n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , 
     n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , 
     n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , 
     n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , 
     n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , 
     n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , 
     n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , 
     n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , 
     n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , 
     n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , 
     n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , 
     n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , 
     n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , 
     n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , 
     n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , 
     n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , 
     n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , 
     n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , 
     n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , 
     n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , 
     n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , 
     n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , 
     n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , 
     n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , 
     n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , 
     n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , 
     n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , 
     n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , 
     n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , 
     n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , 
     n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , 
     n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , 
     n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , 
     n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , 
     n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , 
     n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , 
     n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , 
     n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , 
     n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , 
     n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , 
     n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , 
     n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , 
     n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , 
     n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , 
     n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , 
     n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , 
     n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , 
     n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , 
     n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , 
     n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , 
     n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , 
     n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , 
     n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , 
     n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , 
     n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , 
     n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , 
     n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , 
     n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , 
     n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , 
     n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , 
     n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , 
     n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , 
     n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , 
     n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , 
     n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , 
     n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , 
     n3593 , n3594 , n3595 , n3596 ;
buf ( n513 , n3573 );
buf ( n515 , n3587 );
buf ( n512 , n3591 );
buf ( n516 , n3594 );
buf ( n514 , n3596 );
buf ( n1036 , n244 );
buf ( n1037 , n312 );
buf ( n1038 , n489 );
buf ( n1039 , n494 );
buf ( n1040 , n55 );
buf ( n1041 , n213 );
buf ( n1042 , n68 );
buf ( n1043 , n298 );
buf ( n1044 , n77 );
buf ( n1045 , n38 );
buf ( n1046 , n32 );
buf ( n1047 , n448 );
buf ( n1048 , n388 );
buf ( n1049 , n360 );
buf ( n1050 , n156 );
buf ( n1051 , n286 );
buf ( n1052 , n405 );
buf ( n1053 , n209 );
buf ( n1054 , n472 );
buf ( n1055 , n33 );
buf ( n1056 , n397 );
buf ( n1057 , n101 );
buf ( n1058 , n357 );
buf ( n1059 , n289 );
buf ( n1060 , n498 );
buf ( n1061 , n164 );
buf ( n1062 , n115 );
buf ( n1063 , n103 );
buf ( n1064 , n67 );
buf ( n1065 , n139 );
buf ( n1066 , n121 );
buf ( n1067 , n358 );
buf ( n1068 , n483 );
buf ( n1069 , n131 );
buf ( n1070 , n95 );
buf ( n1071 , n74 );
buf ( n1072 , n221 );
buf ( n1073 , n49 );
buf ( n1074 , n185 );
buf ( n1075 , n206 );
buf ( n1076 , n379 );
buf ( n1077 , n464 );
buf ( n1078 , n75 );
buf ( n1079 , n136 );
buf ( n1080 , n184 );
buf ( n1081 , n203 );
buf ( n1082 , n278 );
buf ( n1083 , n153 );
buf ( n1084 , n178 );
buf ( n1085 , n159 );
buf ( n1086 , n283 );
buf ( n1087 , n255 );
buf ( n1088 , n404 );
buf ( n1089 , n275 );
buf ( n1090 , n353 );
buf ( n1091 , n73 );
buf ( n1092 , n105 );
buf ( n1093 , n462 );
buf ( n1094 , n102 );
buf ( n1095 , n120 );
buf ( n1096 , n249 );
buf ( n1097 , n441 );
buf ( n1098 , n402 );
buf ( n1099 , n225 );
buf ( n1100 , n238 );
buf ( n1101 , n455 );
buf ( n1102 , n363 );
buf ( n1103 , n147 );
buf ( n1104 , n224 );
buf ( n1105 , n128 );
buf ( n1106 , n52 );
buf ( n1107 , n108 );
buf ( n1108 , n486 );
buf ( n1109 , n471 );
buf ( n1110 , n356 );
buf ( n1111 , n276 );
buf ( n1112 , n454 );
buf ( n1113 , n9 );
buf ( n1114 , n281 );
buf ( n1115 , n180 );
buf ( n1116 , n324 );
buf ( n1117 , n340 );
buf ( n1118 , n309 );
buf ( n1119 , n337 );
buf ( n1120 , n484 );
buf ( n1121 , n291 );
buf ( n1122 , n349 );
buf ( n1123 , n375 );
buf ( n1124 , n325 );
buf ( n1125 , n195 );
buf ( n1126 , n425 );
buf ( n1127 , n507 );
buf ( n1128 , n461 );
buf ( n1129 , n460 );
buf ( n1130 , n348 );
buf ( n1131 , n328 );
buf ( n1132 , n467 );
buf ( n1133 , n65 );
buf ( n1134 , n506 );
buf ( n1135 , n208 );
buf ( n1136 , n273 );
buf ( n1137 , n352 );
buf ( n1138 , n84 );
buf ( n1139 , n230 );
buf ( n1140 , n100 );
buf ( n1141 , n346 );
buf ( n1142 , n362 );
buf ( n1143 , n177 );
buf ( n1144 , n509 );
buf ( n1145 , n192 );
buf ( n1146 , n24 );
buf ( n1147 , n22 );
buf ( n1148 , n158 );
buf ( n1149 , n92 );
buf ( n1150 , n411 );
buf ( n1151 , n343 );
buf ( n1152 , n62 );
buf ( n1153 , n459 );
buf ( n1154 , n126 );
buf ( n1155 , n111 );
buf ( n1156 , n58 );
buf ( n1157 , n439 );
buf ( n1158 , n313 );
buf ( n1159 , n130 );
buf ( n1160 , n37 );
buf ( n1161 , n345 );
buf ( n1162 , n135 );
buf ( n1163 , n475 );
buf ( n1164 , n223 );
buf ( n1165 , n233 );
buf ( n1166 , n389 );
buf ( n1167 , n393 );
buf ( n1168 , n236 );
buf ( n1169 , n143 );
buf ( n1170 , n216 );
buf ( n1171 , n430 );
buf ( n1172 , n399 );
buf ( n1173 , n28 );
buf ( n1174 , n378 );
buf ( n1175 , n350 );
buf ( n1176 , n23 );
buf ( n1177 , n246 );
buf ( n1178 , n320 );
buf ( n1179 , n499 );
buf ( n1180 , n112 );
buf ( n1181 , n410 );
buf ( n1182 , n160 );
buf ( n1183 , n386 );
buf ( n1184 , n418 );
buf ( n1185 , n194 );
buf ( n1186 , n318 );
buf ( n1187 , n432 );
buf ( n1188 , n219 );
buf ( n1189 , n477 );
buf ( n1190 , n170 );
buf ( n1191 , n282 );
buf ( n1192 , n331 );
buf ( n1193 , n372 );
buf ( n1194 , n505 );
buf ( n1195 , n6 );
buf ( n1196 , n14 );
buf ( n1197 , n271 );
buf ( n1198 , n168 );
buf ( n1199 , n248 );
buf ( n1200 , n149 );
buf ( n1201 , n0 );
buf ( n1202 , n382 );
buf ( n1203 , n447 );
buf ( n1204 , n56 );
buf ( n1205 , n110 );
buf ( n1206 , n162 );
buf ( n1207 , n150 );
buf ( n1208 , n123 );
buf ( n1209 , n390 );
buf ( n1210 , n323 );
buf ( n1211 , n371 );
buf ( n1212 , n303 );
buf ( n1213 , n34 );
buf ( n1214 , n480 );
buf ( n1215 , n127 );
buf ( n1216 , n429 );
buf ( n1217 , n338 );
buf ( n1218 , n25 );
buf ( n1219 , n82 );
buf ( n1220 , n215 );
buf ( n1221 , n502 );
buf ( n1222 , n450 );
buf ( n1223 , n335 );
buf ( n1224 , n272 );
buf ( n1225 , n446 );
buf ( n1226 , n187 );
buf ( n1227 , n161 );
buf ( n1228 , n361 );
buf ( n1229 , n99 );
buf ( n1230 , n302 );
buf ( n1231 , n334 );
buf ( n1232 , n85 );
buf ( n1233 , n129 );
buf ( n1234 , n481 );
buf ( n1235 , n417 );
buf ( n1236 , n394 );
buf ( n1237 , n193 );
buf ( n1238 , n125 );
buf ( n1239 , n152 );
buf ( n1240 , n88 );
buf ( n1241 , n332 );
buf ( n1242 , n339 );
buf ( n1243 , n122 );
buf ( n1244 , n252 );
buf ( n1245 , n280 );
buf ( n1246 , n458 );
buf ( n1247 , n148 );
buf ( n1248 , n500 );
buf ( n1249 , n235 );
buf ( n1250 , n431 );
buf ( n1251 , n401 );
buf ( n1252 , n277 );
buf ( n1253 , n46 );
buf ( n1254 , n327 );
buf ( n1255 , n189 );
buf ( n1256 , n501 );
buf ( n1257 , n510 );
buf ( n1258 , n40 );
buf ( n1259 , n307 );
buf ( n1260 , n262 );
buf ( n1261 , n300 );
buf ( n1262 , n419 );
buf ( n1263 , n463 );
buf ( n1264 , n17 );
buf ( n1265 , n493 );
buf ( n1266 , n54 );
buf ( n1267 , n288 );
buf ( n1268 , n310 );
buf ( n1269 , n241 );
buf ( n1270 , n336 );
buf ( n1271 , n87 );
buf ( n1272 , n228 );
buf ( n1273 , n78 );
buf ( n1274 , n354 );
buf ( n1275 , n59 );
buf ( n1276 , n265 );
buf ( n1277 , n19 );
buf ( n1278 , n377 );
buf ( n1279 , n412 );
buf ( n1280 , n231 );
buf ( n1281 , n465 );
buf ( n1282 , n250 );
buf ( n1283 , n176 );
buf ( n1284 , n299 );
buf ( n1285 , n259 );
buf ( n1286 , n169 );
buf ( n1287 , n466 );
buf ( n1288 , n31 );
buf ( n1289 , n452 );
buf ( n1290 , n145 );
buf ( n1291 , n47 );
buf ( n1292 , n444 );
buf ( n1293 , n69 );
buf ( n1294 , n5 );
buf ( n1295 , n89 );
buf ( n1296 , n197 );
buf ( n1297 , n98 );
buf ( n1298 , n453 );
buf ( n1299 , n175 );
buf ( n1300 , n217 );
buf ( n1301 , n60 );
buf ( n1302 , n204 );
buf ( n1303 , n293 );
buf ( n1304 , n457 );
buf ( n1305 , n26 );
buf ( n1306 , n306 );
buf ( n1307 , n406 );
buf ( n1308 , n497 );
buf ( n1309 , n391 );
buf ( n1310 , n1 );
buf ( n1311 , n269 );
buf ( n1312 , n44 );
buf ( n1313 , n434 );
buf ( n1314 , n30 );
buf ( n1315 , n474 );
buf ( n1316 , n190 );
buf ( n1317 , n21 );
buf ( n1318 , n72 );
buf ( n1319 , n71 );
buf ( n1320 , n267 );
buf ( n1321 , n119 );
buf ( n1322 , n266 );
buf ( n1323 , n373 );
buf ( n1324 , n487 );
buf ( n1325 , n482 );
buf ( n1326 , n91 );
buf ( n1327 , n146 );
buf ( n1328 , n124 );
buf ( n1329 , n45 );
buf ( n1330 , n329 );
buf ( n1331 , n50 );
buf ( n1332 , n294 );
buf ( n1333 , n254 );
buf ( n1334 , n76 );
buf ( n1335 , n400 );
buf ( n1336 , n261 );
buf ( n1337 , n94 );
buf ( n1338 , n420 );
buf ( n1339 , n264 );
buf ( n1340 , n70 );
buf ( n1341 , n133 );
buf ( n1342 , n199 );
buf ( n1343 , n20 );
buf ( n1344 , n290 );
buf ( n1345 , n93 );
buf ( n1346 , n202 );
buf ( n1347 , n315 );
buf ( n1348 , n468 );
buf ( n1349 , n86 );
buf ( n1350 , n268 );
buf ( n1351 , n495 );
buf ( n1352 , n182 );
buf ( n1353 , n27 );
buf ( n1354 , n220 );
buf ( n1355 , n344 );
buf ( n1356 , n240 );
buf ( n1357 , n81 );
buf ( n1358 , n232 );
buf ( n1359 , n508 );
buf ( n1360 , n2 );
buf ( n1361 , n41 );
buf ( n1362 , n186 );
buf ( n1363 , n351 );
buf ( n1364 , n179 );
buf ( n1365 , n296 );
buf ( n1366 , n243 );
buf ( n1367 , n96 );
buf ( n1368 , n35 );
buf ( n1369 , n287 );
buf ( n1370 , n29 );
buf ( n1371 , n414 );
buf ( n1372 , n415 );
buf ( n1373 , n214 );
buf ( n1374 , n284 );
buf ( n1375 , n395 );
buf ( n1376 , n201 );
buf ( n1377 , n4 );
buf ( n1378 , n333 );
buf ( n1379 , n387 );
buf ( n1380 , n237 );
buf ( n1381 , n392 );
buf ( n1382 , n416 );
buf ( n1383 , n8 );
buf ( n1384 , n188 );
buf ( n1385 , n53 );
buf ( n1386 , n478 );
buf ( n1387 , n359 );
buf ( n1388 , n171 );
buf ( n1389 , n476 );
buf ( n1390 , n163 );
buf ( n1391 , n449 );
buf ( n1392 , n191 );
buf ( n1393 , n227 );
buf ( n1394 , n492 );
buf ( n1395 , n297 );
buf ( n1396 , n245 );
buf ( n1397 , n106 );
buf ( n1398 , n365 );
buf ( n1399 , n274 );
buf ( n1400 , n316 );
buf ( n1401 , n116 );
buf ( n1402 , n157 );
buf ( n1403 , n451 );
buf ( n1404 , n376 );
buf ( n1405 , n155 );
buf ( n1406 , n364 );
buf ( n1407 , n381 );
buf ( n1408 , n426 );
buf ( n1409 , n196 );
buf ( n1410 , n384 );
buf ( n1411 , n256 );
buf ( n1412 , n260 );
buf ( n1413 , n317 );
buf ( n1414 , n270 );
buf ( n1415 , n314 );
buf ( n1416 , n311 );
buf ( n1417 , n183 );
buf ( n1418 , n39 );
buf ( n1419 , n366 );
buf ( n1420 , n212 );
buf ( n1421 , n421 );
buf ( n1422 , n427 );
buf ( n1423 , n239 );
buf ( n1424 , n11 );
buf ( n1425 , n326 );
buf ( n1426 , n369 );
buf ( n1427 , n166 );
buf ( n1428 , n403 );
buf ( n1429 , n470 );
buf ( n1430 , n205 );
buf ( n1431 , n422 );
buf ( n1432 , n174 );
buf ( n1433 , n118 );
buf ( n1434 , n198 );
buf ( n1435 , n57 );
buf ( n1436 , n7 );
buf ( n1437 , n10 );
buf ( n1438 , n251 );
buf ( n1439 , n511 );
buf ( n1440 , n247 );
buf ( n1441 , n42 );
buf ( n1442 , n36 );
buf ( n1443 , n222 );
buf ( n1444 , n367 );
buf ( n1445 , n144 );
buf ( n1446 , n137 );
buf ( n1447 , n134 );
buf ( n1448 , n396 );
buf ( n1449 , n43 );
buf ( n1450 , n321 );
buf ( n1451 , n503 );
buf ( n1452 , n66 );
buf ( n1453 , n479 );
buf ( n1454 , n242 );
buf ( n1455 , n330 );
buf ( n1456 , n107 );
buf ( n1457 , n12 );
buf ( n1458 , n305 );
buf ( n1459 , n490 );
buf ( n1460 , n423 );
buf ( n1461 , n368 );
buf ( n1462 , n117 );
buf ( n1463 , n90 );
buf ( n1464 , n370 );
buf ( n1465 , n342 );
buf ( n1466 , n16 );
buf ( n1467 , n3 );
buf ( n1468 , n109 );
buf ( n1469 , n485 );
buf ( n1470 , n341 );
buf ( n1471 , n295 );
buf ( n1472 , n442 );
buf ( n1473 , n104 );
buf ( n1474 , n473 );
buf ( n1475 , n285 );
buf ( n1476 , n200 );
buf ( n1477 , n140 );
buf ( n1478 , n63 );
buf ( n1479 , n436 );
buf ( n1480 , n438 );
buf ( n1481 , n51 );
buf ( n1482 , n181 );
buf ( n1483 , n226 );
buf ( n1484 , n173 );
buf ( n1485 , n165 );
buf ( n1486 , n263 );
buf ( n1487 , n138 );
buf ( n1488 , n456 );
buf ( n1489 , n304 );
buf ( n1490 , n433 );
buf ( n1491 , n409 );
buf ( n1492 , n218 );
buf ( n1493 , n408 );
buf ( n1494 , n13 );
buf ( n1495 , n61 );
buf ( n1496 , n79 );
buf ( n1497 , n437 );
buf ( n1498 , n234 );
buf ( n1499 , n151 );
buf ( n1500 , n229 );
buf ( n1501 , n258 );
buf ( n1502 , n440 );
buf ( n1503 , n413 );
buf ( n1504 , n383 );
buf ( n1505 , n319 );
buf ( n1506 , n301 );
buf ( n1507 , n380 );
buf ( n1508 , n374 );
buf ( n1509 , n64 );
buf ( n1510 , n424 );
buf ( n1511 , n83 );
buf ( n1512 , n488 );
buf ( n1513 , n496 );
buf ( n1514 , n141 );
buf ( n1515 , n211 );
buf ( n1516 , n15 );
buf ( n1517 , n308 );
buf ( n1518 , n172 );
buf ( n1519 , n398 );
buf ( n1520 , n167 );
buf ( n1521 , n132 );
buf ( n1522 , n253 );
buf ( n1523 , n18 );
buf ( n1524 , n322 );
buf ( n1525 , n114 );
buf ( n1526 , n48 );
buf ( n1527 , n347 );
buf ( n1528 , n154 );
buf ( n1529 , n97 );
buf ( n1530 , n385 );
buf ( n1531 , n292 );
buf ( n1532 , n279 );
buf ( n1533 , n428 );
buf ( n1534 , n445 );
buf ( n1535 , n355 );
buf ( n1536 , n113 );
buf ( n1537 , n491 );
buf ( n1538 , n207 );
buf ( n1539 , n80 );
buf ( n1540 , n504 );
buf ( n1541 , n435 );
buf ( n1542 , n469 );
buf ( n1543 , n142 );
buf ( n1544 , n407 );
buf ( n1545 , n210 );
buf ( n1546 , n257 );
buf ( n1547 , n443 );
and ( n1548 , n1039 , n1167 );
not ( n1549 , n1039 );
not ( n1550 , n1167 );
and ( n1551 , n1549 , n1550 );
nor ( n1552 , n1548 , n1551 );
and ( n1553 , n1295 , n1423 );
not ( n1554 , n1295 );
not ( n1555 , n1423 );
and ( n1556 , n1554 , n1555 );
nor ( n1557 , n1553 , n1556 );
nand ( n1558 , n1552 , n1557 );
not ( n1559 , n1558 );
nor ( n1560 , n1557 , n1552 );
or ( n1561 , n1559 , n1560 );
and ( n1562 , n1038 , n1166 );
not ( n1563 , n1038 );
not ( n1564 , n1166 );
and ( n1565 , n1563 , n1564 );
nor ( n1566 , n1562 , n1565 );
xor ( n1567 , n1294 , n1422 );
not ( n1568 , n1567 );
and ( n1569 , n1566 , n1568 );
not ( n1570 , n1566 );
and ( n1571 , n1570 , n1567 );
nor ( n1572 , n1569 , n1571 );
nand ( n1573 , n1561 , n1572 );
and ( n1574 , n1165 , n1293 );
not ( n1575 , n1165 );
not ( n1576 , n1293 );
and ( n1577 , n1575 , n1576 );
nor ( n1578 , n1574 , n1577 );
and ( n1579 , n1037 , n1421 );
not ( n1580 , n1037 );
not ( n1581 , n1421 );
and ( n1582 , n1580 , n1581 );
nor ( n1583 , n1579 , n1582 );
nand ( n1584 , n1578 , n1583 );
not ( n1585 , n1584 );
nor ( n1586 , n1583 , n1578 );
or ( n1587 , n1585 , n1586 );
and ( n1588 , n1036 , n1164 );
not ( n1589 , n1036 );
not ( n1590 , n1164 );
and ( n1591 , n1589 , n1590 );
nor ( n1592 , n1588 , n1591 );
xor ( n1593 , n1292 , n1420 );
not ( n1594 , n1593 );
and ( n1595 , n1592 , n1594 );
not ( n1596 , n1592 );
and ( n1597 , n1596 , n1593 );
nor ( n1598 , n1595 , n1597 );
nand ( n1599 , n1587 , n1598 );
nor ( n1600 , n1573 , n1599 );
and ( n1601 , n1299 , n1427 );
not ( n1602 , n1299 );
not ( n1603 , n1427 );
and ( n1604 , n1602 , n1603 );
nor ( n1605 , n1601 , n1604 );
not ( n1606 , n1043 );
and ( n1607 , n1171 , n1606 );
not ( n1608 , n1171 );
and ( n1609 , n1608 , n1043 );
nor ( n1610 , n1607 , n1609 );
and ( n1611 , n1605 , n1610 );
not ( n1612 , n1605 );
not ( n1613 , n1610 );
and ( n1614 , n1612 , n1613 );
nor ( n1615 , n1611 , n1614 );
and ( n1616 , n1042 , n1170 );
not ( n1617 , n1042 );
not ( n1618 , n1170 );
and ( n1619 , n1617 , n1618 );
nor ( n1620 , n1616 , n1619 );
not ( n1621 , n1620 );
and ( n1622 , n1298 , n1426 );
not ( n1623 , n1298 );
not ( n1624 , n1426 );
and ( n1625 , n1623 , n1624 );
nor ( n1626 , n1622 , n1625 );
not ( n1627 , n1626 );
or ( n1628 , n1621 , n1627 );
or ( n1629 , n1620 , n1626 );
nand ( n1630 , n1628 , n1629 );
nand ( n1631 , n1615 , n1630 );
and ( n1632 , n1040 , n1168 );
not ( n1633 , n1040 );
not ( n1634 , n1168 );
and ( n1635 , n1633 , n1634 );
nor ( n1636 , n1632 , n1635 );
and ( n1637 , n1296 , n1424 );
not ( n1638 , n1296 );
not ( n1639 , n1424 );
and ( n1640 , n1638 , n1639 );
nor ( n1641 , n1637 , n1640 );
not ( n1642 , n1641 );
and ( n1643 , n1636 , n1642 );
not ( n1644 , n1636 );
and ( n1645 , n1644 , n1641 );
nor ( n1646 , n1643 , n1645 );
and ( n1647 , n1169 , n1297 );
not ( n1648 , n1169 );
not ( n1649 , n1297 );
and ( n1650 , n1648 , n1649 );
nor ( n1651 , n1647 , n1650 );
and ( n1652 , n1041 , n1425 );
not ( n1653 , n1041 );
not ( n1654 , n1425 );
and ( n1655 , n1653 , n1654 );
nor ( n1656 , n1652 , n1655 );
not ( n1657 , n1656 );
and ( n1658 , n1651 , n1657 );
not ( n1659 , n1651 );
and ( n1660 , n1659 , n1656 );
nor ( n1661 , n1658 , n1660 );
nand ( n1662 , n1646 , n1661 );
nor ( n1663 , n1631 , n1662 );
nand ( n1664 , n1600 , n1663 );
and ( n1665 , n1175 , n1303 );
not ( n1666 , n1175 );
not ( n1667 , n1303 );
and ( n1668 , n1666 , n1667 );
nor ( n1669 , n1665 , n1668 );
and ( n1670 , n1047 , n1431 );
not ( n1671 , n1047 );
not ( n1672 , n1431 );
and ( n1673 , n1671 , n1672 );
nor ( n1674 , n1670 , n1673 );
nand ( n1675 , n1669 , n1674 );
not ( n1676 , n1675 );
nor ( n1677 , n1674 , n1669 );
or ( n1678 , n1676 , n1677 );
and ( n1679 , n1046 , n1174 );
not ( n1680 , n1046 );
not ( n1681 , n1174 );
and ( n1682 , n1680 , n1681 );
nor ( n1683 , n1679 , n1682 );
xor ( n1684 , n1302 , n1430 );
not ( n1685 , n1684 );
and ( n1686 , n1683 , n1685 );
not ( n1687 , n1683 );
and ( n1688 , n1687 , n1684 );
nor ( n1689 , n1686 , n1688 );
nand ( n1690 , n1678 , n1689 );
and ( n1691 , n1045 , n1173 );
not ( n1692 , n1045 );
not ( n1693 , n1173 );
and ( n1694 , n1692 , n1693 );
nor ( n1695 , n1691 , n1694 );
and ( n1696 , n1301 , n1429 );
not ( n1697 , n1301 );
not ( n1698 , n1429 );
and ( n1699 , n1697 , n1698 );
nor ( n1700 , n1696 , n1699 );
nand ( n1701 , n1695 , n1700 );
not ( n1702 , n1701 );
not ( n1703 , n1700 );
and ( n1704 , n1045 , n1173 );
not ( n1705 , n1045 );
and ( n1706 , n1705 , n1693 );
nor ( n1707 , n1704 , n1706 );
not ( n1708 , n1707 );
nand ( n1709 , n1703 , n1708 );
not ( n1710 , n1709 );
or ( n1711 , n1702 , n1710 );
not ( n1712 , n1428 );
nand ( n1713 , n1712 , n1044 );
not ( n1714 , n1044 );
nand ( n1715 , n1714 , n1428 );
nand ( n1716 , n1713 , n1715 );
and ( n1717 , n1172 , n1300 );
not ( n1718 , n1172 );
not ( n1719 , n1300 );
and ( n1720 , n1718 , n1719 );
nor ( n1721 , n1717 , n1720 );
or ( n1722 , n1716 , n1721 );
nand ( n1723 , n1714 , n1428 );
not ( n1724 , n1723 );
not ( n1725 , n1713 );
or ( n1726 , n1724 , n1725 );
nand ( n1727 , n1726 , n1721 );
nand ( n1728 , n1722 , n1727 );
nand ( n1729 , n1711 , n1728 );
nor ( n1730 , n1690 , n1729 );
and ( n1731 , n1178 , n1306 );
not ( n1732 , n1178 );
not ( n1733 , n1306 );
and ( n1734 , n1732 , n1733 );
nor ( n1735 , n1731 , n1734 );
and ( n1736 , n1050 , n1434 );
not ( n1737 , n1050 );
not ( n1738 , n1434 );
and ( n1739 , n1737 , n1738 );
nor ( n1740 , n1736 , n1739 );
not ( n1741 , n1740 );
and ( n1742 , n1735 , n1741 );
not ( n1743 , n1735 );
and ( n1744 , n1743 , n1740 );
nor ( n1745 , n1742 , n1744 );
and ( n1746 , n1051 , n1179 );
not ( n1747 , n1051 );
not ( n1748 , n1179 );
and ( n1749 , n1747 , n1748 );
nor ( n1750 , n1746 , n1749 );
and ( n1751 , n1307 , n1435 );
not ( n1752 , n1307 );
not ( n1753 , n1435 );
and ( n1754 , n1752 , n1753 );
nor ( n1755 , n1751 , n1754 );
not ( n1756 , n1755 );
and ( n1757 , n1750 , n1756 );
not ( n1758 , n1750 );
and ( n1759 , n1758 , n1755 );
nor ( n1760 , n1757 , n1759 );
nand ( n1761 , n1745 , n1760 );
not ( n1762 , n1432 );
not ( n1763 , n1304 );
and ( n1764 , n1762 , n1763 );
and ( n1765 , n1304 , n1432 );
nor ( n1766 , n1764 , n1765 );
and ( n1767 , n1048 , n1176 );
not ( n1768 , n1048 );
not ( n1769 , n1176 );
and ( n1770 , n1768 , n1769 );
nor ( n1771 , n1767 , n1770 );
or ( n1772 , n1766 , n1771 );
and ( n1773 , n1304 , n1432 );
not ( n1774 , n1304 );
and ( n1775 , n1774 , n1762 );
nor ( n1776 , n1773 , n1775 );
nand ( n1777 , n1776 , n1771 );
nand ( n1778 , n1772 , n1777 );
and ( n1779 , n1305 , n1433 );
not ( n1780 , n1305 );
not ( n1781 , n1433 );
and ( n1782 , n1780 , n1781 );
nor ( n1783 , n1779 , n1782 );
and ( n1784 , n1049 , n1177 );
not ( n1785 , n1049 );
not ( n1786 , n1177 );
and ( n1787 , n1785 , n1786 );
nor ( n1788 , n1784 , n1787 );
not ( n1789 , n1788 );
and ( n1790 , n1783 , n1789 );
not ( n1791 , n1783 );
and ( n1792 , n1791 , n1788 );
nor ( n1793 , n1790 , n1792 );
nand ( n1794 , n1778 , n1793 );
nor ( n1795 , n1761 , n1794 );
nand ( n1796 , n1730 , n1795 );
nor ( n1797 , n1664 , n1796 );
and ( n1798 , n1311 , n1439 );
not ( n1799 , n1311 );
not ( n1800 , n1439 );
and ( n1801 , n1799 , n1800 );
nor ( n1802 , n1798 , n1801 );
not ( n1803 , n1802 );
and ( n1804 , n1055 , n1183 );
not ( n1805 , n1055 );
not ( n1806 , n1183 );
and ( n1807 , n1805 , n1806 );
nor ( n1808 , n1804 , n1807 );
not ( n1809 , n1808 );
or ( n1810 , n1803 , n1809 );
or ( n1811 , n1808 , n1802 );
nand ( n1812 , n1810 , n1811 );
not ( n1813 , n1054 );
and ( n1814 , n1438 , n1813 );
not ( n1815 , n1438 );
and ( n1816 , n1815 , n1054 );
nor ( n1817 , n1814 , n1816 );
and ( n1818 , n1182 , n1310 );
not ( n1819 , n1182 );
not ( n1820 , n1310 );
and ( n1821 , n1819 , n1820 );
nor ( n1822 , n1818 , n1821 );
and ( n1823 , n1817 , n1822 );
not ( n1824 , n1817 );
not ( n1825 , n1822 );
and ( n1826 , n1824 , n1825 );
nor ( n1827 , n1823 , n1826 );
nand ( n1828 , n1812 , n1827 );
and ( n1829 , n1181 , n1309 );
not ( n1830 , n1181 );
not ( n1831 , n1309 );
and ( n1832 , n1830 , n1831 );
nor ( n1833 , n1829 , n1832 );
and ( n1834 , n1053 , n1437 );
not ( n1835 , n1053 );
not ( n1836 , n1437 );
and ( n1837 , n1835 , n1836 );
nor ( n1838 , n1834 , n1837 );
not ( n1839 , n1838 );
and ( n1840 , n1833 , n1839 );
not ( n1841 , n1833 );
and ( n1842 , n1841 , n1838 );
nor ( n1843 , n1840 , n1842 );
and ( n1844 , n1052 , n1180 );
not ( n1845 , n1052 );
not ( n1846 , n1180 );
and ( n1847 , n1845 , n1846 );
nor ( n1848 , n1844 , n1847 );
xor ( n1849 , n1308 , n1436 );
not ( n1850 , n1849 );
and ( n1851 , n1848 , n1850 );
not ( n1852 , n1848 );
and ( n1853 , n1852 , n1849 );
nor ( n1854 , n1851 , n1853 );
nand ( n1855 , n1843 , n1854 );
nor ( n1856 , n1828 , n1855 );
and ( n1857 , n1313 , n1441 );
not ( n1858 , n1313 );
not ( n1859 , n1441 );
and ( n1860 , n1858 , n1859 );
nor ( n1861 , n1857 , n1860 );
and ( n1862 , n1057 , n1185 );
not ( n1863 , n1057 );
not ( n1864 , n1185 );
and ( n1865 , n1863 , n1864 );
nor ( n1866 , n1862 , n1865 );
nand ( n1867 , n1861 , n1866 );
not ( n1868 , n1867 );
nor ( n1869 , n1861 , n1866 );
or ( n1870 , n1868 , n1869 );
and ( n1871 , n1184 , n1312 );
not ( n1872 , n1184 );
not ( n1873 , n1312 );
and ( n1874 , n1872 , n1873 );
nor ( n1875 , n1871 , n1874 );
xor ( n1876 , n1056 , n1440 );
not ( n1877 , n1876 );
and ( n1878 , n1875 , n1877 );
not ( n1879 , n1875 );
and ( n1880 , n1879 , n1876 );
nor ( n1881 , n1878 , n1880 );
nand ( n1882 , n1870 , n1881 );
and ( n1883 , n1059 , n1187 );
not ( n1884 , n1059 );
not ( n1885 , n1187 );
and ( n1886 , n1884 , n1885 );
nor ( n1887 , n1883 , n1886 );
and ( n1888 , n1315 , n1443 );
not ( n1889 , n1315 );
not ( n1890 , n1443 );
and ( n1891 , n1889 , n1890 );
nor ( n1892 , n1888 , n1891 );
not ( n1893 , n1892 );
and ( n1894 , n1887 , n1893 );
not ( n1895 , n1887 );
and ( n1896 , n1895 , n1892 );
nor ( n1897 , n1894 , n1896 );
and ( n1898 , n1186 , n1314 );
not ( n1899 , n1186 );
not ( n1900 , n1314 );
and ( n1901 , n1899 , n1900 );
nor ( n1902 , n1898 , n1901 );
xor ( n1903 , n1058 , n1442 );
not ( n1904 , n1903 );
and ( n1905 , n1902 , n1904 );
not ( n1906 , n1902 );
and ( n1907 , n1906 , n1903 );
nor ( n1908 , n1905 , n1907 );
nand ( n1909 , n1897 , n1908 );
nor ( n1910 , n1882 , n1909 );
nand ( n1911 , n1856 , n1910 );
and ( n1912 , n1195 , n1323 );
not ( n1913 , n1195 );
not ( n1914 , n1323 );
and ( n1915 , n1913 , n1914 );
nor ( n1916 , n1912 , n1915 );
and ( n1917 , n1067 , n1451 );
not ( n1918 , n1067 );
not ( n1919 , n1451 );
and ( n1920 , n1918 , n1919 );
nor ( n1921 , n1917 , n1920 );
nand ( n1922 , n1916 , n1921 );
not ( n1923 , n1922 );
nor ( n1924 , n1921 , n1916 );
or ( n1925 , n1923 , n1924 );
and ( n1926 , n1066 , n1194 );
not ( n1927 , n1066 );
not ( n1928 , n1194 );
and ( n1929 , n1927 , n1928 );
nor ( n1930 , n1926 , n1929 );
xor ( n1931 , n1322 , n1450 );
not ( n1932 , n1931 );
and ( n1933 , n1930 , n1932 );
not ( n1934 , n1930 );
and ( n1935 , n1934 , n1931 );
nor ( n1936 , n1933 , n1935 );
nand ( n1937 , n1925 , n1936 );
and ( n1938 , n1193 , n1321 );
not ( n1939 , n1193 );
not ( n1940 , n1321 );
and ( n1941 , n1939 , n1940 );
nor ( n1942 , n1938 , n1941 );
and ( n1943 , n1065 , n1449 );
not ( n1944 , n1065 );
not ( n1945 , n1449 );
and ( n1946 , n1944 , n1945 );
nor ( n1947 , n1943 , n1946 );
nand ( n1948 , n1942 , n1947 );
not ( n1949 , n1948 );
not ( n1950 , n1947 );
and ( n1951 , n1193 , n1321 );
not ( n1952 , n1193 );
and ( n1953 , n1952 , n1940 );
nor ( n1954 , n1951 , n1953 );
not ( n1955 , n1954 );
nand ( n1956 , n1950 , n1955 );
not ( n1957 , n1956 );
or ( n1958 , n1949 , n1957 );
not ( n1959 , n1448 );
nand ( n1960 , n1959 , n1320 );
not ( n1961 , n1320 );
nand ( n1962 , n1961 , n1448 );
nand ( n1963 , n1960 , n1962 );
and ( n1964 , n1064 , n1192 );
not ( n1965 , n1064 );
not ( n1966 , n1192 );
and ( n1967 , n1965 , n1966 );
nor ( n1968 , n1964 , n1967 );
or ( n1969 , n1963 , n1968 );
nand ( n1970 , n1961 , n1448 );
not ( n1971 , n1970 );
not ( n1972 , n1960 );
or ( n1973 , n1971 , n1972 );
nand ( n1974 , n1973 , n1968 );
nand ( n1975 , n1969 , n1974 );
nand ( n1976 , n1958 , n1975 );
nor ( n1977 , n1937 , n1976 );
and ( n1978 , n1191 , n1319 );
not ( n1979 , n1191 );
not ( n1980 , n1319 );
and ( n1981 , n1979 , n1980 );
nor ( n1982 , n1978 , n1981 );
and ( n1983 , n1063 , n1447 );
not ( n1984 , n1063 );
not ( n1985 , n1447 );
and ( n1986 , n1984 , n1985 );
nor ( n1987 , n1983 , n1986 );
not ( n1988 , n1987 );
and ( n1989 , n1982 , n1988 );
not ( n1990 , n1982 );
and ( n1991 , n1990 , n1987 );
nor ( n1992 , n1989 , n1991 );
xor ( n1993 , n1062 , n1446 );
xnor ( n1994 , n1190 , n1318 );
and ( n1995 , n1993 , n1994 );
not ( n1996 , n1993 );
xor ( n1997 , n1190 , n1318 );
and ( n1998 , n1996 , n1997 );
nor ( n1999 , n1995 , n1998 );
nand ( n2000 , n1992 , n1999 );
and ( n2001 , n1189 , n1317 );
not ( n2002 , n1189 );
not ( n2003 , n1317 );
and ( n2004 , n2002 , n2003 );
nor ( n2005 , n2001 , n2004 );
not ( n2006 , n1061 );
not ( n2007 , n1445 );
not ( n2008 , n2007 );
or ( n2009 , n2006 , n2008 );
not ( n2010 , n1061 );
nand ( n2011 , n2010 , n1445 );
nand ( n2012 , n2009 , n2011 );
or ( n2013 , n2005 , n2012 );
nand ( n2014 , n2007 , n1061 );
not ( n2015 , n2014 );
not ( n2016 , n2011 );
or ( n2017 , n2015 , n2016 );
and ( n2018 , n1189 , n1317 );
not ( n2019 , n1189 );
and ( n2020 , n2019 , n2003 );
nor ( n2021 , n2018 , n2020 );
nand ( n2022 , n2017 , n2021 );
nand ( n2023 , n2013 , n2022 );
not ( n2024 , n1444 );
and ( n2025 , n1316 , n2024 );
not ( n2026 , n1316 );
and ( n2027 , n2026 , n1444 );
nor ( n2028 , n2025 , n2027 );
and ( n2029 , n1060 , n1188 );
not ( n2030 , n1060 );
not ( n2031 , n1188 );
and ( n2032 , n2030 , n2031 );
nor ( n2033 , n2029 , n2032 );
and ( n2034 , n2028 , n2033 );
not ( n2035 , n2028 );
not ( n2036 , n1060 );
nand ( n2037 , n2036 , n2031 );
nand ( n2038 , n1188 , n1060 );
nand ( n2039 , n2037 , n2038 );
and ( n2040 , n2035 , n2039 );
nor ( n2041 , n2034 , n2040 );
nand ( n2042 , n2023 , n2041 );
nor ( n2043 , n2000 , n2042 );
nand ( n2044 , n1977 , n2043 );
nor ( n2045 , n1911 , n2044 );
nand ( n2046 , n1797 , n2045 );
and ( n2047 , n1202 , n1330 );
not ( n2048 , n1202 );
not ( n2049 , n1330 );
and ( n2050 , n2048 , n2049 );
nor ( n2051 , n2047 , n2050 );
and ( n2052 , n1074 , n1458 );
not ( n2053 , n1074 );
not ( n2054 , n1458 );
and ( n2055 , n2053 , n2054 );
nor ( n2056 , n2052 , n2055 );
not ( n2057 , n2056 );
and ( n2058 , n2051 , n2057 );
not ( n2059 , n2051 );
and ( n2060 , n2059 , n2056 );
nor ( n2061 , n2058 , n2060 );
and ( n2062 , n1203 , n1331 );
not ( n2063 , n1203 );
not ( n2064 , n1331 );
and ( n2065 , n2063 , n2064 );
nor ( n2066 , n2062 , n2065 );
and ( n2067 , n1075 , n1459 );
not ( n2068 , n1075 );
not ( n2069 , n1459 );
and ( n2070 , n2068 , n2069 );
nor ( n2071 , n2067 , n2070 );
not ( n2072 , n2071 );
and ( n2073 , n2066 , n2072 );
not ( n2074 , n2066 );
and ( n2075 , n2074 , n2071 );
nor ( n2076 , n2073 , n2075 );
nand ( n2077 , n2061 , n2076 );
not ( n2078 , n1072 );
and ( n2079 , n1456 , n2078 );
not ( n2080 , n1456 );
and ( n2081 , n2080 , n1072 );
nor ( n2082 , n2079 , n2081 );
and ( n2083 , n1200 , n1328 );
not ( n2084 , n1200 );
not ( n2085 , n1328 );
and ( n2086 , n2084 , n2085 );
nor ( n2087 , n2083 , n2086 );
and ( n2088 , n2082 , n2087 );
not ( n2089 , n2082 );
not ( n2090 , n2087 );
and ( n2091 , n2089 , n2090 );
nor ( n2092 , n2088 , n2091 );
and ( n2093 , n1073 , n1457 );
not ( n2094 , n1073 );
not ( n2095 , n1457 );
and ( n2096 , n2094 , n2095 );
nor ( n2097 , n2093 , n2096 );
and ( n2098 , n1201 , n1329 );
not ( n2099 , n1201 );
not ( n2100 , n1329 );
and ( n2101 , n2099 , n2100 );
nor ( n2102 , n2098 , n2101 );
not ( n2103 , n2102 );
and ( n2104 , n2097 , n2103 );
not ( n2105 , n2097 );
and ( n2106 , n2105 , n2102 );
nor ( n2107 , n2104 , n2106 );
nand ( n2108 , n2092 , n2107 );
nor ( n2109 , n2077 , n2108 );
and ( n2110 , n1071 , n1455 );
not ( n2111 , n1071 );
not ( n2112 , n1455 );
and ( n2113 , n2111 , n2112 );
nor ( n2114 , n2110 , n2113 );
and ( n2115 , n1199 , n1327 );
not ( n2116 , n1199 );
not ( n2117 , n1327 );
and ( n2118 , n2116 , n2117 );
nor ( n2119 , n2115 , n2118 );
not ( n2120 , n2119 );
and ( n2121 , n2114 , n2120 );
not ( n2122 , n2114 );
and ( n2123 , n2122 , n2119 );
nor ( n2124 , n2121 , n2123 );
and ( n2125 , n1198 , n1326 );
not ( n2126 , n1198 );
not ( n2127 , n1326 );
and ( n2128 , n2126 , n2127 );
nor ( n2129 , n2125 , n2128 );
xor ( n2130 , n1070 , n1454 );
not ( n2131 , n2130 );
and ( n2132 , n2129 , n2131 );
not ( n2133 , n2129 );
and ( n2134 , n2133 , n2130 );
nor ( n2135 , n2132 , n2134 );
nand ( n2136 , n2124 , n2135 );
and ( n2137 , n1453 , n1325 );
not ( n2138 , n1453 );
not ( n2139 , n1325 );
and ( n2140 , n2138 , n2139 );
nor ( n2141 , n2137 , n2140 );
and ( n2142 , n1069 , n1197 );
not ( n2143 , n1069 );
not ( n2144 , n1197 );
and ( n2145 , n2143 , n2144 );
nor ( n2146 , n2142 , n2145 );
nand ( n2147 , n2141 , n2146 );
not ( n2148 , n2147 );
not ( n2149 , n2141 );
not ( n2150 , n2144 );
not ( n2151 , n1069 );
and ( n2152 , n2150 , n2151 );
and ( n2153 , n2144 , n1069 );
nor ( n2154 , n2152 , n2153 );
nand ( n2155 , n2149 , n2154 );
not ( n2156 , n2155 );
or ( n2157 , n2148 , n2156 );
not ( n2158 , n1324 );
not ( n2159 , n1452 );
not ( n2160 , n2159 );
or ( n2161 , n2158 , n2160 );
not ( n2162 , n1324 );
nand ( n2163 , n2162 , n1452 );
nand ( n2164 , n2161 , n2163 );
and ( n2165 , n1068 , n1196 );
not ( n2166 , n1068 );
not ( n2167 , n1196 );
and ( n2168 , n2166 , n2167 );
nor ( n2169 , n2165 , n2168 );
or ( n2170 , n2164 , n2169 );
not ( n2171 , n1324 );
not ( n2172 , n2159 );
or ( n2173 , n2171 , n2172 );
nand ( n2174 , n2173 , n2163 );
nand ( n2175 , n2174 , n2169 );
nand ( n2176 , n2170 , n2175 );
nand ( n2177 , n2157 , n2176 );
nor ( n2178 , n2136 , n2177 );
nand ( n2179 , n2109 , n2178 );
and ( n2180 , n1094 , n1222 );
not ( n2181 , n1094 );
not ( n2182 , n1222 );
and ( n2183 , n2181 , n2182 );
nor ( n2184 , n2180 , n2183 );
not ( n2185 , n1350 );
not ( n2186 , n2185 );
not ( n2187 , n1478 );
or ( n2188 , n2186 , n2187 );
not ( n2189 , n1478 );
nand ( n2190 , n2189 , n1350 );
nand ( n2191 , n2188 , n2190 );
or ( n2192 , n2184 , n2191 );
nand ( n2193 , n2185 , n1478 );
not ( n2194 , n2193 );
not ( n2195 , n2190 );
or ( n2196 , n2194 , n2195 );
and ( n2197 , n1094 , n1222 );
not ( n2198 , n1094 );
and ( n2199 , n2198 , n2182 );
nor ( n2200 , n2197 , n2199 );
nand ( n2201 , n2196 , n2200 );
nand ( n2202 , n2192 , n2201 );
and ( n2203 , n1095 , n1223 );
not ( n2204 , n1095 );
not ( n2205 , n1223 );
and ( n2206 , n2204 , n2205 );
nor ( n2207 , n2203 , n2206 );
not ( n2208 , n1479 );
and ( n2209 , n2208 , n1351 );
not ( n2210 , n1351 );
and ( n2211 , n2210 , n1479 );
nor ( n2212 , n2209 , n2211 );
and ( n2213 , n2207 , n2212 );
not ( n2214 , n2207 );
not ( n2215 , n1351 );
not ( n2216 , n2208 );
or ( n2217 , n2215 , n2216 );
nand ( n2218 , n2210 , n1479 );
nand ( n2219 , n2217 , n2218 );
and ( n2220 , n2214 , n2219 );
nor ( n2221 , n2213 , n2220 );
nand ( n2222 , n2202 , n2221 );
and ( n2223 , n1092 , n1220 );
not ( n2224 , n1092 );
not ( n2225 , n1220 );
and ( n2226 , n2224 , n2225 );
nor ( n2227 , n2223 , n2226 );
not ( n2228 , n1348 );
and ( n2229 , n2228 , n1476 );
not ( n2230 , n1476 );
and ( n2231 , n2230 , n1348 );
nor ( n2232 , n2229 , n2231 );
and ( n2233 , n2227 , n2232 );
not ( n2234 , n2227 );
not ( n2235 , n2228 );
not ( n2236 , n1476 );
or ( n2237 , n2235 , n2236 );
nand ( n2238 , n2230 , n1348 );
nand ( n2239 , n2237 , n2238 );
and ( n2240 , n2234 , n2239 );
nor ( n2241 , n2233 , n2240 );
and ( n2242 , n1349 , n1477 );
not ( n2243 , n1349 );
not ( n2244 , n1477 );
and ( n2245 , n2243 , n2244 );
nor ( n2246 , n2242 , n2245 );
xnor ( n2247 , n1221 , n1093 );
and ( n2248 , n2246 , n2247 );
not ( n2249 , n2246 );
xor ( n2250 , n1093 , n1221 );
and ( n2251 , n2249 , n2250 );
nor ( n2252 , n2248 , n2251 );
nand ( n2253 , n2241 , n2252 );
nor ( n2254 , n2222 , n2253 );
and ( n2255 , n1227 , n1355 );
not ( n2256 , n1227 );
not ( n2257 , n1355 );
and ( n2258 , n2256 , n2257 );
nor ( n2259 , n2255 , n2258 );
and ( n2260 , n1099 , n1483 );
not ( n2261 , n1099 );
not ( n2262 , n1483 );
and ( n2263 , n2261 , n2262 );
nor ( n2264 , n2260 , n2263 );
nand ( n2265 , n2259 , n2264 );
not ( n2266 , n2265 );
not ( n2267 , n2264 );
and ( n2268 , n1227 , n1355 );
not ( n2269 , n1227 );
and ( n2270 , n2269 , n2257 );
nor ( n2271 , n2268 , n2270 );
not ( n2272 , n2271 );
nand ( n2273 , n2267 , n2272 );
not ( n2274 , n2273 );
or ( n2275 , n2266 , n2274 );
not ( n2276 , n1354 );
not ( n2277 , n1482 );
not ( n2278 , n2277 );
or ( n2279 , n2276 , n2278 );
not ( n2280 , n1354 );
nand ( n2281 , n2280 , n1482 );
nand ( n2282 , n2279 , n2281 );
and ( n2283 , n1098 , n1226 );
not ( n2284 , n1098 );
not ( n2285 , n1226 );
and ( n2286 , n2284 , n2285 );
nor ( n2287 , n2283 , n2286 );
or ( n2288 , n2282 , n2287 );
not ( n2289 , n1354 );
not ( n2290 , n2277 );
or ( n2291 , n2289 , n2290 );
nand ( n2292 , n2291 , n2281 );
nand ( n2293 , n2292 , n2287 );
nand ( n2294 , n2288 , n2293 );
nand ( n2295 , n2275 , n2294 );
xor ( n2296 , n1481 , n1353 );
and ( n2297 , n1097 , n1225 );
not ( n2298 , n1097 );
not ( n2299 , n1225 );
and ( n2300 , n2298 , n2299 );
nor ( n2301 , n2297 , n2300 );
nand ( n2302 , n2296 , n2301 );
not ( n2303 , n2302 );
xnor ( n2304 , n1353 , n1481 );
not ( n2305 , n2299 );
not ( n2306 , n1097 );
and ( n2307 , n2305 , n2306 );
not ( n2308 , n1225 );
and ( n2309 , n2308 , n1097 );
nor ( n2310 , n2307 , n2309 );
nand ( n2311 , n2304 , n2310 );
not ( n2312 , n2311 );
or ( n2313 , n2303 , n2312 );
xor ( n2314 , n1096 , n1224 );
xor ( n2315 , n1352 , n1480 );
or ( n2316 , n2314 , n2315 );
xor ( n2317 , n1352 , n1480 );
xor ( n2318 , n1096 , n1224 );
nand ( n2319 , n2317 , n2318 );
nand ( n2320 , n2316 , n2319 );
nand ( n2321 , n2313 , n2320 );
nor ( n2322 , n2295 , n2321 );
nand ( n2323 , n2254 , n2322 );
nor ( n2324 , n2179 , n2323 );
and ( n2325 , n1344 , n1472 );
not ( n2326 , n1344 );
not ( n2327 , n1472 );
and ( n2328 , n2326 , n2327 );
nor ( n2329 , n2325 , n2328 );
not ( n2330 , n2329 );
and ( n2331 , n1088 , n1216 );
not ( n2332 , n1088 );
not ( n2333 , n1216 );
and ( n2334 , n2332 , n2333 );
nor ( n2335 , n2331 , n2334 );
not ( n2336 , n2335 );
or ( n2337 , n2330 , n2336 );
and ( n2338 , n1088 , n1216 );
not ( n2339 , n1088 );
and ( n2340 , n2339 , n2333 );
nor ( n2341 , n2338 , n2340 );
or ( n2342 , n2341 , n2329 );
nand ( n2343 , n2337 , n2342 );
not ( n2344 , n1089 );
and ( n2345 , n1217 , n2344 );
not ( n2346 , n1217 );
and ( n2347 , n2346 , n1089 );
nor ( n2348 , n2345 , n2347 );
and ( n2349 , n1345 , n1473 );
not ( n2350 , n1345 );
not ( n2351 , n1473 );
and ( n2352 , n2350 , n2351 );
nor ( n2353 , n2349 , n2352 );
and ( n2354 , n2348 , n2353 );
not ( n2355 , n2348 );
not ( n2356 , n2353 );
and ( n2357 , n2355 , n2356 );
nor ( n2358 , n2354 , n2357 );
nand ( n2359 , n2343 , n2358 );
not ( n2360 , n1347 );
and ( n2361 , n1475 , n2360 );
not ( n2362 , n1475 );
and ( n2363 , n2362 , n1347 );
nor ( n2364 , n2361 , n2363 );
and ( n2365 , n1091 , n1219 );
not ( n2366 , n1091 );
not ( n2367 , n1219 );
and ( n2368 , n2366 , n2367 );
nor ( n2369 , n2365 , n2368 );
and ( n2370 , n2364 , n2369 );
not ( n2371 , n2364 );
not ( n2372 , n2369 );
and ( n2373 , n2371 , n2372 );
nor ( n2374 , n2370 , n2373 );
and ( n2375 , n1218 , n1346 );
not ( n2376 , n1218 );
not ( n2377 , n1346 );
and ( n2378 , n2376 , n2377 );
nor ( n2379 , n2375 , n2378 );
xor ( n2380 , n1090 , n1474 );
not ( n2381 , n2380 );
and ( n2382 , n2379 , n2381 );
not ( n2383 , n2379 );
and ( n2384 , n2383 , n2380 );
nor ( n2385 , n2382 , n2384 );
nand ( n2386 , n2374 , n2385 );
nor ( n2387 , n2359 , n2386 );
and ( n2388 , n1087 , n1215 );
not ( n2389 , n1087 );
not ( n2390 , n1215 );
and ( n2391 , n2389 , n2390 );
nor ( n2392 , n2388 , n2391 );
not ( n2393 , n2392 );
xor ( n2394 , n1343 , n1471 );
not ( n2395 , n2394 );
or ( n2396 , n2393 , n2395 );
or ( n2397 , n2394 , n2392 );
nand ( n2398 , n2396 , n2397 );
xor ( n2399 , n1342 , n1470 );
xnor ( n2400 , n1086 , n1214 );
and ( n2401 , n2399 , n2400 );
not ( n2402 , n2399 );
xor ( n2403 , n1086 , n1214 );
and ( n2404 , n2402 , n2403 );
nor ( n2405 , n2401 , n2404 );
nand ( n2406 , n2398 , n2405 );
xor ( n2407 , n1212 , n1340 );
not ( n2408 , n1084 );
nand ( n2409 , n2408 , n1468 );
not ( n2410 , n1468 );
nand ( n2411 , n2410 , n1084 );
nand ( n2412 , n2409 , n2411 );
or ( n2413 , n2407 , n2412 );
not ( n2414 , n2411 );
not ( n2415 , n2409 );
or ( n2416 , n2414 , n2415 );
xor ( n2417 , n1212 , n1340 );
nand ( n2418 , n2416 , n2417 );
nand ( n2419 , n2413 , n2418 );
not ( n2420 , n1085 );
not ( n2421 , n1469 );
not ( n2422 , n2421 );
or ( n2423 , n2420 , n2422 );
not ( n2424 , n1085 );
nand ( n2425 , n2424 , n1469 );
nand ( n2426 , n2423 , n2425 );
not ( n2427 , n1213 );
or ( n2428 , n2427 , n1341 );
not ( n2429 , n1341 );
or ( n2430 , n2429 , n1213 );
nand ( n2431 , n2428 , n2430 );
or ( n2432 , n2426 , n2431 );
nand ( n2433 , n2421 , n1085 );
not ( n2434 , n2433 );
not ( n2435 , n2425 );
or ( n2436 , n2434 , n2435 );
xor ( n2437 , n1341 , n1213 );
nand ( n2438 , n2436 , n2437 );
nand ( n2439 , n2432 , n2438 );
nand ( n2440 , n2419 , n2439 );
nor ( n2441 , n2406 , n2440 );
nand ( n2442 , n2387 , n2441 );
xor ( n2443 , n1207 , n1079 );
and ( n2444 , n1335 , n1463 );
not ( n2445 , n1335 );
not ( n2446 , n1463 );
and ( n2447 , n2445 , n2446 );
nor ( n2448 , n2444 , n2447 );
nand ( n2449 , n2443 , n2448 );
not ( n2450 , n2449 );
not ( n2451 , n2448 );
xnor ( n2452 , n1079 , n1207 );
nand ( n2453 , n2451 , n2452 );
not ( n2454 , n2453 );
or ( n2455 , n2450 , n2454 );
not ( n2456 , n1078 );
not ( n2457 , n1462 );
not ( n2458 , n2457 );
or ( n2459 , n2456 , n2458 );
not ( n2460 , n1078 );
nand ( n2461 , n2460 , n1462 );
nand ( n2462 , n2459 , n2461 );
and ( n2463 , n1206 , n1334 );
not ( n2464 , n1206 );
not ( n2465 , n1334 );
and ( n2466 , n2464 , n2465 );
nor ( n2467 , n2463 , n2466 );
or ( n2468 , n2462 , n2467 );
not ( n2469 , n1078 );
not ( n2470 , n2457 );
or ( n2471 , n2469 , n2470 );
nand ( n2472 , n2471 , n2461 );
nand ( n2473 , n2472 , n2467 );
nand ( n2474 , n2468 , n2473 );
nand ( n2475 , n2455 , n2474 );
and ( n2476 , n1205 , n1333 );
not ( n2477 , n1205 );
not ( n2478 , n1333 );
and ( n2479 , n2477 , n2478 );
nor ( n2480 , n2476 , n2479 );
and ( n2481 , n1077 , n1461 );
not ( n2482 , n1077 );
not ( n2483 , n1461 );
and ( n2484 , n2482 , n2483 );
nor ( n2485 , n2481 , n2484 );
nand ( n2486 , n2480 , n2485 );
not ( n2487 , n2486 );
xnor ( n2488 , n1461 , n1077 );
and ( n2489 , n1333 , n1205 );
not ( n2490 , n1333 );
not ( n2491 , n1205 );
and ( n2492 , n2490 , n2491 );
nor ( n2493 , n2489 , n2492 );
not ( n2494 , n2493 );
nand ( n2495 , n2488 , n2494 );
not ( n2496 , n2495 );
or ( n2497 , n2487 , n2496 );
and ( n2498 , n1204 , n1332 );
not ( n2499 , n1204 );
not ( n2500 , n1332 );
and ( n2501 , n2499 , n2500 );
nor ( n2502 , n2498 , n2501 );
xnor ( n2503 , n1076 , n1460 );
and ( n2504 , n2502 , n2503 );
not ( n2505 , n2502 );
xor ( n2506 , n1076 , n1460 );
and ( n2507 , n2505 , n2506 );
nor ( n2508 , n2504 , n2507 );
nand ( n2509 , n2497 , n2508 );
nor ( n2510 , n2475 , n2509 );
xor ( n2511 , n1466 , n1338 );
and ( n2512 , n1082 , n1210 );
not ( n2513 , n1082 );
not ( n2514 , n1210 );
and ( n2515 , n2513 , n2514 );
nor ( n2516 , n2512 , n2515 );
or ( n2517 , n2511 , n2516 );
xor ( n2518 , n1338 , n1466 );
nand ( n2519 , n2518 , n2516 );
nand ( n2520 , n2517 , n2519 );
not ( n2521 , n1083 );
and ( n2522 , n1211 , n2521 );
not ( n2523 , n1211 );
and ( n2524 , n2523 , n1083 );
nor ( n2525 , n2522 , n2524 );
and ( n2526 , n1339 , n1467 );
not ( n2527 , n1339 );
not ( n2528 , n1467 );
and ( n2529 , n2527 , n2528 );
nor ( n2530 , n2526 , n2529 );
and ( n2531 , n2525 , n2530 );
not ( n2532 , n2525 );
and ( n2533 , n1339 , n1467 );
not ( n2534 , n1339 );
and ( n2535 , n2534 , n2528 );
nor ( n2536 , n2533 , n2535 );
not ( n2537 , n2536 );
and ( n2538 , n2532 , n2537 );
nor ( n2539 , n2531 , n2538 );
nand ( n2540 , n2520 , n2539 );
and ( n2541 , n1336 , n1464 );
not ( n2542 , n1336 );
not ( n2543 , n1464 );
and ( n2544 , n2542 , n2543 );
nor ( n2545 , n2541 , n2544 );
xnor ( n2546 , n1208 , n1080 );
and ( n2547 , n2545 , n2546 );
not ( n2548 , n2545 );
and ( n2549 , n1080 , n1208 );
not ( n2550 , n1080 );
not ( n2551 , n1208 );
and ( n2552 , n2550 , n2551 );
nor ( n2553 , n2549 , n2552 );
and ( n2554 , n2548 , n2553 );
nor ( n2555 , n2547 , n2554 );
and ( n2556 , n1081 , n1465 );
not ( n2557 , n1081 );
not ( n2558 , n1465 );
and ( n2559 , n2557 , n2558 );
nor ( n2560 , n2556 , n2559 );
xnor ( n2561 , n1337 , n1209 );
and ( n2562 , n2560 , n2561 );
not ( n2563 , n2560 );
and ( n2564 , n1209 , n1337 );
not ( n2565 , n1209 );
not ( n2566 , n1337 );
and ( n2567 , n2565 , n2566 );
nor ( n2568 , n2564 , n2567 );
and ( n2569 , n2563 , n2568 );
nor ( n2570 , n2562 , n2569 );
nand ( n2571 , n2555 , n2570 );
nor ( n2572 , n2540 , n2571 );
nand ( n2573 , n2510 , n2572 );
nor ( n2574 , n2442 , n2573 );
nand ( n2575 , n2324 , n2574 );
nor ( n2576 , n2046 , n2575 );
xor ( n2577 , n1103 , n1487 );
not ( n2578 , n2577 );
and ( n2579 , n1231 , n1359 );
not ( n2580 , n1231 );
not ( n2581 , n1359 );
and ( n2582 , n2580 , n2581 );
nor ( n2583 , n2579 , n2582 );
not ( n2584 , n2583 );
or ( n2585 , n2578 , n2584 );
or ( n2586 , n2583 , n2577 );
nand ( n2587 , n2585 , n2586 );
and ( n2588 , n1358 , n1486 );
not ( n2589 , n1358 );
not ( n2590 , n1486 );
and ( n2591 , n2589 , n2590 );
nor ( n2592 , n2588 , n2591 );
not ( n2593 , n2592 );
and ( n2594 , n1102 , n1230 );
not ( n2595 , n1102 );
not ( n2596 , n1230 );
and ( n2597 , n2595 , n2596 );
nor ( n2598 , n2594 , n2597 );
not ( n2599 , n2598 );
or ( n2600 , n2593 , n2599 );
or ( n2601 , n2592 , n2598 );
nand ( n2602 , n2600 , n2601 );
nand ( n2603 , n2587 , n2602 );
xor ( n2604 , n1100 , n1484 );
not ( n2605 , n2604 );
and ( n2606 , n1228 , n1356 );
not ( n2607 , n1228 );
not ( n2608 , n1356 );
and ( n2609 , n2607 , n2608 );
nor ( n2610 , n2606 , n2609 );
not ( n2611 , n2610 );
or ( n2612 , n2605 , n2611 );
or ( n2613 , n2604 , n2610 );
nand ( n2614 , n2612 , n2613 );
and ( n2615 , n1101 , n1229 );
not ( n2616 , n1101 );
not ( n2617 , n1229 );
and ( n2618 , n2616 , n2617 );
nor ( n2619 , n2615 , n2618 );
xor ( n2620 , n1357 , n1485 );
not ( n2621 , n2620 );
and ( n2622 , n2619 , n2621 );
not ( n2623 , n2619 );
and ( n2624 , n2623 , n2620 );
nor ( n2625 , n2622 , n2624 );
nand ( n2626 , n2614 , n2625 );
nor ( n2627 , n2603 , n2626 );
and ( n2628 , n1363 , n1491 );
not ( n2629 , n1363 );
not ( n2630 , n1491 );
and ( n2631 , n2629 , n2630 );
nor ( n2632 , n2628 , n2631 );
not ( n2633 , n2632 );
and ( n2634 , n1107 , n1235 );
not ( n2635 , n1107 );
not ( n2636 , n1235 );
and ( n2637 , n2635 , n2636 );
nor ( n2638 , n2634 , n2637 );
not ( n2639 , n2638 );
or ( n2640 , n2633 , n2639 );
or ( n2641 , n2638 , n2632 );
nand ( n2642 , n2640 , n2641 );
xor ( n2643 , n1106 , n1490 );
not ( n2644 , n2643 );
and ( n2645 , n1234 , n1362 );
not ( n2646 , n1234 );
not ( n2647 , n1362 );
and ( n2648 , n2646 , n2647 );
nor ( n2649 , n2645 , n2648 );
not ( n2650 , n2649 );
or ( n2651 , n2644 , n2650 );
or ( n2652 , n2649 , n2643 );
nand ( n2653 , n2651 , n2652 );
nand ( n2654 , n2642 , n2653 );
and ( n2655 , n1104 , n1488 );
not ( n2656 , n1104 );
not ( n2657 , n1488 );
and ( n2658 , n2656 , n2657 );
nor ( n2659 , n2655 , n2658 );
not ( n2660 , n2659 );
and ( n2661 , n1232 , n1360 );
not ( n2662 , n1232 );
not ( n2663 , n1360 );
and ( n2664 , n2662 , n2663 );
nor ( n2665 , n2661 , n2664 );
not ( n2666 , n2665 );
or ( n2667 , n2660 , n2666 );
or ( n2668 , n2659 , n2665 );
nand ( n2669 , n2667 , n2668 );
not ( n2670 , n1233 );
and ( n2671 , n1361 , n2670 );
not ( n2672 , n1361 );
and ( n2673 , n2672 , n1233 );
nor ( n2674 , n2671 , n2673 );
and ( n2675 , n1105 , n1489 );
not ( n2676 , n1105 );
not ( n2677 , n1489 );
and ( n2678 , n2676 , n2677 );
nor ( n2679 , n2675 , n2678 );
and ( n2680 , n2674 , n2679 );
not ( n2681 , n2674 );
not ( n2682 , n2679 );
and ( n2683 , n2681 , n2682 );
nor ( n2684 , n2680 , n2683 );
nand ( n2685 , n2669 , n2684 );
nor ( n2686 , n2654 , n2685 );
nand ( n2687 , n2627 , n2686 );
xor ( n2688 , n1108 , n1492 );
and ( n2689 , n1236 , n1364 );
not ( n2690 , n1236 );
not ( n2691 , n1364 );
and ( n2692 , n2690 , n2691 );
nor ( n2693 , n2689 , n2692 );
not ( n2694 , n2693 );
and ( n2695 , n2688 , n2694 );
not ( n2696 , n2688 );
and ( n2697 , n2696 , n2693 );
nor ( n2698 , n2695 , n2697 );
xor ( n2699 , n1365 , n1493 );
and ( n2700 , n1109 , n1237 );
not ( n2701 , n1109 );
not ( n2702 , n1237 );
and ( n2703 , n2701 , n2702 );
nor ( n2704 , n2700 , n2703 );
not ( n2705 , n2704 );
and ( n2706 , n2699 , n2705 );
not ( n2707 , n2699 );
and ( n2708 , n2707 , n2704 );
nor ( n2709 , n2706 , n2708 );
nand ( n2710 , n2698 , n2709 );
and ( n2711 , n1111 , n1239 );
not ( n2712 , n1111 );
not ( n2713 , n1239 );
and ( n2714 , n2712 , n2713 );
nor ( n2715 , n2711 , n2714 );
xor ( n2716 , n1367 , n1495 );
not ( n2717 , n2716 );
and ( n2718 , n2715 , n2717 );
not ( n2719 , n2715 );
and ( n2720 , n2719 , n2716 );
nor ( n2721 , n2718 , n2720 );
and ( n2722 , n1110 , n1238 );
not ( n2723 , n1110 );
not ( n2724 , n1238 );
and ( n2725 , n2723 , n2724 );
nor ( n2726 , n2722 , n2725 );
xor ( n2727 , n1366 , n1494 );
not ( n2728 , n2727 );
and ( n2729 , n2726 , n2728 );
not ( n2730 , n2726 );
and ( n2731 , n2730 , n2727 );
nor ( n2732 , n2729 , n2731 );
nand ( n2733 , n2721 , n2732 );
nor ( n2734 , n2710 , n2733 );
and ( n2735 , n1112 , n1240 );
not ( n2736 , n1112 );
not ( n2737 , n1240 );
and ( n2738 , n2736 , n2737 );
nor ( n2739 , n2735 , n2738 );
xor ( n2740 , n1368 , n1496 );
nand ( n2741 , n2739 , n2740 );
not ( n2742 , n2741 );
not ( n2743 , n2739 );
not ( n2744 , n2740 );
nand ( n2745 , n2743 , n2744 );
not ( n2746 , n2745 );
or ( n2747 , n2742 , n2746 );
not ( n2748 , n1113 );
and ( n2749 , n1241 , n2748 );
not ( n2750 , n1241 );
and ( n2751 , n2750 , n1113 );
nor ( n2752 , n2749 , n2751 );
and ( n2753 , n1369 , n1497 );
not ( n2754 , n1369 );
not ( n2755 , n1497 );
and ( n2756 , n2754 , n2755 );
nor ( n2757 , n2753 , n2756 );
and ( n2758 , n2752 , n2757 );
not ( n2759 , n2752 );
not ( n2760 , n2757 );
and ( n2761 , n2759 , n2760 );
nor ( n2762 , n2758 , n2761 );
nand ( n2763 , n2747 , n2762 );
and ( n2764 , n1114 , n1242 );
not ( n2765 , n1114 );
not ( n2766 , n1242 );
and ( n2767 , n2765 , n2766 );
nor ( n2768 , n2764 , n2767 );
xor ( n2769 , n1370 , n1498 );
not ( n2770 , n2769 );
and ( n2771 , n2768 , n2770 );
not ( n2772 , n2768 );
and ( n2773 , n2772 , n2769 );
nor ( n2774 , n2771 , n2773 );
and ( n2775 , n1371 , n1499 );
not ( n2776 , n1371 );
not ( n2777 , n1499 );
and ( n2778 , n2776 , n2777 );
nor ( n2779 , n2775 , n2778 );
and ( n2780 , n1115 , n1243 );
not ( n2781 , n1115 );
not ( n2782 , n1243 );
and ( n2783 , n2781 , n2782 );
nor ( n2784 , n2780 , n2783 );
not ( n2785 , n2784 );
and ( n2786 , n2779 , n2785 );
not ( n2787 , n2779 );
and ( n2788 , n2787 , n2784 );
nor ( n2789 , n2786 , n2788 );
nand ( n2790 , n2774 , n2789 );
nor ( n2791 , n2763 , n2790 );
nand ( n2792 , n2734 , n2791 );
nor ( n2793 , n2687 , n2792 );
and ( n2794 , n1379 , n1507 );
not ( n2795 , n1379 );
not ( n2796 , n1507 );
and ( n2797 , n2795 , n2796 );
nor ( n2798 , n2794 , n2797 );
not ( n2799 , n2798 );
and ( n2800 , n1123 , n1251 );
not ( n2801 , n1123 );
not ( n2802 , n1251 );
and ( n2803 , n2801 , n2802 );
nor ( n2804 , n2800 , n2803 );
not ( n2805 , n2804 );
or ( n2806 , n2799 , n2805 );
or ( n2807 , n2798 , n2804 );
nand ( n2808 , n2806 , n2807 );
and ( n2809 , n1378 , n1506 );
not ( n2810 , n1378 );
not ( n2811 , n1506 );
and ( n2812 , n2810 , n2811 );
nor ( n2813 , n2809 , n2812 );
not ( n2814 , n2813 );
and ( n2815 , n1122 , n1250 );
not ( n2816 , n1122 );
not ( n2817 , n1250 );
and ( n2818 , n2816 , n2817 );
nor ( n2819 , n2815 , n2818 );
not ( n2820 , n2819 );
or ( n2821 , n2814 , n2820 );
or ( n2822 , n2813 , n2819 );
nand ( n2823 , n2821 , n2822 );
nand ( n2824 , n2808 , n2823 );
xor ( n2825 , n1376 , n1504 );
not ( n2826 , n2825 );
and ( n2827 , n1120 , n1248 );
not ( n2828 , n1120 );
not ( n2829 , n1248 );
and ( n2830 , n2828 , n2829 );
nor ( n2831 , n2827 , n2830 );
not ( n2832 , n2831 );
or ( n2833 , n2826 , n2832 );
or ( n2834 , n2831 , n2825 );
nand ( n2835 , n2833 , n2834 );
and ( n2836 , n1121 , n1249 );
not ( n2837 , n1121 );
not ( n2838 , n1249 );
and ( n2839 , n2837 , n2838 );
nor ( n2840 , n2836 , n2839 );
xor ( n2841 , n1377 , n1505 );
not ( n2842 , n2841 );
and ( n2843 , n2840 , n2842 );
not ( n2844 , n2840 );
and ( n2845 , n2844 , n2841 );
nor ( n2846 , n2843 , n2845 );
nand ( n2847 , n2835 , n2846 );
nor ( n2848 , n2824 , n2847 );
and ( n2849 , n1117 , n1245 );
not ( n2850 , n1117 );
not ( n2851 , n1245 );
and ( n2852 , n2850 , n2851 );
nor ( n2853 , n2849 , n2852 );
and ( n2854 , n1373 , n1501 );
not ( n2855 , n1373 );
not ( n2856 , n1501 );
and ( n2857 , n2855 , n2856 );
nor ( n2858 , n2854 , n2857 );
not ( n2859 , n2858 );
and ( n2860 , n2853 , n2859 );
not ( n2861 , n2853 );
and ( n2862 , n2861 , n2858 );
nor ( n2863 , n2860 , n2862 );
xor ( n2864 , n1116 , n1500 );
and ( n2865 , n1244 , n1372 );
not ( n2866 , n1244 );
not ( n2867 , n1372 );
and ( n2868 , n2866 , n2867 );
nor ( n2869 , n2865 , n2868 );
not ( n2870 , n2869 );
and ( n2871 , n2864 , n2870 );
not ( n2872 , n2864 );
and ( n2873 , n2872 , n2869 );
nor ( n2874 , n2871 , n2873 );
nand ( n2875 , n2863 , n2874 );
and ( n2876 , n1118 , n1246 );
not ( n2877 , n1118 );
not ( n2878 , n1246 );
and ( n2879 , n2877 , n2878 );
nor ( n2880 , n2876 , n2879 );
and ( n2881 , n1374 , n1502 );
not ( n2882 , n1374 );
not ( n2883 , n1502 );
and ( n2884 , n2882 , n2883 );
nor ( n2885 , n2881 , n2884 );
nand ( n2886 , n2880 , n2885 );
not ( n2887 , n2886 );
nor ( n2888 , n2885 , n2880 );
or ( n2889 , n2887 , n2888 );
and ( n2890 , n1119 , n1247 );
not ( n2891 , n1119 );
not ( n2892 , n1247 );
and ( n2893 , n2891 , n2892 );
nor ( n2894 , n2890 , n2893 );
xor ( n2895 , n1375 , n1503 );
or ( n2896 , n2894 , n2895 );
and ( n2897 , n1119 , n1247 );
not ( n2898 , n1119 );
and ( n2899 , n2898 , n2892 );
nor ( n2900 , n2897 , n2899 );
nand ( n2901 , n2900 , n2895 );
nand ( n2902 , n2896 , n2901 );
nand ( n2903 , n2889 , n2902 );
nor ( n2904 , n2875 , n2903 );
nand ( n2905 , n2848 , n2904 );
and ( n2906 , n1387 , n1515 );
not ( n2907 , n1387 );
not ( n2908 , n1515 );
and ( n2909 , n2907 , n2908 );
nor ( n2910 , n2906 , n2909 );
not ( n2911 , n2910 );
and ( n2912 , n1131 , n1259 );
not ( n2913 , n1131 );
not ( n2914 , n1259 );
and ( n2915 , n2913 , n2914 );
nor ( n2916 , n2912 , n2915 );
not ( n2917 , n2916 );
or ( n2918 , n2911 , n2917 );
or ( n2919 , n2916 , n2910 );
nand ( n2920 , n2918 , n2919 );
and ( n2921 , n1130 , n1258 );
not ( n2922 , n1130 );
not ( n2923 , n1258 );
and ( n2924 , n2922 , n2923 );
nor ( n2925 , n2921 , n2924 );
not ( n2926 , n2925 );
xor ( n2927 , n1386 , n1514 );
not ( n2928 , n2927 );
or ( n2929 , n2926 , n2928 );
or ( n2930 , n2927 , n2925 );
nand ( n2931 , n2929 , n2930 );
nand ( n2932 , n2920 , n2931 );
xor ( n2933 , n1385 , n1513 );
and ( n2934 , n1129 , n1257 );
not ( n2935 , n1129 );
not ( n2936 , n1257 );
and ( n2937 , n2935 , n2936 );
nor ( n2938 , n2934 , n2937 );
not ( n2939 , n2938 );
and ( n2940 , n2933 , n2939 );
not ( n2941 , n2933 );
and ( n2942 , n2941 , n2938 );
nor ( n2943 , n2940 , n2942 );
xor ( n2944 , n1384 , n1512 );
and ( n2945 , n1128 , n1256 );
not ( n2946 , n1128 );
not ( n2947 , n1256 );
and ( n2948 , n2946 , n2947 );
nor ( n2949 , n2945 , n2948 );
not ( n2950 , n2949 );
and ( n2951 , n2944 , n2950 );
not ( n2952 , n2944 );
and ( n2953 , n2952 , n2949 );
nor ( n2954 , n2951 , n2953 );
nand ( n2955 , n2943 , n2954 );
nor ( n2956 , n2932 , n2955 );
and ( n2957 , n1509 , n1125 );
not ( n2958 , n1509 );
not ( n2959 , n1125 );
and ( n2960 , n2958 , n2959 );
nor ( n2961 , n2957 , n2960 );
and ( n2962 , n1253 , n1381 );
not ( n2963 , n1253 );
not ( n2964 , n1381 );
and ( n2965 , n2963 , n2964 );
nor ( n2966 , n2962 , n2965 );
nand ( n2967 , n2961 , n2966 );
not ( n2968 , n2967 );
not ( n2969 , n2966 );
and ( n2970 , n1509 , n1125 );
not ( n2971 , n1509 );
and ( n2972 , n2971 , n2959 );
nor ( n2973 , n2970 , n2972 );
not ( n2974 , n2973 );
nand ( n2975 , n2969 , n2974 );
not ( n2976 , n2975 );
or ( n2977 , n2968 , n2976 );
not ( n2978 , n1380 );
nand ( n2979 , n2978 , n1508 );
not ( n2980 , n1508 );
nand ( n2981 , n2980 , n1380 );
nand ( n2982 , n2979 , n2981 );
and ( n2983 , n1124 , n1252 );
not ( n2984 , n1124 );
not ( n2985 , n1252 );
and ( n2986 , n2984 , n2985 );
nor ( n2987 , n2983 , n2986 );
or ( n2988 , n2982 , n2987 );
nand ( n2989 , n2982 , n2987 );
nand ( n2990 , n2988 , n2989 );
nand ( n2991 , n2977 , n2990 );
and ( n2992 , n1255 , n1383 );
not ( n2993 , n1255 );
not ( n2994 , n1383 );
and ( n2995 , n2993 , n2994 );
nor ( n2996 , n2992 , n2995 );
xor ( n2997 , n1127 , n1511 );
not ( n2998 , n2997 );
and ( n2999 , n2996 , n2998 );
not ( n3000 , n2996 );
and ( n3001 , n3000 , n2997 );
nor ( n3002 , n2999 , n3001 );
and ( n3003 , n1126 , n1254 );
not ( n3004 , n1126 );
not ( n3005 , n1254 );
and ( n3006 , n3004 , n3005 );
nor ( n3007 , n3003 , n3006 );
xor ( n3008 , n1382 , n1510 );
not ( n3009 , n3008 );
and ( n3010 , n3007 , n3009 );
not ( n3011 , n3007 );
and ( n3012 , n3011 , n3008 );
nor ( n3013 , n3010 , n3012 );
nand ( n3014 , n3002 , n3013 );
nor ( n3015 , n2991 , n3014 );
nand ( n3016 , n2956 , n3015 );
nor ( n3017 , n2905 , n3016 );
nand ( n3018 , n2793 , n3017 );
not ( n3019 , n3018 );
not ( n3020 , n1139 );
and ( n3021 , n1267 , n3020 );
not ( n3022 , n1267 );
and ( n3023 , n3022 , n1139 );
nor ( n3024 , n3021 , n3023 );
and ( n3025 , n1395 , n1523 );
not ( n3026 , n1395 );
not ( n3027 , n1523 );
and ( n3028 , n3026 , n3027 );
nor ( n3029 , n3025 , n3028 );
and ( n3030 , n3024 , n3029 );
not ( n3031 , n3024 );
not ( n3032 , n3029 );
and ( n3033 , n3031 , n3032 );
nor ( n3034 , n3030 , n3033 );
and ( n3035 , n1138 , n1266 );
not ( n3036 , n1138 );
not ( n3037 , n1266 );
and ( n3038 , n3036 , n3037 );
nor ( n3039 , n3035 , n3038 );
and ( n3040 , n1394 , n1522 );
not ( n3041 , n1394 );
not ( n3042 , n1522 );
and ( n3043 , n3041 , n3042 );
nor ( n3044 , n3040 , n3043 );
not ( n3045 , n3044 );
and ( n3046 , n3039 , n3045 );
not ( n3047 , n3039 );
and ( n3048 , n3047 , n3044 );
nor ( n3049 , n3046 , n3048 );
nand ( n3050 , n3034 , n3049 );
and ( n3051 , n1136 , n1264 );
not ( n3052 , n1136 );
not ( n3053 , n1264 );
and ( n3054 , n3052 , n3053 );
nor ( n3055 , n3051 , n3054 );
xor ( n3056 , n1392 , n1520 );
nand ( n3057 , n3055 , n3056 );
not ( n3058 , n3057 );
and ( n3059 , n1136 , n1264 );
not ( n3060 , n1136 );
and ( n3061 , n3060 , n3053 );
or ( n3062 , n3059 , n3061 );
not ( n3063 , n3056 );
nand ( n3064 , n3062 , n3063 );
not ( n3065 , n3064 );
or ( n3066 , n3058 , n3065 );
not ( n3067 , n1265 );
and ( n3068 , n1393 , n3067 );
not ( n3069 , n1393 );
and ( n3070 , n3069 , n1265 );
nor ( n3071 , n3068 , n3070 );
and ( n3072 , n1137 , n1521 );
not ( n3073 , n1137 );
not ( n3074 , n1521 );
and ( n3075 , n3073 , n3074 );
nor ( n3076 , n3072 , n3075 );
and ( n3077 , n3071 , n3076 );
not ( n3078 , n3071 );
not ( n3079 , n3076 );
and ( n3080 , n3078 , n3079 );
nor ( n3081 , n3077 , n3080 );
nand ( n3082 , n3066 , n3081 );
nor ( n3083 , n3050 , n3082 );
and ( n3084 , n1263 , n1391 );
not ( n3085 , n1263 );
not ( n3086 , n1391 );
and ( n3087 , n3085 , n3086 );
nor ( n3088 , n3084 , n3087 );
not ( n3089 , n3088 );
xor ( n3090 , n1135 , n1519 );
not ( n3091 , n3090 );
or ( n3092 , n3089 , n3091 );
or ( n3093 , n3090 , n3088 );
nand ( n3094 , n3092 , n3093 );
and ( n3095 , n1390 , n1518 );
not ( n3096 , n1390 );
not ( n3097 , n1518 );
and ( n3098 , n3096 , n3097 );
nor ( n3099 , n3095 , n3098 );
not ( n3100 , n3099 );
and ( n3101 , n1134 , n1262 );
not ( n3102 , n1134 );
not ( n3103 , n1262 );
and ( n3104 , n3102 , n3103 );
nor ( n3105 , n3101 , n3104 );
not ( n3106 , n3105 );
or ( n3107 , n3100 , n3106 );
and ( n3108 , n1134 , n1262 );
not ( n3109 , n1134 );
and ( n3110 , n3109 , n3103 );
nor ( n3111 , n3108 , n3110 );
or ( n3112 , n3111 , n3099 );
nand ( n3113 , n3107 , n3112 );
nand ( n3114 , n3094 , n3113 );
xor ( n3115 , n1133 , n1517 );
and ( n3116 , n1261 , n1389 );
not ( n3117 , n1261 );
not ( n3118 , n1389 );
and ( n3119 , n3117 , n3118 );
nor ( n3120 , n3116 , n3119 );
not ( n3121 , n3120 );
and ( n3122 , n3115 , n3121 );
not ( n3123 , n3115 );
and ( n3124 , n3123 , n3120 );
nor ( n3125 , n3122 , n3124 );
xor ( n3126 , n1132 , n1516 );
and ( n3127 , n1260 , n1388 );
not ( n3128 , n1260 );
not ( n3129 , n1388 );
and ( n3130 , n3128 , n3129 );
nor ( n3131 , n3127 , n3130 );
not ( n3132 , n3131 );
and ( n3133 , n3126 , n3132 );
not ( n3134 , n3126 );
and ( n3135 , n3134 , n3131 );
nor ( n3136 , n3133 , n3135 );
nand ( n3137 , n3125 , n3136 );
nor ( n3138 , n3114 , n3137 );
nand ( n3139 , n3083 , n3138 );
not ( n3140 , n1402 );
nand ( n3141 , n3140 , n1530 );
not ( n3142 , n1530 );
nand ( n3143 , n3142 , n1402 );
nand ( n3144 , n3141 , n3143 );
and ( n3145 , n1146 , n1274 );
not ( n3146 , n1146 );
not ( n3147 , n1274 );
and ( n3148 , n3146 , n3147 );
nor ( n3149 , n3145 , n3148 );
or ( n3150 , n3144 , n3149 );
not ( n3151 , n3143 );
not ( n3152 , n3141 );
or ( n3153 , n3151 , n3152 );
nand ( n3154 , n3153 , n3149 );
nand ( n3155 , n3150 , n3154 );
and ( n3156 , n1403 , n1531 );
not ( n3157 , n1403 );
not ( n3158 , n1531 );
and ( n3159 , n3157 , n3158 );
nor ( n3160 , n3156 , n3159 );
and ( n3161 , n1147 , n1275 );
not ( n3162 , n1147 );
not ( n3163 , n1275 );
and ( n3164 , n3162 , n3163 );
nor ( n3165 , n3161 , n3164 );
not ( n3166 , n3165 );
and ( n3167 , n3160 , n3166 );
not ( n3168 , n3160 );
and ( n3169 , n3168 , n3165 );
nor ( n3170 , n3167 , n3169 );
nand ( n3171 , n3155 , n3170 );
and ( n3172 , n1529 , n1401 );
not ( n3173 , n1529 );
not ( n3174 , n1401 );
and ( n3175 , n3173 , n3174 );
nor ( n3176 , n3172 , n3175 );
not ( n3177 , n3176 );
and ( n3178 , n1273 , n1145 );
not ( n3179 , n1273 );
not ( n3180 , n1145 );
and ( n3181 , n3179 , n3180 );
nor ( n3182 , n3178 , n3181 );
not ( n3183 , n3182 );
or ( n3184 , n3177 , n3183 );
and ( n3185 , n1145 , n1273 );
not ( n3186 , n1145 );
not ( n3187 , n1273 );
and ( n3188 , n3186 , n3187 );
nor ( n3189 , n3185 , n3188 );
and ( n3190 , n1401 , n1529 );
not ( n3191 , n1401 );
not ( n3192 , n1529 );
and ( n3193 , n3191 , n3192 );
nor ( n3194 , n3190 , n3193 );
or ( n3195 , n3189 , n3194 );
nand ( n3196 , n3184 , n3195 );
not ( n3197 , n1400 );
not ( n3198 , n1528 );
not ( n3199 , n3198 );
or ( n3200 , n3197 , n3199 );
not ( n3201 , n1400 );
nand ( n3202 , n3201 , n1528 );
nand ( n3203 , n3200 , n3202 );
and ( n3204 , n1144 , n1272 );
not ( n3205 , n1144 );
not ( n3206 , n1272 );
and ( n3207 , n3205 , n3206 );
nor ( n3208 , n3204 , n3207 );
or ( n3209 , n3203 , n3208 );
not ( n3210 , n3202 );
nand ( n3211 , n3198 , n1400 );
not ( n3212 , n3211 );
or ( n3213 , n3210 , n3212 );
nand ( n3214 , n3213 , n3208 );
nand ( n3215 , n3209 , n3214 );
nand ( n3216 , n3196 , n3215 );
nor ( n3217 , n3171 , n3216 );
and ( n3218 , n1143 , n1271 );
not ( n3219 , n1143 );
not ( n3220 , n1271 );
and ( n3221 , n3219 , n3220 );
nor ( n3222 , n3218 , n3221 );
not ( n3223 , n1399 );
not ( n3224 , n1527 );
not ( n3225 , n3224 );
or ( n3226 , n3223 , n3225 );
not ( n3227 , n1399 );
nand ( n3228 , n3227 , n1527 );
nand ( n3229 , n3226 , n3228 );
or ( n3230 , n3222 , n3229 );
not ( n3231 , n3228 );
nand ( n3232 , n3224 , n1399 );
not ( n3233 , n3232 );
or ( n3234 , n3231 , n3233 );
nand ( n3235 , n3234 , n3222 );
nand ( n3236 , n3230 , n3235 );
not ( n3237 , n1526 );
and ( n3238 , n1142 , n3237 );
not ( n3239 , n1142 );
and ( n3240 , n3239 , n1526 );
nor ( n3241 , n3238 , n3240 );
and ( n3242 , n1270 , n1398 );
not ( n3243 , n1270 );
not ( n3244 , n1398 );
and ( n3245 , n3243 , n3244 );
nor ( n3246 , n3242 , n3245 );
and ( n3247 , n3241 , n3246 );
not ( n3248 , n3241 );
not ( n3249 , n3246 );
and ( n3250 , n3248 , n3249 );
nor ( n3251 , n3247 , n3250 );
nand ( n3252 , n3236 , n3251 );
not ( n3253 , n1525 );
nand ( n3254 , n3253 , n1141 );
not ( n3255 , n1141 );
nand ( n3256 , n3255 , n1525 );
nand ( n3257 , n3254 , n3256 );
and ( n3258 , n1269 , n1397 );
not ( n3259 , n1269 );
not ( n3260 , n1397 );
and ( n3261 , n3259 , n3260 );
nor ( n3262 , n3258 , n3261 );
or ( n3263 , n3257 , n3262 );
nand ( n3264 , n3255 , n1525 );
not ( n3265 , n3264 );
not ( n3266 , n3254 );
or ( n3267 , n3265 , n3266 );
nand ( n3268 , n3267 , n3262 );
nand ( n3269 , n3263 , n3268 );
not ( n3270 , n1396 );
not ( n3271 , n3270 );
not ( n3272 , n1524 );
or ( n3273 , n3271 , n3272 );
not ( n3274 , n1524 );
nand ( n3275 , n3274 , n1396 );
nand ( n3276 , n3273 , n3275 );
and ( n3277 , n1140 , n1268 );
not ( n3278 , n1140 );
not ( n3279 , n1268 );
and ( n3280 , n3278 , n3279 );
nor ( n3281 , n3277 , n3280 );
or ( n3282 , n3276 , n3281 );
nand ( n3283 , n3274 , n1396 );
not ( n3284 , n3283 );
nand ( n3285 , n3270 , n1524 );
not ( n3286 , n3285 );
or ( n3287 , n3284 , n3286 );
nand ( n3288 , n3287 , n3281 );
nand ( n3289 , n3282 , n3288 );
nand ( n3290 , n3269 , n3289 );
nor ( n3291 , n3252 , n3290 );
nand ( n3292 , n3217 , n3291 );
nor ( n3293 , n3139 , n3292 );
and ( n3294 , n1155 , n1283 );
not ( n3295 , n1155 );
not ( n3296 , n1283 );
and ( n3297 , n3295 , n3296 );
nor ( n3298 , n3294 , n3297 );
not ( n3299 , n3298 );
xor ( n3300 , n1411 , n1539 );
not ( n3301 , n3300 );
or ( n3302 , n3299 , n3301 );
or ( n3303 , n3298 , n3300 );
nand ( n3304 , n3302 , n3303 );
and ( n3305 , n1282 , n1410 );
not ( n3306 , n1282 );
not ( n3307 , n1410 );
and ( n3308 , n3306 , n3307 );
nor ( n3309 , n3305 , n3308 );
not ( n3310 , n3309 );
xor ( n3311 , n1154 , n1538 );
not ( n3312 , n3311 );
or ( n3313 , n3310 , n3312 );
or ( n3314 , n3309 , n3311 );
nand ( n3315 , n3313 , n3314 );
nand ( n3316 , n3304 , n3315 );
not ( n3317 , n1153 );
not ( n3318 , n1537 );
not ( n3319 , n3318 );
or ( n3320 , n3317 , n3319 );
not ( n3321 , n1153 );
nand ( n3322 , n3321 , n1537 );
nand ( n3323 , n3320 , n3322 );
not ( n3324 , n3323 );
and ( n3325 , n1281 , n1409 );
not ( n3326 , n1281 );
not ( n3327 , n1409 );
and ( n3328 , n3326 , n3327 );
nor ( n3329 , n3325 , n3328 );
not ( n3330 , n3329 );
or ( n3331 , n3324 , n3330 );
and ( n3332 , n1281 , n1409 );
not ( n3333 , n1281 );
and ( n3334 , n3333 , n3327 );
nor ( n3335 , n3332 , n3334 );
not ( n3336 , n1153 );
not ( n3337 , n3318 );
or ( n3338 , n3336 , n3337 );
nand ( n3339 , n3338 , n3322 );
or ( n3340 , n3335 , n3339 );
nand ( n3341 , n3331 , n3340 );
not ( n3342 , n1536 );
and ( n3343 , n1152 , n3342 );
not ( n3344 , n1152 );
and ( n3345 , n3344 , n1536 );
nor ( n3346 , n3343 , n3345 );
and ( n3347 , n1280 , n1408 );
not ( n3348 , n1280 );
not ( n3349 , n1408 );
and ( n3350 , n3348 , n3349 );
nor ( n3351 , n3347 , n3350 );
and ( n3352 , n3346 , n3351 );
not ( n3353 , n3346 );
not ( n3354 , n3351 );
and ( n3355 , n3353 , n3354 );
nor ( n3356 , n3352 , n3355 );
nand ( n3357 , n3341 , n3356 );
nor ( n3358 , n3316 , n3357 );
xor ( n3359 , n1532 , n1404 );
and ( n3360 , n1148 , n1276 );
not ( n3361 , n1148 );
not ( n3362 , n1276 );
and ( n3363 , n3361 , n3362 );
nor ( n3364 , n3360 , n3363 );
not ( n3365 , n3364 );
and ( n3366 , n3359 , n3365 );
not ( n3367 , n3359 );
and ( n3368 , n3367 , n3364 );
nor ( n3369 , n3366 , n3368 );
and ( n3370 , n1533 , n1405 );
not ( n3371 , n1533 );
not ( n3372 , n1405 );
and ( n3373 , n3371 , n3372 );
nor ( n3374 , n3370 , n3373 );
and ( n3375 , n1149 , n1277 );
not ( n3376 , n1149 );
not ( n3377 , n1277 );
and ( n3378 , n3376 , n3377 );
nor ( n3379 , n3375 , n3378 );
not ( n3380 , n3379 );
and ( n3381 , n3374 , n3380 );
not ( n3382 , n3374 );
and ( n3383 , n3382 , n3379 );
nor ( n3384 , n3381 , n3383 );
nand ( n3385 , n3369 , n3384 );
xor ( n3386 , n1407 , n1535 );
not ( n3387 , n3386 );
and ( n3388 , n1151 , n1279 );
not ( n3389 , n1151 );
not ( n3390 , n1279 );
and ( n3391 , n3389 , n3390 );
nor ( n3392 , n3388 , n3391 );
not ( n3393 , n3392 );
or ( n3394 , n3387 , n3393 );
and ( n3395 , n1151 , n1279 );
not ( n3396 , n1151 );
and ( n3397 , n3396 , n3390 );
nor ( n3398 , n3395 , n3397 );
or ( n3399 , n3398 , n3386 );
nand ( n3400 , n3394 , n3399 );
not ( n3401 , n1150 );
and ( n3402 , n1278 , n3401 );
not ( n3403 , n1278 );
and ( n3404 , n3403 , n1150 );
nor ( n3405 , n3402 , n3404 );
and ( n3406 , n1406 , n1534 );
not ( n3407 , n1406 );
not ( n3408 , n1534 );
and ( n3409 , n3407 , n3408 );
nor ( n3410 , n3406 , n3409 );
and ( n3411 , n3405 , n3410 );
not ( n3412 , n3405 );
not ( n3413 , n3410 );
and ( n3414 , n3412 , n3413 );
nor ( n3415 , n3411 , n3414 );
nand ( n3416 , n3400 , n3415 );
nor ( n3417 , n3385 , n3416 );
nand ( n3418 , n3358 , n3417 );
not ( n3419 , n1414 );
nand ( n3420 , n3419 , n1542 );
not ( n3421 , n1542 );
nand ( n3422 , n3421 , n1414 );
nand ( n3423 , n3420 , n3422 );
and ( n3424 , n1158 , n1286 );
not ( n3425 , n1158 );
not ( n3426 , n1286 );
and ( n3427 , n3425 , n3426 );
nor ( n3428 , n3424 , n3427 );
or ( n3429 , n3423 , n3428 );
not ( n3430 , n3422 );
not ( n3431 , n3420 );
or ( n3432 , n3430 , n3431 );
nand ( n3433 , n3432 , n3428 );
nand ( n3434 , n3429 , n3433 );
and ( n3435 , n1159 , n1287 );
not ( n3436 , n1159 );
not ( n3437 , n1287 );
and ( n3438 , n3436 , n3437 );
nor ( n3439 , n3435 , n3438 );
not ( n3440 , n3439 );
not ( n3441 , n1415 );
nand ( n3442 , n3441 , n1543 );
not ( n3443 , n1543 );
nand ( n3444 , n3443 , n1415 );
nand ( n3445 , n3442 , n3444 );
not ( n3446 , n3445 );
or ( n3447 , n3440 , n3446 );
and ( n3448 , n1159 , n1287 );
not ( n3449 , n1159 );
and ( n3450 , n3449 , n3437 );
nor ( n3451 , n3448 , n3450 );
nand ( n3452 , n3444 , n3442 );
or ( n3453 , n3451 , n3452 );
nand ( n3454 , n3447 , n3453 );
nand ( n3455 , n3434 , n3454 );
not ( n3456 , n1156 );
nand ( n3457 , n3456 , n1540 );
not ( n3458 , n1540 );
nand ( n3459 , n3458 , n1156 );
nand ( n3460 , n3457 , n3459 );
and ( n3461 , n1284 , n1412 );
not ( n3462 , n1284 );
not ( n3463 , n1412 );
and ( n3464 , n3462 , n3463 );
nor ( n3465 , n3461 , n3464 );
or ( n3466 , n3460 , n3465 );
not ( n3467 , n1156 );
not ( n3468 , n3458 );
or ( n3469 , n3467 , n3468 );
nand ( n3470 , n3469 , n3457 );
nand ( n3471 , n3470 , n3465 );
nand ( n3472 , n3466 , n3471 );
and ( n3473 , n1157 , n1285 );
not ( n3474 , n1157 );
not ( n3475 , n1285 );
and ( n3476 , n3474 , n3475 );
nor ( n3477 , n3473 , n3476 );
not ( n3478 , n3477 );
xor ( n3479 , n1413 , n1541 );
not ( n3480 , n3479 );
or ( n3481 , n3478 , n3480 );
and ( n3482 , n1157 , n1285 );
not ( n3483 , n1157 );
and ( n3484 , n3483 , n3475 );
nor ( n3485 , n3482 , n3484 );
xor ( n3486 , n1413 , n1541 );
or ( n3487 , n3485 , n3486 );
nand ( n3488 , n3481 , n3487 );
nand ( n3489 , n3472 , n3488 );
nor ( n3490 , n3455 , n3489 );
not ( n3491 , n1163 );
nand ( n3492 , n3491 , n1547 );
not ( n3493 , n1547 );
nand ( n3494 , n3493 , n1163 );
nand ( n3495 , n3492 , n3494 );
and ( n3496 , n1291 , n1419 );
not ( n3497 , n1291 );
not ( n3498 , n1419 );
and ( n3499 , n3497 , n3498 );
nor ( n3500 , n3496 , n3499 );
or ( n3501 , n3495 , n3500 );
not ( n3502 , n3494 );
not ( n3503 , n3492 );
or ( n3504 , n3502 , n3503 );
nand ( n3505 , n3504 , n3500 );
nand ( n3506 , n3501 , n3505 );
not ( n3507 , n1290 );
and ( n3508 , n1418 , n3507 );
not ( n3509 , n1418 );
and ( n3510 , n3509 , n1290 );
nor ( n3511 , n3508 , n3510 );
and ( n3512 , n1546 , n1162 );
not ( n3513 , n1546 );
not ( n3514 , n1162 );
and ( n3515 , n3513 , n3514 );
nor ( n3516 , n3512 , n3515 );
and ( n3517 , n3511 , n3516 );
not ( n3518 , n3511 );
not ( n3519 , n3516 );
and ( n3520 , n3518 , n3519 );
nor ( n3521 , n3517 , n3520 );
nand ( n3522 , n3506 , n3521 );
xor ( n3523 , n1289 , n1417 );
not ( n3524 , n1161 );
not ( n3525 , n1545 );
not ( n3526 , n3525 );
or ( n3527 , n3524 , n3526 );
not ( n3528 , n1161 );
nand ( n3529 , n3528 , n1545 );
nand ( n3530 , n3527 , n3529 );
or ( n3531 , n3523 , n3530 );
xor ( n3532 , n1417 , n1289 );
not ( n3533 , n1161 );
not ( n3534 , n3525 );
or ( n3535 , n3533 , n3534 );
nand ( n3536 , n3535 , n3529 );
nand ( n3537 , n3532 , n3536 );
nand ( n3538 , n3531 , n3537 );
and ( n3539 , n1288 , n1416 );
not ( n3540 , n1288 );
not ( n3541 , n1416 );
and ( n3542 , n3540 , n3541 );
nor ( n3543 , n3539 , n3542 );
not ( n3544 , n3543 );
and ( n3545 , n1160 , n1544 );
not ( n3546 , n1160 );
not ( n3547 , n1544 );
and ( n3548 , n3546 , n3547 );
nor ( n3549 , n3545 , n3548 );
not ( n3550 , n3549 );
or ( n3551 , n3544 , n3550 );
and ( n3552 , n1288 , n1416 );
not ( n3553 , n1288 );
and ( n3554 , n3553 , n3541 );
nor ( n3555 , n3552 , n3554 );
and ( n3556 , n1160 , n1544 );
not ( n3557 , n1160 );
and ( n3558 , n3557 , n3547 );
nor ( n3559 , n3556 , n3558 );
or ( n3560 , n3555 , n3559 );
nand ( n3561 , n3551 , n3560 );
nand ( n3562 , n3538 , n3561 );
nor ( n3563 , n3522 , n3562 );
nand ( n3564 , n3490 , n3563 );
nor ( n3565 , n3418 , n3564 );
nand ( n3566 , n3293 , n3565 );
not ( n3567 , n3566 );
and ( n3568 , n2576 , n3019 , n3567 );
not ( n3569 , n1406 );
nand ( n3570 , n3569 , n1269 );
nor ( n3571 , n3568 , n3570 );
buf ( n3572 , n3571 );
buf ( n3573 , n3572 );
not ( n3574 , n2442 );
not ( n3575 , n2323 );
or ( n3576 , n1160 , n1546 );
nand ( n3577 , n3574 , n3575 , n3576 );
not ( n3578 , n2179 );
not ( n3579 , n2573 );
nand ( n3580 , n3578 , n3579 );
nor ( n3581 , n3577 , n3580 );
nand ( n3582 , n3581 , n3019 );
not ( n3583 , n2046 );
nand ( n3584 , n3567 , n3583 );
nor ( n3585 , n3582 , n3584 );
buf ( n3586 , n3585 );
buf ( n3587 , n3586 );
nor ( n3588 , n3018 , n3566 );
nand ( n3589 , n3588 , n2576 );
buf ( n3590 , n3589 );
buf ( n3591 , n3590 );
not ( n3592 , n3589 );
buf ( n3593 , n3592 );
buf ( n3594 , n3593 );
buf ( n3595 , n3592 );
buf ( n3596 , n3595 );
endmodule

