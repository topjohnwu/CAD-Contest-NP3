//
// Conformal-LEC Version 15.20-d250 ( 18-Apr-2016) ( 64 bit executable)
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n12345 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 ;
output n12345 ;

wire n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , 
     n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , 
     n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , 
     n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , 
     n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , 
     n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , 
     n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , 
     n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , 
     n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , 
     n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , 
     n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , 
     n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , 
     n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , 
     n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , 
     n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , 
     n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , 
     n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , 
     n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , 
     n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , 
     n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , 
     n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , 
     n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , 
     n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , 
     n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , 
     n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , 
     n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , 
     n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , 
     n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , 
     n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , 
     n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , 
     n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , 
     n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , 
     n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , 
     n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , 
     n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , 
     n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , 
     n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , 
     n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , 
     n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , 
     n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , 
     n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , 
     n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , 
     n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , 
     n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , 
     n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , 
     n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , 
     n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , 
     n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , 
     n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , 
     n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , 
     n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , 
     n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , 
     n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , 
     n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , 
     n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , 
     n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , 
     n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , 
     n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , 
     n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , 
     n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , 
     n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , 
     n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , 
     n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , 
     n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , 
     n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , 
     n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , 
     n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , 
     n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , 
     n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , 
     n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , 
     n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , 
     n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , 
     n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , 
     n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , 
     n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , 
     n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , 
     n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , 
     n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , 
     n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , 
     n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , 
     n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , 
     n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , 
     n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , 
     n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , 
     n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , 
     n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , 
     n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , 
     n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , 
     n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , 
     n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , 
     n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , 
     n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , 
     n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , 
     n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , 
     n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , 
     n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , 
     n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , 
     n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , 
     n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , 
     n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , 
     n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , 
     n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , 
     n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , 
     n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , 
     n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , 
     n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , 
     n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , 
     n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , 
     n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , 
     n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , 
     n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , 
     n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , 
     n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , 
     n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , 
     n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , 
     n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , 
     n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , 
     n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , 
     n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , 
     n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , 
     n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , 
     n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , 
     n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , 
     n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , 
     n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , 
     n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , 
     n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , 
     n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , 
     n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , 
     n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , 
     n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , 
     n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , 
     n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , 
     n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , 
     n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , 
     n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , 
     n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , 
     n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , 
     n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , 
     n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , 
     n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , 
     n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , 
     n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , 
     n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , 
     n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , 
     n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , 
     n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , 
     n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , 
     n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , 
     n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , 
     n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , 
     n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , 
     n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , 
     n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , 
     n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , 
     n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , 
     n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , 
     n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , 
     n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , 
     n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , 
     n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , 
     n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , 
     n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , 
     n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , 
     n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , 
     n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , 
     n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , 
     n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , 
     n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , 
     n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , 
     n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , 
     n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , 
     n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , 
     n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , 
     n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , 
     n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , 
     n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , 
     n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , 
     n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , 
     n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , 
     n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , 
     n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , 
     n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , 
     n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , 
     n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , 
     n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , 
     n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , 
     n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , 
     n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , 
     n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , 
     n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , 
     n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , 
     n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , 
     n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , 
     n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , 
     n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , 
     n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , 
     n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , 
     n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , 
     n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , 
     n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , 
     n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , 
     n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , 
     n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , 
     n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , 
     n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , 
     n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , 
     n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , 
     n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , 
     n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , 
     n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , 
     n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , 
     n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , 
     n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , 
     n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , 
     n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , 
     n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , 
     n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , 
     n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , 
     n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , 
     n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , 
     n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , 
     n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , 
     n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , 
     n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , 
     n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , 
     n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , 
     n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , 
     n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , 
     n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , 
     n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , 
     n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , 
     n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , 
     n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , 
     n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , 
     n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , 
     n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , 
     n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , 
     n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , 
     n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , 
     n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , 
     n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , 
     n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , 
     n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , 
     n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , 
     n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , 
     n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , 
     n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , 
     n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , 
     n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , 
     n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , 
     n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , 
     n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , 
     n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , 
     n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , 
     n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , 
     n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , 
     n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , 
     n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , 
     n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , 
     n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , 
     n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , 
     n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , 
     n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , 
     n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , 
     n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , 
     n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , 
     n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , 
     n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , 
     n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , 
     n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , 
     n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , 
     n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , 
     n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , 
     n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , 
     n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , 
     n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , 
     n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , 
     n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , 
     n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , 
     n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , 
     n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , 
     n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , 
     n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , 
     n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , 
     n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , 
     n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , 
     n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , 
     n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , 
     n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , 
     n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , 
     n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , 
     n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , 
     n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , 
     n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , 
     n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , 
     n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , 
     n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , 
     n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , 
     n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , 
     n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , 
     n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , 
     n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , 
     n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , 
     n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , 
     n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , 
     n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 ;
buf ( n12345 , n4090 );
buf ( n1026 , n322 );
buf ( n1027 , n504 );
buf ( n1028 , n37 );
buf ( n1029 , n287 );
buf ( n1030 , n365 );
buf ( n1031 , n499 );
buf ( n1032 , n47 );
buf ( n1033 , n95 );
buf ( n1034 , n8 );
buf ( n1035 , n87 );
buf ( n1036 , n470 );
buf ( n1037 , n507 );
buf ( n1038 , n410 );
buf ( n1039 , n58 );
buf ( n1040 , n361 );
buf ( n1041 , n479 );
buf ( n1042 , n320 );
buf ( n1043 , n221 );
buf ( n1044 , n466 );
buf ( n1045 , n492 );
buf ( n1046 , n211 );
buf ( n1047 , n483 );
buf ( n1048 , n426 );
buf ( n1049 , n55 );
buf ( n1050 , n321 );
buf ( n1051 , n458 );
buf ( n1052 , n50 );
buf ( n1053 , n510 );
buf ( n1054 , n407 );
buf ( n1055 , n427 );
buf ( n1056 , n378 );
buf ( n1057 , n461 );
buf ( n1058 , n175 );
buf ( n1059 , n350 );
buf ( n1060 , n445 );
buf ( n1061 , n398 );
buf ( n1062 , n255 );
buf ( n1063 , n425 );
buf ( n1064 , n292 );
buf ( n1065 , n105 );
buf ( n1066 , n220 );
buf ( n1067 , n157 );
buf ( n1068 , n3 );
buf ( n1069 , n178 );
buf ( n1070 , n282 );
buf ( n1071 , n450 );
buf ( n1072 , n349 );
buf ( n1073 , n477 );
buf ( n1074 , n207 );
buf ( n1075 , n100 );
buf ( n1076 , n63 );
buf ( n1077 , n143 );
buf ( n1078 , n132 );
buf ( n1079 , n21 );
buf ( n1080 , n66 );
buf ( n1081 , n366 );
buf ( n1082 , n163 );
buf ( n1083 , n460 );
buf ( n1084 , n12 );
buf ( n1085 , n311 );
buf ( n1086 , n43 );
buf ( n1087 , n198 );
buf ( n1088 , n503 );
buf ( n1089 , n242 );
buf ( n1090 , n338 );
buf ( n1091 , n179 );
buf ( n1092 , n284 );
buf ( n1093 , n181 );
buf ( n1094 , n167 );
buf ( n1095 , n414 );
buf ( n1096 , n363 );
buf ( n1097 , n120 );
buf ( n1098 , n229 );
buf ( n1099 , n44 );
buf ( n1100 , n233 );
buf ( n1101 , n454 );
buf ( n1102 , n155 );
buf ( n1103 , n62 );
buf ( n1104 , n502 );
buf ( n1105 , n191 );
buf ( n1106 , n131 );
buf ( n1107 , n85 );
buf ( n1108 , n272 );
buf ( n1109 , n468 );
buf ( n1110 , n144 );
buf ( n1111 , n230 );
buf ( n1112 , n437 );
buf ( n1113 , n319 );
buf ( n1114 , n441 );
buf ( n1115 , n164 );
buf ( n1116 , n374 );
buf ( n1117 , n283 );
buf ( n1118 , n145 );
buf ( n1119 , n362 );
buf ( n1120 , n395 );
buf ( n1121 , n423 );
buf ( n1122 , n11 );
buf ( n1123 , n182 );
buf ( n1124 , n253 );
buf ( n1125 , n23 );
buf ( n1126 , n343 );
buf ( n1127 , n420 );
buf ( n1128 , n278 );
buf ( n1129 , n259 );
buf ( n1130 , n422 );
buf ( n1131 , n86 );
buf ( n1132 , n109 );
buf ( n1133 , n367 );
buf ( n1134 , n162 );
buf ( n1135 , n188 );
buf ( n1136 , n108 );
buf ( n1137 , n302 );
buf ( n1138 , n34 );
buf ( n1139 , n210 );
buf ( n1140 , n315 );
buf ( n1141 , n435 );
buf ( n1142 , n462 );
buf ( n1143 , n99 );
buf ( n1144 , n139 );
buf ( n1145 , n56 );
buf ( n1146 , n61 );
buf ( n1147 , n430 );
buf ( n1148 , n506 );
buf ( n1149 , n476 );
buf ( n1150 , n102 );
buf ( n1151 , n224 );
buf ( n1152 , n176 );
buf ( n1153 , n324 );
buf ( n1154 , n300 );
buf ( n1155 , n478 );
buf ( n1156 , n29 );
buf ( n1157 , n485 );
buf ( n1158 , n303 );
buf ( n1159 , n40 );
buf ( n1160 , n455 );
buf ( n1161 , n383 );
buf ( n1162 , n281 );
buf ( n1163 , n151 );
buf ( n1164 , n413 );
buf ( n1165 , n399 );
buf ( n1166 , n74 );
buf ( n1167 , n314 );
buf ( n1168 , n228 );
buf ( n1169 , n28 );
buf ( n1170 , n4 );
buf ( n1171 , n20 );
buf ( n1172 , n152 );
buf ( n1173 , n391 );
buf ( n1174 , n490 );
buf ( n1175 , n469 );
buf ( n1176 , n463 );
buf ( n1177 , n439 );
buf ( n1178 , n204 );
buf ( n1179 , n360 );
buf ( n1180 , n273 );
buf ( n1181 , n190 );
buf ( n1182 , n46 );
buf ( n1183 , n444 );
buf ( n1184 , n429 );
buf ( n1185 , n341 );
buf ( n1186 , n72 );
buf ( n1187 , n16 );
buf ( n1188 , n354 );
buf ( n1189 , n71 );
buf ( n1190 , n205 );
buf ( n1191 , n262 );
buf ( n1192 , n345 );
buf ( n1193 , n70 );
buf ( n1194 , n482 );
buf ( n1195 , n505 );
buf ( n1196 , n417 );
buf ( n1197 , n370 );
buf ( n1198 , n474 );
buf ( n1199 , n51 );
buf ( n1200 , n150 );
buf ( n1201 , n161 );
buf ( n1202 , n305 );
buf ( n1203 , n243 );
buf ( n1204 , n187 );
buf ( n1205 , n307 );
buf ( n1206 , n432 );
buf ( n1207 , n472 );
buf ( n1208 , n235 );
buf ( n1209 , n236 );
buf ( n1210 , n298 );
buf ( n1211 , n271 );
buf ( n1212 , n177 );
buf ( n1213 , n434 );
buf ( n1214 , n484 );
buf ( n1215 , n285 );
buf ( n1216 , n133 );
buf ( n1217 , n0 );
buf ( n1218 , n369 );
buf ( n1219 , n380 );
buf ( n1220 , n418 );
buf ( n1221 , n270 );
buf ( n1222 , n291 );
buf ( n1223 , n156 );
buf ( n1224 , n39 );
buf ( n1225 , n306 );
buf ( n1226 , n327 );
buf ( n1227 , n339 );
buf ( n1228 , n401 );
buf ( n1229 , n333 );
buf ( n1230 , n489 );
buf ( n1231 , n388 );
buf ( n1232 , n27 );
buf ( n1233 , n83 );
buf ( n1234 , n421 );
buf ( n1235 , n377 );
buf ( n1236 , n41 );
buf ( n1237 , n433 );
buf ( n1238 , n397 );
buf ( n1239 , n215 );
buf ( n1240 , n405 );
buf ( n1241 , n128 );
buf ( n1242 , n153 );
buf ( n1243 , n326 );
buf ( n1244 , n265 );
buf ( n1245 , n53 );
buf ( n1246 , n185 );
buf ( n1247 , n473 );
buf ( n1248 , n386 );
buf ( n1249 , n332 );
buf ( n1250 , n57 );
buf ( n1251 , n192 );
buf ( n1252 , n238 );
buf ( n1253 , n330 );
buf ( n1254 , n389 );
buf ( n1255 , n15 );
buf ( n1256 , n25 );
buf ( n1257 , n5 );
buf ( n1258 , n246 );
buf ( n1259 , n487 );
buf ( n1260 , n411 );
buf ( n1261 , n36 );
buf ( n1262 , n353 );
buf ( n1263 , n250 );
buf ( n1264 , n45 );
buf ( n1265 , n475 );
buf ( n1266 , n309 );
buf ( n1267 , n344 );
buf ( n1268 , n486 );
buf ( n1269 , n9 );
buf ( n1270 , n125 );
buf ( n1271 , n500 );
buf ( n1272 , n31 );
buf ( n1273 , n301 );
buf ( n1274 , n275 );
buf ( n1275 , n358 );
buf ( n1276 , n313 );
buf ( n1277 , n464 );
buf ( n1278 , n480 );
buf ( n1279 , n196 );
buf ( n1280 , n440 );
buf ( n1281 , n154 );
buf ( n1282 , n7 );
buf ( n1283 , n206 );
buf ( n1284 , n184 );
buf ( n1285 , n19 );
buf ( n1286 , n82 );
buf ( n1287 , n328 );
buf ( n1288 , n356 );
buf ( n1289 , n64 );
buf ( n1290 , n295 );
buf ( n1291 , n274 );
buf ( n1292 , n497 );
buf ( n1293 , n113 );
buf ( n1294 , n160 );
buf ( n1295 , n222 );
buf ( n1296 , n142 );
buf ( n1297 , n32 );
buf ( n1298 , n80 );
buf ( n1299 , n194 );
buf ( n1300 , n171 );
buf ( n1301 , n90 );
buf ( n1302 , n213 );
buf ( n1303 , n260 );
buf ( n1304 , n403 );
buf ( n1305 , n118 );
buf ( n1306 , n357 );
buf ( n1307 , n467 );
buf ( n1308 , n508 );
buf ( n1309 , n289 );
buf ( n1310 , n38 );
buf ( n1311 , n111 );
buf ( n1312 , n304 );
buf ( n1313 , n141 );
buf ( n1314 , n384 );
buf ( n1315 , n294 );
buf ( n1316 , n376 );
buf ( n1317 , n225 );
buf ( n1318 , n481 );
buf ( n1319 , n355 );
buf ( n1320 , n130 );
buf ( n1321 , n104 );
buf ( n1322 , n112 );
buf ( n1323 , n135 );
buf ( n1324 , n195 );
buf ( n1325 , n138 );
buf ( n1326 , n134 );
buf ( n1327 , n453 );
buf ( n1328 , n79 );
buf ( n1329 , n310 );
buf ( n1330 , n340 );
buf ( n1331 , n402 );
buf ( n1332 , n52 );
buf ( n1333 , n494 );
buf ( n1334 , n200 );
buf ( n1335 , n73 );
buf ( n1336 , n452 );
buf ( n1337 , n96 );
buf ( n1338 , n335 );
buf ( n1339 , n269 );
buf ( n1340 , n256 );
buf ( n1341 , n258 );
buf ( n1342 , n148 );
buf ( n1343 , n416 );
buf ( n1344 , n347 );
buf ( n1345 , n122 );
buf ( n1346 , n312 );
buf ( n1347 , n251 );
buf ( n1348 , n35 );
buf ( n1349 , n202 );
buf ( n1350 , n495 );
buf ( n1351 , n442 );
buf ( n1352 , n170 );
buf ( n1353 , n216 );
buf ( n1354 , n448 );
buf ( n1355 , n237 );
buf ( n1356 , n17 );
buf ( n1357 , n183 );
buf ( n1358 , n18 );
buf ( n1359 , n121 );
buf ( n1360 , n438 );
buf ( n1361 , n174 );
buf ( n1362 , n14 );
buf ( n1363 , n498 );
buf ( n1364 , n231 );
buf ( n1365 , n446 );
buf ( n1366 , n373 );
buf ( n1367 , n60 );
buf ( n1368 , n436 );
buf ( n1369 , n81 );
buf ( n1370 , n78 );
buf ( n1371 , n197 );
buf ( n1372 , n77 );
buf ( n1373 , n124 );
buf ( n1374 , n30 );
buf ( n1375 , n232 );
buf ( n1376 , n227 );
buf ( n1377 , n173 );
buf ( n1378 , n263 );
buf ( n1379 , n189 );
buf ( n1380 , n234 );
buf ( n1381 , n290 );
buf ( n1382 , n293 );
buf ( n1383 , n49 );
buf ( n1384 , n98 );
buf ( n1385 , n158 );
buf ( n1386 , n254 );
buf ( n1387 , n409 );
buf ( n1388 , n68 );
buf ( n1389 , n299 );
buf ( n1390 , n115 );
buf ( n1391 , n123 );
buf ( n1392 , n396 );
buf ( n1393 , n65 );
buf ( n1394 , n449 );
buf ( n1395 , n511 );
buf ( n1396 , n13 );
buf ( n1397 , n400 );
buf ( n1398 , n10 );
buf ( n1399 , n316 );
buf ( n1400 , n336 );
buf ( n1401 , n91 );
buf ( n1402 , n146 );
buf ( n1403 , n509 );
buf ( n1404 , n193 );
buf ( n1405 , n149 );
buf ( n1406 , n266 );
buf ( n1407 , n59 );
buf ( n1408 , n267 );
buf ( n1409 , n408 );
buf ( n1410 , n218 );
buf ( n1411 , n471 );
buf ( n1412 , n415 );
buf ( n1413 , n404 );
buf ( n1414 , n257 );
buf ( n1415 , n296 );
buf ( n1416 , n75 );
buf ( n1417 , n465 );
buf ( n1418 , n346 );
buf ( n1419 , n491 );
buf ( n1420 , n371 );
buf ( n1421 , n223 );
buf ( n1422 , n217 );
buf ( n1423 , n342 );
buf ( n1424 , n240 );
buf ( n1425 , n394 );
buf ( n1426 , n372 );
buf ( n1427 , n93 );
buf ( n1428 , n103 );
buf ( n1429 , n387 );
buf ( n1430 , n268 );
buf ( n1431 , n114 );
buf ( n1432 , n459 );
buf ( n1433 , n219 );
buf ( n1434 , n101 );
buf ( n1435 , n126 );
buf ( n1436 , n501 );
buf ( n1437 , n48 );
buf ( n1438 , n119 );
buf ( n1439 , n172 );
buf ( n1440 , n42 );
buf ( n1441 , n24 );
buf ( n1442 , n385 );
buf ( n1443 , n168 );
buf ( n1444 , n456 );
buf ( n1445 , n226 );
buf ( n1446 , n488 );
buf ( n1447 , n140 );
buf ( n1448 , n247 );
buf ( n1449 , n214 );
buf ( n1450 , n106 );
buf ( n1451 , n352 );
buf ( n1452 , n428 );
buf ( n1453 , n412 );
buf ( n1454 , n348 );
buf ( n1455 , n212 );
buf ( n1456 , n379 );
buf ( n1457 , n241 );
buf ( n1458 , n166 );
buf ( n1459 , n286 );
buf ( n1460 , n84 );
buf ( n1461 , n248 );
buf ( n1462 , n89 );
buf ( n1463 , n390 );
buf ( n1464 , n6 );
buf ( n1465 , n244 );
buf ( n1466 , n451 );
buf ( n1467 , n264 );
buf ( n1468 , n2 );
buf ( n1469 , n277 );
buf ( n1470 , n199 );
buf ( n1471 , n26 );
buf ( n1472 , n67 );
buf ( n1473 , n165 );
buf ( n1474 , n186 );
buf ( n1475 , n239 );
buf ( n1476 , n159 );
buf ( n1477 , n443 );
buf ( n1478 , n447 );
buf ( n1479 , n208 );
buf ( n1480 , n318 );
buf ( n1481 , n457 );
buf ( n1482 , n169 );
buf ( n1483 , n107 );
buf ( n1484 , n368 );
buf ( n1485 , n297 );
buf ( n1486 , n1 );
buf ( n1487 , n92 );
buf ( n1488 , n392 );
buf ( n1489 , n203 );
buf ( n1490 , n88 );
buf ( n1491 , n496 );
buf ( n1492 , n382 );
buf ( n1493 , n279 );
buf ( n1494 , n331 );
buf ( n1495 , n393 );
buf ( n1496 , n280 );
buf ( n1497 , n249 );
buf ( n1498 , n97 );
buf ( n1499 , n325 );
buf ( n1500 , n261 );
buf ( n1501 , n406 );
buf ( n1502 , n334 );
buf ( n1503 , n117 );
buf ( n1504 , n375 );
buf ( n1505 , n351 );
buf ( n1506 , n137 );
buf ( n1507 , n129 );
buf ( n1508 , n76 );
buf ( n1509 , n317 );
buf ( n1510 , n337 );
buf ( n1511 , n329 );
buf ( n1512 , n381 );
buf ( n1513 , n209 );
buf ( n1514 , n22 );
buf ( n1515 , n94 );
buf ( n1516 , n136 );
buf ( n1517 , n245 );
buf ( n1518 , n201 );
buf ( n1519 , n33 );
buf ( n1520 , n493 );
buf ( n1521 , n180 );
buf ( n1522 , n431 );
buf ( n1523 , n252 );
buf ( n1524 , n359 );
buf ( n1525 , n276 );
buf ( n1526 , n110 );
buf ( n1527 , n323 );
buf ( n1528 , n419 );
buf ( n1529 , n69 );
buf ( n1530 , n308 );
buf ( n1531 , n424 );
buf ( n1532 , n147 );
buf ( n1533 , n54 );
buf ( n1534 , n364 );
buf ( n1535 , n288 );
buf ( n1536 , n116 );
buf ( n1537 , n127 );
buf ( n1538 , n1026 );
buf ( n1539 , n1282 );
xor ( n1540 , n1538 , n1539 );
buf ( n1541 , n1027 );
buf ( n1542 , n1283 );
and ( n1543 , n1541 , n1542 );
buf ( n1544 , n1028 );
buf ( n1545 , n1284 );
and ( n1546 , n1544 , n1545 );
buf ( n1547 , n1029 );
buf ( n1548 , n1285 );
and ( n1549 , n1547 , n1548 );
buf ( n1550 , n1030 );
buf ( n1551 , n1286 );
and ( n1552 , n1550 , n1551 );
buf ( n1553 , n1031 );
buf ( n1554 , n1287 );
and ( n1555 , n1553 , n1554 );
buf ( n1556 , n1032 );
buf ( n1557 , n1288 );
and ( n1558 , n1556 , n1557 );
buf ( n1559 , n1033 );
buf ( n1560 , n1289 );
and ( n1561 , n1559 , n1560 );
buf ( n1562 , n1034 );
buf ( n1563 , n1290 );
and ( n1564 , n1562 , n1563 );
buf ( n1565 , n1035 );
buf ( n1566 , n1291 );
and ( n1567 , n1565 , n1566 );
buf ( n1568 , n1036 );
buf ( n1569 , n1292 );
and ( n1570 , n1568 , n1569 );
buf ( n1571 , n1037 );
buf ( n1572 , n1293 );
and ( n1573 , n1571 , n1572 );
buf ( n1574 , n1038 );
buf ( n1575 , n1294 );
and ( n1576 , n1574 , n1575 );
buf ( n1577 , n1039 );
buf ( n1578 , n1295 );
and ( n1579 , n1577 , n1578 );
buf ( n1580 , n1040 );
buf ( n1581 , n1296 );
and ( n1582 , n1580 , n1581 );
buf ( n1583 , n1041 );
buf ( n1584 , n1297 );
and ( n1585 , n1583 , n1584 );
buf ( n1586 , n1042 );
buf ( n1587 , n1298 );
and ( n1588 , n1586 , n1587 );
buf ( n1589 , n1043 );
buf ( n1590 , n1299 );
and ( n1591 , n1589 , n1590 );
buf ( n1592 , n1044 );
buf ( n1593 , n1300 );
and ( n1594 , n1592 , n1593 );
buf ( n1595 , n1045 );
buf ( n1596 , n1301 );
and ( n1597 , n1595 , n1596 );
buf ( n1598 , n1046 );
buf ( n1599 , n1302 );
and ( n1600 , n1598 , n1599 );
buf ( n1601 , n1047 );
buf ( n1602 , n1303 );
and ( n1603 , n1601 , n1602 );
buf ( n1604 , n1048 );
buf ( n1605 , n1304 );
and ( n1606 , n1604 , n1605 );
buf ( n1607 , n1049 );
buf ( n1608 , n1305 );
and ( n1609 , n1607 , n1608 );
buf ( n1610 , n1050 );
buf ( n1611 , n1306 );
and ( n1612 , n1610 , n1611 );
buf ( n1613 , n1051 );
buf ( n1614 , n1307 );
and ( n1615 , n1613 , n1614 );
buf ( n1616 , n1052 );
buf ( n1617 , n1308 );
and ( n1618 , n1616 , n1617 );
buf ( n1619 , n1053 );
buf ( n1620 , n1309 );
and ( n1621 , n1619 , n1620 );
buf ( n1622 , n1054 );
buf ( n1623 , n1310 );
and ( n1624 , n1622 , n1623 );
buf ( n1625 , n1055 );
buf ( n1626 , n1311 );
and ( n1627 , n1625 , n1626 );
buf ( n1628 , n1056 );
buf ( n1629 , n1312 );
and ( n1630 , n1628 , n1629 );
buf ( n1631 , n1057 );
buf ( n1632 , n1313 );
and ( n1633 , n1631 , n1632 );
buf ( n1634 , n1058 );
buf ( n1635 , n1314 );
and ( n1636 , n1634 , n1635 );
buf ( n1637 , n1059 );
buf ( n1638 , n1315 );
and ( n1639 , n1637 , n1638 );
buf ( n1640 , n1060 );
buf ( n1641 , n1316 );
and ( n1642 , n1640 , n1641 );
buf ( n1643 , n1061 );
buf ( n1644 , n1317 );
and ( n1645 , n1643 , n1644 );
buf ( n1646 , n1062 );
buf ( n1647 , n1318 );
and ( n1648 , n1646 , n1647 );
buf ( n1649 , n1063 );
buf ( n1650 , n1319 );
and ( n1651 , n1649 , n1650 );
buf ( n1652 , n1064 );
buf ( n1653 , n1320 );
and ( n1654 , n1652 , n1653 );
buf ( n1655 , n1065 );
buf ( n1656 , n1321 );
and ( n1657 , n1655 , n1656 );
buf ( n1658 , n1066 );
buf ( n1659 , n1322 );
and ( n1660 , n1658 , n1659 );
buf ( n1661 , n1067 );
buf ( n1662 , n1323 );
and ( n1663 , n1661 , n1662 );
buf ( n1664 , n1068 );
buf ( n1665 , n1324 );
and ( n1666 , n1664 , n1665 );
buf ( n1667 , n1069 );
buf ( n1668 , n1325 );
and ( n1669 , n1667 , n1668 );
buf ( n1670 , n1070 );
buf ( n1671 , n1326 );
and ( n1672 , n1670 , n1671 );
buf ( n1673 , n1071 );
buf ( n1674 , n1327 );
and ( n1675 , n1673 , n1674 );
buf ( n1676 , n1072 );
buf ( n1677 , n1328 );
and ( n1678 , n1676 , n1677 );
buf ( n1679 , n1073 );
buf ( n1680 , n1329 );
and ( n1681 , n1679 , n1680 );
buf ( n1682 , n1074 );
buf ( n1683 , n1330 );
and ( n1684 , n1682 , n1683 );
buf ( n1685 , n1075 );
buf ( n1686 , n1331 );
and ( n1687 , n1685 , n1686 );
buf ( n1688 , n1076 );
buf ( n1689 , n1332 );
and ( n1690 , n1688 , n1689 );
buf ( n1691 , n1077 );
buf ( n1692 , n1333 );
and ( n1693 , n1691 , n1692 );
buf ( n1694 , n1078 );
buf ( n1695 , n1334 );
and ( n1696 , n1694 , n1695 );
buf ( n1697 , n1079 );
buf ( n1698 , n1335 );
and ( n1699 , n1697 , n1698 );
buf ( n1700 , n1080 );
buf ( n1701 , n1336 );
and ( n1702 , n1700 , n1701 );
buf ( n1703 , n1081 );
buf ( n1704 , n1337 );
and ( n1705 , n1703 , n1704 );
buf ( n1706 , n1082 );
buf ( n1707 , n1338 );
and ( n1708 , n1706 , n1707 );
buf ( n1709 , n1083 );
buf ( n1710 , n1339 );
and ( n1711 , n1709 , n1710 );
buf ( n1712 , n1084 );
buf ( n1713 , n1340 );
and ( n1714 , n1712 , n1713 );
buf ( n1715 , n1085 );
buf ( n1716 , n1341 );
and ( n1717 , n1715 , n1716 );
buf ( n1718 , n1086 );
buf ( n1719 , n1342 );
and ( n1720 , n1718 , n1719 );
buf ( n1721 , n1087 );
buf ( n1722 , n1343 );
and ( n1723 , n1721 , n1722 );
buf ( n1724 , n1088 );
buf ( n1725 , n1344 );
and ( n1726 , n1724 , n1725 );
buf ( n1727 , n1089 );
buf ( n1728 , n1345 );
and ( n1729 , n1727 , n1728 );
buf ( n1730 , n1090 );
buf ( n1731 , n1346 );
and ( n1732 , n1730 , n1731 );
buf ( n1733 , n1091 );
buf ( n1734 , n1347 );
and ( n1735 , n1733 , n1734 );
buf ( n1736 , n1092 );
buf ( n1737 , n1348 );
and ( n1738 , n1736 , n1737 );
buf ( n1739 , n1093 );
buf ( n1740 , n1349 );
and ( n1741 , n1739 , n1740 );
buf ( n1742 , n1094 );
buf ( n1743 , n1350 );
and ( n1744 , n1742 , n1743 );
buf ( n1745 , n1095 );
buf ( n1746 , n1351 );
and ( n1747 , n1745 , n1746 );
buf ( n1748 , n1096 );
buf ( n1749 , n1352 );
and ( n1750 , n1748 , n1749 );
buf ( n1751 , n1097 );
buf ( n1752 , n1353 );
and ( n1753 , n1751 , n1752 );
buf ( n1754 , n1098 );
buf ( n1755 , n1354 );
and ( n1756 , n1754 , n1755 );
buf ( n1757 , n1099 );
buf ( n1758 , n1355 );
and ( n1759 , n1757 , n1758 );
buf ( n1760 , n1100 );
buf ( n1761 , n1356 );
and ( n1762 , n1760 , n1761 );
buf ( n1763 , n1101 );
buf ( n1764 , n1357 );
and ( n1765 , n1763 , n1764 );
buf ( n1766 , n1102 );
buf ( n1767 , n1358 );
and ( n1768 , n1766 , n1767 );
buf ( n1769 , n1103 );
buf ( n1770 , n1359 );
and ( n1771 , n1769 , n1770 );
buf ( n1772 , n1104 );
buf ( n1773 , n1360 );
and ( n1774 , n1772 , n1773 );
buf ( n1775 , n1105 );
buf ( n1776 , n1361 );
and ( n1777 , n1775 , n1776 );
buf ( n1778 , n1106 );
buf ( n1779 , n1362 );
and ( n1780 , n1778 , n1779 );
buf ( n1781 , n1107 );
buf ( n1782 , n1363 );
and ( n1783 , n1781 , n1782 );
buf ( n1784 , n1108 );
buf ( n1785 , n1364 );
and ( n1786 , n1784 , n1785 );
buf ( n1787 , n1109 );
buf ( n1788 , n1365 );
and ( n1789 , n1787 , n1788 );
buf ( n1790 , n1110 );
buf ( n1791 , n1366 );
and ( n1792 , n1790 , n1791 );
buf ( n1793 , n1111 );
buf ( n1794 , n1367 );
and ( n1795 , n1793 , n1794 );
buf ( n1796 , n1112 );
buf ( n1797 , n1368 );
and ( n1798 , n1796 , n1797 );
buf ( n1799 , n1113 );
buf ( n1800 , n1369 );
and ( n1801 , n1799 , n1800 );
buf ( n1802 , n1114 );
buf ( n1803 , n1370 );
and ( n1804 , n1802 , n1803 );
buf ( n1805 , n1115 );
buf ( n1806 , n1371 );
and ( n1807 , n1805 , n1806 );
buf ( n1808 , n1116 );
buf ( n1809 , n1372 );
and ( n1810 , n1808 , n1809 );
buf ( n1811 , n1117 );
buf ( n1812 , n1373 );
and ( n1813 , n1811 , n1812 );
buf ( n1814 , n1118 );
buf ( n1815 , n1374 );
and ( n1816 , n1814 , n1815 );
buf ( n1817 , n1119 );
buf ( n1818 , n1375 );
and ( n1819 , n1817 , n1818 );
buf ( n1820 , n1120 );
buf ( n1821 , n1376 );
and ( n1822 , n1820 , n1821 );
buf ( n1823 , n1121 );
buf ( n1824 , n1377 );
and ( n1825 , n1823 , n1824 );
buf ( n1826 , n1122 );
buf ( n1827 , n1378 );
and ( n1828 , n1826 , n1827 );
buf ( n1829 , n1123 );
buf ( n1830 , n1379 );
and ( n1831 , n1829 , n1830 );
buf ( n1832 , n1124 );
buf ( n1833 , n1380 );
and ( n1834 , n1832 , n1833 );
buf ( n1835 , n1125 );
buf ( n1836 , n1381 );
and ( n1837 , n1835 , n1836 );
buf ( n1838 , n1126 );
buf ( n1839 , n1382 );
and ( n1840 , n1838 , n1839 );
buf ( n1841 , n1127 );
buf ( n1842 , n1383 );
and ( n1843 , n1841 , n1842 );
buf ( n1844 , n1128 );
buf ( n1845 , n1384 );
and ( n1846 , n1844 , n1845 );
buf ( n1847 , n1129 );
buf ( n1848 , n1385 );
and ( n1849 , n1847 , n1848 );
buf ( n1850 , n1130 );
buf ( n1851 , n1386 );
and ( n1852 , n1850 , n1851 );
buf ( n1853 , n1131 );
buf ( n1854 , n1387 );
and ( n1855 , n1853 , n1854 );
buf ( n1856 , n1132 );
buf ( n1857 , n1388 );
and ( n1858 , n1856 , n1857 );
buf ( n1859 , n1133 );
buf ( n1860 , n1389 );
and ( n1861 , n1859 , n1860 );
buf ( n1862 , n1134 );
buf ( n1863 , n1390 );
and ( n1864 , n1862 , n1863 );
buf ( n1865 , n1135 );
buf ( n1866 , n1391 );
and ( n1867 , n1865 , n1866 );
buf ( n1868 , n1136 );
buf ( n1869 , n1392 );
and ( n1870 , n1868 , n1869 );
buf ( n1871 , n1137 );
buf ( n1872 , n1393 );
and ( n1873 , n1871 , n1872 );
buf ( n1874 , n1138 );
buf ( n1875 , n1394 );
and ( n1876 , n1874 , n1875 );
buf ( n1877 , n1139 );
buf ( n1878 , n1395 );
and ( n1879 , n1877 , n1878 );
buf ( n1880 , n1140 );
buf ( n1881 , n1396 );
and ( n1882 , n1880 , n1881 );
buf ( n1883 , n1141 );
buf ( n1884 , n1397 );
and ( n1885 , n1883 , n1884 );
buf ( n1886 , n1142 );
buf ( n1887 , n1398 );
and ( n1888 , n1886 , n1887 );
buf ( n1889 , n1143 );
buf ( n1890 , n1399 );
and ( n1891 , n1889 , n1890 );
buf ( n1892 , n1144 );
buf ( n1893 , n1400 );
and ( n1894 , n1892 , n1893 );
buf ( n1895 , n1145 );
buf ( n1896 , n1401 );
and ( n1897 , n1895 , n1896 );
buf ( n1898 , n1146 );
buf ( n1899 , n1402 );
and ( n1900 , n1898 , n1899 );
buf ( n1901 , n1147 );
buf ( n1902 , n1403 );
and ( n1903 , n1901 , n1902 );
buf ( n1904 , n1148 );
buf ( n1905 , n1404 );
and ( n1906 , n1904 , n1905 );
buf ( n1907 , n1149 );
buf ( n1908 , n1405 );
and ( n1909 , n1907 , n1908 );
buf ( n1910 , n1150 );
buf ( n1911 , n1406 );
and ( n1912 , n1910 , n1911 );
buf ( n1913 , n1151 );
buf ( n1914 , n1407 );
and ( n1915 , n1913 , n1914 );
buf ( n1916 , n1152 );
buf ( n1917 , n1408 );
and ( n1918 , n1916 , n1917 );
buf ( n1919 , n1153 );
buf ( n1920 , n1409 );
and ( n1921 , n1919 , n1920 );
buf ( n1922 , n1154 );
buf ( n1923 , n1410 );
and ( n1924 , n1922 , n1923 );
buf ( n1925 , n1155 );
buf ( n1926 , n1411 );
and ( n1927 , n1925 , n1926 );
buf ( n1928 , n1156 );
buf ( n1929 , n1412 );
and ( n1930 , n1928 , n1929 );
buf ( n1931 , n1157 );
buf ( n1932 , n1413 );
and ( n1933 , n1931 , n1932 );
buf ( n1934 , n1158 );
buf ( n1935 , n1414 );
and ( n1936 , n1934 , n1935 );
buf ( n1937 , n1159 );
buf ( n1938 , n1415 );
and ( n1939 , n1937 , n1938 );
buf ( n1940 , n1160 );
buf ( n1941 , n1416 );
and ( n1942 , n1940 , n1941 );
buf ( n1943 , n1161 );
buf ( n1944 , n1417 );
and ( n1945 , n1943 , n1944 );
buf ( n1946 , n1162 );
buf ( n1947 , n1418 );
and ( n1948 , n1946 , n1947 );
buf ( n1949 , n1163 );
buf ( n1950 , n1419 );
and ( n1951 , n1949 , n1950 );
buf ( n1952 , n1164 );
buf ( n1953 , n1420 );
and ( n1954 , n1952 , n1953 );
buf ( n1955 , n1165 );
buf ( n1956 , n1421 );
and ( n1957 , n1955 , n1956 );
buf ( n1958 , n1166 );
buf ( n1959 , n1422 );
and ( n1960 , n1958 , n1959 );
buf ( n1961 , n1167 );
buf ( n1962 , n1423 );
and ( n1963 , n1961 , n1962 );
buf ( n1964 , n1168 );
buf ( n1965 , n1424 );
and ( n1966 , n1964 , n1965 );
buf ( n1967 , n1169 );
buf ( n1968 , n1425 );
and ( n1969 , n1967 , n1968 );
buf ( n1970 , n1170 );
buf ( n1971 , n1426 );
and ( n1972 , n1970 , n1971 );
buf ( n1973 , n1171 );
buf ( n1974 , n1427 );
and ( n1975 , n1973 , n1974 );
buf ( n1976 , n1172 );
buf ( n1977 , n1428 );
and ( n1978 , n1976 , n1977 );
buf ( n1979 , n1173 );
buf ( n1980 , n1429 );
and ( n1981 , n1979 , n1980 );
buf ( n1982 , n1174 );
buf ( n1983 , n1430 );
and ( n1984 , n1982 , n1983 );
buf ( n1985 , n1175 );
buf ( n1986 , n1431 );
and ( n1987 , n1985 , n1986 );
buf ( n1988 , n1176 );
buf ( n1989 , n1432 );
and ( n1990 , n1988 , n1989 );
buf ( n1991 , n1177 );
buf ( n1992 , n1433 );
and ( n1993 , n1991 , n1992 );
buf ( n1994 , n1178 );
buf ( n1995 , n1434 );
and ( n1996 , n1994 , n1995 );
buf ( n1997 , n1179 );
buf ( n1998 , n1435 );
and ( n1999 , n1997 , n1998 );
buf ( n2000 , n1180 );
buf ( n2001 , n1436 );
and ( n2002 , n2000 , n2001 );
buf ( n2003 , n1181 );
buf ( n2004 , n1437 );
and ( n2005 , n2003 , n2004 );
buf ( n2006 , n1182 );
buf ( n2007 , n1438 );
and ( n2008 , n2006 , n2007 );
buf ( n2009 , n1183 );
buf ( n2010 , n1439 );
and ( n2011 , n2009 , n2010 );
buf ( n2012 , n1184 );
buf ( n2013 , n1440 );
and ( n2014 , n2012 , n2013 );
buf ( n2015 , n1185 );
buf ( n2016 , n1441 );
and ( n2017 , n2015 , n2016 );
buf ( n2018 , n1186 );
buf ( n2019 , n1442 );
and ( n2020 , n2018 , n2019 );
buf ( n2021 , n1187 );
buf ( n2022 , n1443 );
and ( n2023 , n2021 , n2022 );
buf ( n2024 , n1188 );
buf ( n2025 , n1444 );
and ( n2026 , n2024 , n2025 );
buf ( n2027 , n1189 );
buf ( n2028 , n1445 );
and ( n2029 , n2027 , n2028 );
buf ( n2030 , n1190 );
buf ( n2031 , n1446 );
and ( n2032 , n2030 , n2031 );
buf ( n2033 , n1191 );
buf ( n2034 , n1447 );
and ( n2035 , n2033 , n2034 );
buf ( n2036 , n1192 );
buf ( n2037 , n1448 );
and ( n2038 , n2036 , n2037 );
buf ( n2039 , n1193 );
buf ( n2040 , n1449 );
and ( n2041 , n2039 , n2040 );
buf ( n2042 , n1194 );
buf ( n2043 , n1450 );
and ( n2044 , n2042 , n2043 );
buf ( n2045 , n1195 );
buf ( n2046 , n1451 );
and ( n2047 , n2045 , n2046 );
buf ( n2048 , n1196 );
buf ( n2049 , n1452 );
and ( n2050 , n2048 , n2049 );
buf ( n2051 , n1197 );
buf ( n2052 , n1453 );
and ( n2053 , n2051 , n2052 );
buf ( n2054 , n1198 );
buf ( n2055 , n1454 );
and ( n2056 , n2054 , n2055 );
buf ( n2057 , n1199 );
buf ( n2058 , n1455 );
and ( n2059 , n2057 , n2058 );
buf ( n2060 , n1200 );
buf ( n2061 , n1456 );
and ( n2062 , n2060 , n2061 );
buf ( n2063 , n1201 );
buf ( n2064 , n1457 );
and ( n2065 , n2063 , n2064 );
buf ( n2066 , n1202 );
buf ( n2067 , n1458 );
and ( n2068 , n2066 , n2067 );
buf ( n2069 , n1203 );
buf ( n2070 , n1459 );
and ( n2071 , n2069 , n2070 );
buf ( n2072 , n1204 );
buf ( n2073 , n1460 );
and ( n2074 , n2072 , n2073 );
buf ( n2075 , n1205 );
buf ( n2076 , n1461 );
and ( n2077 , n2075 , n2076 );
buf ( n2078 , n1206 );
buf ( n2079 , n1462 );
and ( n2080 , n2078 , n2079 );
buf ( n2081 , n1207 );
buf ( n2082 , n1463 );
and ( n2083 , n2081 , n2082 );
buf ( n2084 , n1208 );
buf ( n2085 , n1464 );
and ( n2086 , n2084 , n2085 );
buf ( n2087 , n1209 );
buf ( n2088 , n1465 );
and ( n2089 , n2087 , n2088 );
buf ( n2090 , n1210 );
buf ( n2091 , n1466 );
and ( n2092 , n2090 , n2091 );
buf ( n2093 , n1211 );
buf ( n2094 , n1467 );
and ( n2095 , n2093 , n2094 );
buf ( n2096 , n1212 );
buf ( n2097 , n1468 );
and ( n2098 , n2096 , n2097 );
buf ( n2099 , n1213 );
buf ( n2100 , n1469 );
and ( n2101 , n2099 , n2100 );
buf ( n2102 , n1214 );
buf ( n2103 , n1470 );
and ( n2104 , n2102 , n2103 );
buf ( n2105 , n1215 );
buf ( n2106 , n1471 );
and ( n2107 , n2105 , n2106 );
buf ( n2108 , n1216 );
buf ( n2109 , n1472 );
and ( n2110 , n2108 , n2109 );
buf ( n2111 , n1217 );
buf ( n2112 , n1473 );
and ( n2113 , n2111 , n2112 );
buf ( n2114 , n1218 );
buf ( n2115 , n1474 );
and ( n2116 , n2114 , n2115 );
buf ( n2117 , n1219 );
buf ( n2118 , n1475 );
and ( n2119 , n2117 , n2118 );
buf ( n2120 , n1220 );
buf ( n2121 , n1476 );
and ( n2122 , n2120 , n2121 );
buf ( n2123 , n1221 );
buf ( n2124 , n1477 );
and ( n2125 , n2123 , n2124 );
buf ( n2126 , n1222 );
buf ( n2127 , n1478 );
and ( n2128 , n2126 , n2127 );
buf ( n2129 , n1223 );
buf ( n2130 , n1479 );
and ( n2131 , n2129 , n2130 );
buf ( n2132 , n1224 );
buf ( n2133 , n1480 );
and ( n2134 , n2132 , n2133 );
buf ( n2135 , n1225 );
buf ( n2136 , n1481 );
and ( n2137 , n2135 , n2136 );
buf ( n2138 , n1226 );
buf ( n2139 , n1482 );
and ( n2140 , n2138 , n2139 );
buf ( n2141 , n1227 );
buf ( n2142 , n1483 );
and ( n2143 , n2141 , n2142 );
buf ( n2144 , n1228 );
buf ( n2145 , n1484 );
and ( n2146 , n2144 , n2145 );
buf ( n2147 , n1229 );
buf ( n2148 , n1485 );
and ( n2149 , n2147 , n2148 );
buf ( n2150 , n1230 );
buf ( n2151 , n1486 );
and ( n2152 , n2150 , n2151 );
buf ( n2153 , n1231 );
buf ( n2154 , n1487 );
and ( n2155 , n2153 , n2154 );
buf ( n2156 , n1232 );
buf ( n2157 , n1488 );
and ( n2158 , n2156 , n2157 );
buf ( n2159 , n1233 );
buf ( n2160 , n1489 );
and ( n2161 , n2159 , n2160 );
buf ( n2162 , n1234 );
buf ( n2163 , n1490 );
and ( n2164 , n2162 , n2163 );
buf ( n2165 , n1235 );
buf ( n2166 , n1491 );
and ( n2167 , n2165 , n2166 );
buf ( n2168 , n1236 );
buf ( n2169 , n1492 );
and ( n2170 , n2168 , n2169 );
buf ( n2171 , n1237 );
buf ( n2172 , n1493 );
and ( n2173 , n2171 , n2172 );
buf ( n2174 , n1238 );
buf ( n2175 , n1494 );
and ( n2176 , n2174 , n2175 );
buf ( n2177 , n1239 );
buf ( n2178 , n1495 );
and ( n2179 , n2177 , n2178 );
buf ( n2180 , n1240 );
buf ( n2181 , n1496 );
and ( n2182 , n2180 , n2181 );
buf ( n2183 , n1241 );
buf ( n2184 , n1497 );
and ( n2185 , n2183 , n2184 );
buf ( n2186 , n1242 );
buf ( n2187 , n1498 );
and ( n2188 , n2186 , n2187 );
buf ( n2189 , n1243 );
buf ( n2190 , n1499 );
and ( n2191 , n2189 , n2190 );
buf ( n2192 , n1244 );
buf ( n2193 , n1500 );
and ( n2194 , n2192 , n2193 );
buf ( n2195 , n1245 );
buf ( n2196 , n1501 );
and ( n2197 , n2195 , n2196 );
buf ( n2198 , n1246 );
buf ( n2199 , n1502 );
and ( n2200 , n2198 , n2199 );
buf ( n2201 , n1247 );
buf ( n2202 , n1503 );
and ( n2203 , n2201 , n2202 );
buf ( n2204 , n1248 );
buf ( n2205 , n1504 );
and ( n2206 , n2204 , n2205 );
buf ( n2207 , n1249 );
buf ( n2208 , n1505 );
and ( n2209 , n2207 , n2208 );
buf ( n2210 , n1250 );
buf ( n2211 , n1506 );
and ( n2212 , n2210 , n2211 );
buf ( n2213 , n1251 );
buf ( n2214 , n1507 );
and ( n2215 , n2213 , n2214 );
buf ( n2216 , n1252 );
buf ( n2217 , n1508 );
and ( n2218 , n2216 , n2217 );
buf ( n2219 , n1253 );
buf ( n2220 , n1509 );
and ( n2221 , n2219 , n2220 );
buf ( n2222 , n1254 );
buf ( n2223 , n1510 );
and ( n2224 , n2222 , n2223 );
buf ( n2225 , n1255 );
buf ( n2226 , n1511 );
and ( n2227 , n2225 , n2226 );
buf ( n2228 , n1256 );
buf ( n2229 , n1512 );
and ( n2230 , n2228 , n2229 );
buf ( n2231 , n1257 );
buf ( n2232 , n1513 );
and ( n2233 , n2231 , n2232 );
buf ( n2234 , n1258 );
buf ( n2235 , n1514 );
and ( n2236 , n2234 , n2235 );
buf ( n2237 , n1259 );
buf ( n2238 , n1515 );
and ( n2239 , n2237 , n2238 );
buf ( n2240 , n1260 );
buf ( n2241 , n1516 );
and ( n2242 , n2240 , n2241 );
buf ( n2243 , n1261 );
buf ( n2244 , n1517 );
and ( n2245 , n2243 , n2244 );
buf ( n2246 , n1262 );
buf ( n2247 , n1518 );
and ( n2248 , n2246 , n2247 );
buf ( n2249 , n1263 );
buf ( n2250 , n1519 );
and ( n2251 , n2249 , n2250 );
buf ( n2252 , n1264 );
buf ( n2253 , n1520 );
and ( n2254 , n2252 , n2253 );
buf ( n2255 , n1265 );
buf ( n2256 , n1521 );
and ( n2257 , n2255 , n2256 );
buf ( n2258 , n1266 );
buf ( n2259 , n1522 );
and ( n2260 , n2258 , n2259 );
buf ( n2261 , n1267 );
buf ( n2262 , n1523 );
and ( n2263 , n2261 , n2262 );
buf ( n2264 , n1268 );
buf ( n2265 , n1524 );
and ( n2266 , n2264 , n2265 );
buf ( n2267 , n1269 );
buf ( n2268 , n1525 );
and ( n2269 , n2267 , n2268 );
buf ( n2270 , n1270 );
buf ( n2271 , n1526 );
and ( n2272 , n2270 , n2271 );
buf ( n2273 , n1271 );
buf ( n2274 , n1527 );
and ( n2275 , n2273 , n2274 );
buf ( n2276 , n1272 );
buf ( n2277 , n1528 );
and ( n2278 , n2276 , n2277 );
buf ( n2279 , n1273 );
buf ( n2280 , n1529 );
and ( n2281 , n2279 , n2280 );
buf ( n2282 , n1274 );
buf ( n2283 , n1530 );
and ( n2284 , n2282 , n2283 );
buf ( n2285 , n1275 );
buf ( n2286 , n1531 );
and ( n2287 , n2285 , n2286 );
buf ( n2288 , n1276 );
buf ( n2289 , n1532 );
and ( n2290 , n2288 , n2289 );
buf ( n2291 , n1277 );
buf ( n2292 , n1533 );
and ( n2293 , n2291 , n2292 );
buf ( n2294 , n1278 );
buf ( n2295 , n1534 );
and ( n2296 , n2294 , n2295 );
buf ( n2297 , n1279 );
buf ( n2298 , n1535 );
and ( n2299 , n2297 , n2298 );
buf ( n2300 , n1280 );
buf ( n2301 , n1536 );
and ( n2302 , n2300 , n2301 );
buf ( n2303 , n1281 );
buf ( n2304 , n1537 );
and ( n2305 , n2303 , n2304 );
and ( n2306 , n2301 , n2305 );
and ( n2307 , n2300 , n2305 );
or ( n2308 , n2302 , n2306 , n2307 );
and ( n2309 , n2298 , n2308 );
and ( n2310 , n2297 , n2308 );
or ( n2311 , n2299 , n2309 , n2310 );
and ( n2312 , n2295 , n2311 );
and ( n2313 , n2294 , n2311 );
or ( n2314 , n2296 , n2312 , n2313 );
and ( n2315 , n2292 , n2314 );
and ( n2316 , n2291 , n2314 );
or ( n2317 , n2293 , n2315 , n2316 );
and ( n2318 , n2289 , n2317 );
and ( n2319 , n2288 , n2317 );
or ( n2320 , n2290 , n2318 , n2319 );
and ( n2321 , n2286 , n2320 );
and ( n2322 , n2285 , n2320 );
or ( n2323 , n2287 , n2321 , n2322 );
and ( n2324 , n2283 , n2323 );
and ( n2325 , n2282 , n2323 );
or ( n2326 , n2284 , n2324 , n2325 );
and ( n2327 , n2280 , n2326 );
and ( n2328 , n2279 , n2326 );
or ( n2329 , n2281 , n2327 , n2328 );
and ( n2330 , n2277 , n2329 );
and ( n2331 , n2276 , n2329 );
or ( n2332 , n2278 , n2330 , n2331 );
and ( n2333 , n2274 , n2332 );
and ( n2334 , n2273 , n2332 );
or ( n2335 , n2275 , n2333 , n2334 );
and ( n2336 , n2271 , n2335 );
and ( n2337 , n2270 , n2335 );
or ( n2338 , n2272 , n2336 , n2337 );
and ( n2339 , n2268 , n2338 );
and ( n2340 , n2267 , n2338 );
or ( n2341 , n2269 , n2339 , n2340 );
and ( n2342 , n2265 , n2341 );
and ( n2343 , n2264 , n2341 );
or ( n2344 , n2266 , n2342 , n2343 );
and ( n2345 , n2262 , n2344 );
and ( n2346 , n2261 , n2344 );
or ( n2347 , n2263 , n2345 , n2346 );
and ( n2348 , n2259 , n2347 );
and ( n2349 , n2258 , n2347 );
or ( n2350 , n2260 , n2348 , n2349 );
and ( n2351 , n2256 , n2350 );
and ( n2352 , n2255 , n2350 );
or ( n2353 , n2257 , n2351 , n2352 );
and ( n2354 , n2253 , n2353 );
and ( n2355 , n2252 , n2353 );
or ( n2356 , n2254 , n2354 , n2355 );
and ( n2357 , n2250 , n2356 );
and ( n2358 , n2249 , n2356 );
or ( n2359 , n2251 , n2357 , n2358 );
and ( n2360 , n2247 , n2359 );
and ( n2361 , n2246 , n2359 );
or ( n2362 , n2248 , n2360 , n2361 );
and ( n2363 , n2244 , n2362 );
and ( n2364 , n2243 , n2362 );
or ( n2365 , n2245 , n2363 , n2364 );
and ( n2366 , n2241 , n2365 );
and ( n2367 , n2240 , n2365 );
or ( n2368 , n2242 , n2366 , n2367 );
and ( n2369 , n2238 , n2368 );
and ( n2370 , n2237 , n2368 );
or ( n2371 , n2239 , n2369 , n2370 );
and ( n2372 , n2235 , n2371 );
and ( n2373 , n2234 , n2371 );
or ( n2374 , n2236 , n2372 , n2373 );
and ( n2375 , n2232 , n2374 );
and ( n2376 , n2231 , n2374 );
or ( n2377 , n2233 , n2375 , n2376 );
and ( n2378 , n2229 , n2377 );
and ( n2379 , n2228 , n2377 );
or ( n2380 , n2230 , n2378 , n2379 );
and ( n2381 , n2226 , n2380 );
and ( n2382 , n2225 , n2380 );
or ( n2383 , n2227 , n2381 , n2382 );
and ( n2384 , n2223 , n2383 );
and ( n2385 , n2222 , n2383 );
or ( n2386 , n2224 , n2384 , n2385 );
and ( n2387 , n2220 , n2386 );
and ( n2388 , n2219 , n2386 );
or ( n2389 , n2221 , n2387 , n2388 );
and ( n2390 , n2217 , n2389 );
and ( n2391 , n2216 , n2389 );
or ( n2392 , n2218 , n2390 , n2391 );
and ( n2393 , n2214 , n2392 );
and ( n2394 , n2213 , n2392 );
or ( n2395 , n2215 , n2393 , n2394 );
and ( n2396 , n2211 , n2395 );
and ( n2397 , n2210 , n2395 );
or ( n2398 , n2212 , n2396 , n2397 );
and ( n2399 , n2208 , n2398 );
and ( n2400 , n2207 , n2398 );
or ( n2401 , n2209 , n2399 , n2400 );
and ( n2402 , n2205 , n2401 );
and ( n2403 , n2204 , n2401 );
or ( n2404 , n2206 , n2402 , n2403 );
and ( n2405 , n2202 , n2404 );
and ( n2406 , n2201 , n2404 );
or ( n2407 , n2203 , n2405 , n2406 );
and ( n2408 , n2199 , n2407 );
and ( n2409 , n2198 , n2407 );
or ( n2410 , n2200 , n2408 , n2409 );
and ( n2411 , n2196 , n2410 );
and ( n2412 , n2195 , n2410 );
or ( n2413 , n2197 , n2411 , n2412 );
and ( n2414 , n2193 , n2413 );
and ( n2415 , n2192 , n2413 );
or ( n2416 , n2194 , n2414 , n2415 );
and ( n2417 , n2190 , n2416 );
and ( n2418 , n2189 , n2416 );
or ( n2419 , n2191 , n2417 , n2418 );
and ( n2420 , n2187 , n2419 );
and ( n2421 , n2186 , n2419 );
or ( n2422 , n2188 , n2420 , n2421 );
and ( n2423 , n2184 , n2422 );
and ( n2424 , n2183 , n2422 );
or ( n2425 , n2185 , n2423 , n2424 );
and ( n2426 , n2181 , n2425 );
and ( n2427 , n2180 , n2425 );
or ( n2428 , n2182 , n2426 , n2427 );
and ( n2429 , n2178 , n2428 );
and ( n2430 , n2177 , n2428 );
or ( n2431 , n2179 , n2429 , n2430 );
and ( n2432 , n2175 , n2431 );
and ( n2433 , n2174 , n2431 );
or ( n2434 , n2176 , n2432 , n2433 );
and ( n2435 , n2172 , n2434 );
and ( n2436 , n2171 , n2434 );
or ( n2437 , n2173 , n2435 , n2436 );
and ( n2438 , n2169 , n2437 );
and ( n2439 , n2168 , n2437 );
or ( n2440 , n2170 , n2438 , n2439 );
and ( n2441 , n2166 , n2440 );
and ( n2442 , n2165 , n2440 );
or ( n2443 , n2167 , n2441 , n2442 );
and ( n2444 , n2163 , n2443 );
and ( n2445 , n2162 , n2443 );
or ( n2446 , n2164 , n2444 , n2445 );
and ( n2447 , n2160 , n2446 );
and ( n2448 , n2159 , n2446 );
or ( n2449 , n2161 , n2447 , n2448 );
and ( n2450 , n2157 , n2449 );
and ( n2451 , n2156 , n2449 );
or ( n2452 , n2158 , n2450 , n2451 );
and ( n2453 , n2154 , n2452 );
and ( n2454 , n2153 , n2452 );
or ( n2455 , n2155 , n2453 , n2454 );
and ( n2456 , n2151 , n2455 );
and ( n2457 , n2150 , n2455 );
or ( n2458 , n2152 , n2456 , n2457 );
and ( n2459 , n2148 , n2458 );
and ( n2460 , n2147 , n2458 );
or ( n2461 , n2149 , n2459 , n2460 );
and ( n2462 , n2145 , n2461 );
and ( n2463 , n2144 , n2461 );
or ( n2464 , n2146 , n2462 , n2463 );
and ( n2465 , n2142 , n2464 );
and ( n2466 , n2141 , n2464 );
or ( n2467 , n2143 , n2465 , n2466 );
and ( n2468 , n2139 , n2467 );
and ( n2469 , n2138 , n2467 );
or ( n2470 , n2140 , n2468 , n2469 );
and ( n2471 , n2136 , n2470 );
and ( n2472 , n2135 , n2470 );
or ( n2473 , n2137 , n2471 , n2472 );
and ( n2474 , n2133 , n2473 );
and ( n2475 , n2132 , n2473 );
or ( n2476 , n2134 , n2474 , n2475 );
and ( n2477 , n2130 , n2476 );
and ( n2478 , n2129 , n2476 );
or ( n2479 , n2131 , n2477 , n2478 );
and ( n2480 , n2127 , n2479 );
and ( n2481 , n2126 , n2479 );
or ( n2482 , n2128 , n2480 , n2481 );
and ( n2483 , n2124 , n2482 );
and ( n2484 , n2123 , n2482 );
or ( n2485 , n2125 , n2483 , n2484 );
and ( n2486 , n2121 , n2485 );
and ( n2487 , n2120 , n2485 );
or ( n2488 , n2122 , n2486 , n2487 );
and ( n2489 , n2118 , n2488 );
and ( n2490 , n2117 , n2488 );
or ( n2491 , n2119 , n2489 , n2490 );
and ( n2492 , n2115 , n2491 );
and ( n2493 , n2114 , n2491 );
or ( n2494 , n2116 , n2492 , n2493 );
and ( n2495 , n2112 , n2494 );
and ( n2496 , n2111 , n2494 );
or ( n2497 , n2113 , n2495 , n2496 );
and ( n2498 , n2109 , n2497 );
and ( n2499 , n2108 , n2497 );
or ( n2500 , n2110 , n2498 , n2499 );
and ( n2501 , n2106 , n2500 );
and ( n2502 , n2105 , n2500 );
or ( n2503 , n2107 , n2501 , n2502 );
and ( n2504 , n2103 , n2503 );
and ( n2505 , n2102 , n2503 );
or ( n2506 , n2104 , n2504 , n2505 );
and ( n2507 , n2100 , n2506 );
and ( n2508 , n2099 , n2506 );
or ( n2509 , n2101 , n2507 , n2508 );
and ( n2510 , n2097 , n2509 );
and ( n2511 , n2096 , n2509 );
or ( n2512 , n2098 , n2510 , n2511 );
and ( n2513 , n2094 , n2512 );
and ( n2514 , n2093 , n2512 );
or ( n2515 , n2095 , n2513 , n2514 );
and ( n2516 , n2091 , n2515 );
and ( n2517 , n2090 , n2515 );
or ( n2518 , n2092 , n2516 , n2517 );
and ( n2519 , n2088 , n2518 );
and ( n2520 , n2087 , n2518 );
or ( n2521 , n2089 , n2519 , n2520 );
and ( n2522 , n2085 , n2521 );
and ( n2523 , n2084 , n2521 );
or ( n2524 , n2086 , n2522 , n2523 );
and ( n2525 , n2082 , n2524 );
and ( n2526 , n2081 , n2524 );
or ( n2527 , n2083 , n2525 , n2526 );
and ( n2528 , n2079 , n2527 );
and ( n2529 , n2078 , n2527 );
or ( n2530 , n2080 , n2528 , n2529 );
and ( n2531 , n2076 , n2530 );
and ( n2532 , n2075 , n2530 );
or ( n2533 , n2077 , n2531 , n2532 );
and ( n2534 , n2073 , n2533 );
and ( n2535 , n2072 , n2533 );
or ( n2536 , n2074 , n2534 , n2535 );
and ( n2537 , n2070 , n2536 );
and ( n2538 , n2069 , n2536 );
or ( n2539 , n2071 , n2537 , n2538 );
and ( n2540 , n2067 , n2539 );
and ( n2541 , n2066 , n2539 );
or ( n2542 , n2068 , n2540 , n2541 );
and ( n2543 , n2064 , n2542 );
and ( n2544 , n2063 , n2542 );
or ( n2545 , n2065 , n2543 , n2544 );
and ( n2546 , n2061 , n2545 );
and ( n2547 , n2060 , n2545 );
or ( n2548 , n2062 , n2546 , n2547 );
and ( n2549 , n2058 , n2548 );
and ( n2550 , n2057 , n2548 );
or ( n2551 , n2059 , n2549 , n2550 );
and ( n2552 , n2055 , n2551 );
and ( n2553 , n2054 , n2551 );
or ( n2554 , n2056 , n2552 , n2553 );
and ( n2555 , n2052 , n2554 );
and ( n2556 , n2051 , n2554 );
or ( n2557 , n2053 , n2555 , n2556 );
and ( n2558 , n2049 , n2557 );
and ( n2559 , n2048 , n2557 );
or ( n2560 , n2050 , n2558 , n2559 );
and ( n2561 , n2046 , n2560 );
and ( n2562 , n2045 , n2560 );
or ( n2563 , n2047 , n2561 , n2562 );
and ( n2564 , n2043 , n2563 );
and ( n2565 , n2042 , n2563 );
or ( n2566 , n2044 , n2564 , n2565 );
and ( n2567 , n2040 , n2566 );
and ( n2568 , n2039 , n2566 );
or ( n2569 , n2041 , n2567 , n2568 );
and ( n2570 , n2037 , n2569 );
and ( n2571 , n2036 , n2569 );
or ( n2572 , n2038 , n2570 , n2571 );
and ( n2573 , n2034 , n2572 );
and ( n2574 , n2033 , n2572 );
or ( n2575 , n2035 , n2573 , n2574 );
and ( n2576 , n2031 , n2575 );
and ( n2577 , n2030 , n2575 );
or ( n2578 , n2032 , n2576 , n2577 );
and ( n2579 , n2028 , n2578 );
and ( n2580 , n2027 , n2578 );
or ( n2581 , n2029 , n2579 , n2580 );
and ( n2582 , n2025 , n2581 );
and ( n2583 , n2024 , n2581 );
or ( n2584 , n2026 , n2582 , n2583 );
and ( n2585 , n2022 , n2584 );
and ( n2586 , n2021 , n2584 );
or ( n2587 , n2023 , n2585 , n2586 );
and ( n2588 , n2019 , n2587 );
and ( n2589 , n2018 , n2587 );
or ( n2590 , n2020 , n2588 , n2589 );
and ( n2591 , n2016 , n2590 );
and ( n2592 , n2015 , n2590 );
or ( n2593 , n2017 , n2591 , n2592 );
and ( n2594 , n2013 , n2593 );
and ( n2595 , n2012 , n2593 );
or ( n2596 , n2014 , n2594 , n2595 );
and ( n2597 , n2010 , n2596 );
and ( n2598 , n2009 , n2596 );
or ( n2599 , n2011 , n2597 , n2598 );
and ( n2600 , n2007 , n2599 );
and ( n2601 , n2006 , n2599 );
or ( n2602 , n2008 , n2600 , n2601 );
and ( n2603 , n2004 , n2602 );
and ( n2604 , n2003 , n2602 );
or ( n2605 , n2005 , n2603 , n2604 );
and ( n2606 , n2001 , n2605 );
and ( n2607 , n2000 , n2605 );
or ( n2608 , n2002 , n2606 , n2607 );
and ( n2609 , n1998 , n2608 );
and ( n2610 , n1997 , n2608 );
or ( n2611 , n1999 , n2609 , n2610 );
and ( n2612 , n1995 , n2611 );
and ( n2613 , n1994 , n2611 );
or ( n2614 , n1996 , n2612 , n2613 );
and ( n2615 , n1992 , n2614 );
and ( n2616 , n1991 , n2614 );
or ( n2617 , n1993 , n2615 , n2616 );
and ( n2618 , n1989 , n2617 );
and ( n2619 , n1988 , n2617 );
or ( n2620 , n1990 , n2618 , n2619 );
and ( n2621 , n1986 , n2620 );
and ( n2622 , n1985 , n2620 );
or ( n2623 , n1987 , n2621 , n2622 );
and ( n2624 , n1983 , n2623 );
and ( n2625 , n1982 , n2623 );
or ( n2626 , n1984 , n2624 , n2625 );
and ( n2627 , n1980 , n2626 );
and ( n2628 , n1979 , n2626 );
or ( n2629 , n1981 , n2627 , n2628 );
and ( n2630 , n1977 , n2629 );
and ( n2631 , n1976 , n2629 );
or ( n2632 , n1978 , n2630 , n2631 );
and ( n2633 , n1974 , n2632 );
and ( n2634 , n1973 , n2632 );
or ( n2635 , n1975 , n2633 , n2634 );
and ( n2636 , n1971 , n2635 );
and ( n2637 , n1970 , n2635 );
or ( n2638 , n1972 , n2636 , n2637 );
and ( n2639 , n1968 , n2638 );
and ( n2640 , n1967 , n2638 );
or ( n2641 , n1969 , n2639 , n2640 );
and ( n2642 , n1965 , n2641 );
and ( n2643 , n1964 , n2641 );
or ( n2644 , n1966 , n2642 , n2643 );
and ( n2645 , n1962 , n2644 );
and ( n2646 , n1961 , n2644 );
or ( n2647 , n1963 , n2645 , n2646 );
and ( n2648 , n1959 , n2647 );
and ( n2649 , n1958 , n2647 );
or ( n2650 , n1960 , n2648 , n2649 );
and ( n2651 , n1956 , n2650 );
and ( n2652 , n1955 , n2650 );
or ( n2653 , n1957 , n2651 , n2652 );
and ( n2654 , n1953 , n2653 );
and ( n2655 , n1952 , n2653 );
or ( n2656 , n1954 , n2654 , n2655 );
and ( n2657 , n1950 , n2656 );
and ( n2658 , n1949 , n2656 );
or ( n2659 , n1951 , n2657 , n2658 );
and ( n2660 , n1947 , n2659 );
and ( n2661 , n1946 , n2659 );
or ( n2662 , n1948 , n2660 , n2661 );
and ( n2663 , n1944 , n2662 );
and ( n2664 , n1943 , n2662 );
or ( n2665 , n1945 , n2663 , n2664 );
and ( n2666 , n1941 , n2665 );
and ( n2667 , n1940 , n2665 );
or ( n2668 , n1942 , n2666 , n2667 );
and ( n2669 , n1938 , n2668 );
and ( n2670 , n1937 , n2668 );
or ( n2671 , n1939 , n2669 , n2670 );
and ( n2672 , n1935 , n2671 );
and ( n2673 , n1934 , n2671 );
or ( n2674 , n1936 , n2672 , n2673 );
and ( n2675 , n1932 , n2674 );
and ( n2676 , n1931 , n2674 );
or ( n2677 , n1933 , n2675 , n2676 );
and ( n2678 , n1929 , n2677 );
and ( n2679 , n1928 , n2677 );
or ( n2680 , n1930 , n2678 , n2679 );
and ( n2681 , n1926 , n2680 );
and ( n2682 , n1925 , n2680 );
or ( n2683 , n1927 , n2681 , n2682 );
and ( n2684 , n1923 , n2683 );
and ( n2685 , n1922 , n2683 );
or ( n2686 , n1924 , n2684 , n2685 );
and ( n2687 , n1920 , n2686 );
and ( n2688 , n1919 , n2686 );
or ( n2689 , n1921 , n2687 , n2688 );
and ( n2690 , n1917 , n2689 );
and ( n2691 , n1916 , n2689 );
or ( n2692 , n1918 , n2690 , n2691 );
and ( n2693 , n1914 , n2692 );
and ( n2694 , n1913 , n2692 );
or ( n2695 , n1915 , n2693 , n2694 );
and ( n2696 , n1911 , n2695 );
and ( n2697 , n1910 , n2695 );
or ( n2698 , n1912 , n2696 , n2697 );
and ( n2699 , n1908 , n2698 );
and ( n2700 , n1907 , n2698 );
or ( n2701 , n1909 , n2699 , n2700 );
and ( n2702 , n1905 , n2701 );
and ( n2703 , n1904 , n2701 );
or ( n2704 , n1906 , n2702 , n2703 );
and ( n2705 , n1902 , n2704 );
and ( n2706 , n1901 , n2704 );
or ( n2707 , n1903 , n2705 , n2706 );
and ( n2708 , n1899 , n2707 );
and ( n2709 , n1898 , n2707 );
or ( n2710 , n1900 , n2708 , n2709 );
and ( n2711 , n1896 , n2710 );
and ( n2712 , n1895 , n2710 );
or ( n2713 , n1897 , n2711 , n2712 );
and ( n2714 , n1893 , n2713 );
and ( n2715 , n1892 , n2713 );
or ( n2716 , n1894 , n2714 , n2715 );
and ( n2717 , n1890 , n2716 );
and ( n2718 , n1889 , n2716 );
or ( n2719 , n1891 , n2717 , n2718 );
and ( n2720 , n1887 , n2719 );
and ( n2721 , n1886 , n2719 );
or ( n2722 , n1888 , n2720 , n2721 );
and ( n2723 , n1884 , n2722 );
and ( n2724 , n1883 , n2722 );
or ( n2725 , n1885 , n2723 , n2724 );
and ( n2726 , n1881 , n2725 );
and ( n2727 , n1880 , n2725 );
or ( n2728 , n1882 , n2726 , n2727 );
and ( n2729 , n1878 , n2728 );
and ( n2730 , n1877 , n2728 );
or ( n2731 , n1879 , n2729 , n2730 );
and ( n2732 , n1875 , n2731 );
and ( n2733 , n1874 , n2731 );
or ( n2734 , n1876 , n2732 , n2733 );
and ( n2735 , n1872 , n2734 );
and ( n2736 , n1871 , n2734 );
or ( n2737 , n1873 , n2735 , n2736 );
and ( n2738 , n1869 , n2737 );
and ( n2739 , n1868 , n2737 );
or ( n2740 , n1870 , n2738 , n2739 );
and ( n2741 , n1866 , n2740 );
and ( n2742 , n1865 , n2740 );
or ( n2743 , n1867 , n2741 , n2742 );
and ( n2744 , n1863 , n2743 );
and ( n2745 , n1862 , n2743 );
or ( n2746 , n1864 , n2744 , n2745 );
and ( n2747 , n1860 , n2746 );
and ( n2748 , n1859 , n2746 );
or ( n2749 , n1861 , n2747 , n2748 );
and ( n2750 , n1857 , n2749 );
and ( n2751 , n1856 , n2749 );
or ( n2752 , n1858 , n2750 , n2751 );
and ( n2753 , n1854 , n2752 );
and ( n2754 , n1853 , n2752 );
or ( n2755 , n1855 , n2753 , n2754 );
and ( n2756 , n1851 , n2755 );
and ( n2757 , n1850 , n2755 );
or ( n2758 , n1852 , n2756 , n2757 );
and ( n2759 , n1848 , n2758 );
and ( n2760 , n1847 , n2758 );
or ( n2761 , n1849 , n2759 , n2760 );
and ( n2762 , n1845 , n2761 );
and ( n2763 , n1844 , n2761 );
or ( n2764 , n1846 , n2762 , n2763 );
and ( n2765 , n1842 , n2764 );
and ( n2766 , n1841 , n2764 );
or ( n2767 , n1843 , n2765 , n2766 );
and ( n2768 , n1839 , n2767 );
and ( n2769 , n1838 , n2767 );
or ( n2770 , n1840 , n2768 , n2769 );
and ( n2771 , n1836 , n2770 );
and ( n2772 , n1835 , n2770 );
or ( n2773 , n1837 , n2771 , n2772 );
and ( n2774 , n1833 , n2773 );
and ( n2775 , n1832 , n2773 );
or ( n2776 , n1834 , n2774 , n2775 );
and ( n2777 , n1830 , n2776 );
and ( n2778 , n1829 , n2776 );
or ( n2779 , n1831 , n2777 , n2778 );
and ( n2780 , n1827 , n2779 );
and ( n2781 , n1826 , n2779 );
or ( n2782 , n1828 , n2780 , n2781 );
and ( n2783 , n1824 , n2782 );
and ( n2784 , n1823 , n2782 );
or ( n2785 , n1825 , n2783 , n2784 );
and ( n2786 , n1821 , n2785 );
and ( n2787 , n1820 , n2785 );
or ( n2788 , n1822 , n2786 , n2787 );
and ( n2789 , n1818 , n2788 );
and ( n2790 , n1817 , n2788 );
or ( n2791 , n1819 , n2789 , n2790 );
and ( n2792 , n1815 , n2791 );
and ( n2793 , n1814 , n2791 );
or ( n2794 , n1816 , n2792 , n2793 );
and ( n2795 , n1812 , n2794 );
and ( n2796 , n1811 , n2794 );
or ( n2797 , n1813 , n2795 , n2796 );
and ( n2798 , n1809 , n2797 );
and ( n2799 , n1808 , n2797 );
or ( n2800 , n1810 , n2798 , n2799 );
and ( n2801 , n1806 , n2800 );
and ( n2802 , n1805 , n2800 );
or ( n2803 , n1807 , n2801 , n2802 );
and ( n2804 , n1803 , n2803 );
and ( n2805 , n1802 , n2803 );
or ( n2806 , n1804 , n2804 , n2805 );
and ( n2807 , n1800 , n2806 );
and ( n2808 , n1799 , n2806 );
or ( n2809 , n1801 , n2807 , n2808 );
and ( n2810 , n1797 , n2809 );
and ( n2811 , n1796 , n2809 );
or ( n2812 , n1798 , n2810 , n2811 );
and ( n2813 , n1794 , n2812 );
and ( n2814 , n1793 , n2812 );
or ( n2815 , n1795 , n2813 , n2814 );
and ( n2816 , n1791 , n2815 );
and ( n2817 , n1790 , n2815 );
or ( n2818 , n1792 , n2816 , n2817 );
and ( n2819 , n1788 , n2818 );
and ( n2820 , n1787 , n2818 );
or ( n2821 , n1789 , n2819 , n2820 );
and ( n2822 , n1785 , n2821 );
and ( n2823 , n1784 , n2821 );
or ( n2824 , n1786 , n2822 , n2823 );
and ( n2825 , n1782 , n2824 );
and ( n2826 , n1781 , n2824 );
or ( n2827 , n1783 , n2825 , n2826 );
and ( n2828 , n1779 , n2827 );
and ( n2829 , n1778 , n2827 );
or ( n2830 , n1780 , n2828 , n2829 );
and ( n2831 , n1776 , n2830 );
and ( n2832 , n1775 , n2830 );
or ( n2833 , n1777 , n2831 , n2832 );
and ( n2834 , n1773 , n2833 );
and ( n2835 , n1772 , n2833 );
or ( n2836 , n1774 , n2834 , n2835 );
and ( n2837 , n1770 , n2836 );
and ( n2838 , n1769 , n2836 );
or ( n2839 , n1771 , n2837 , n2838 );
and ( n2840 , n1767 , n2839 );
and ( n2841 , n1766 , n2839 );
or ( n2842 , n1768 , n2840 , n2841 );
and ( n2843 , n1764 , n2842 );
and ( n2844 , n1763 , n2842 );
or ( n2845 , n1765 , n2843 , n2844 );
and ( n2846 , n1761 , n2845 );
and ( n2847 , n1760 , n2845 );
or ( n2848 , n1762 , n2846 , n2847 );
and ( n2849 , n1758 , n2848 );
and ( n2850 , n1757 , n2848 );
or ( n2851 , n1759 , n2849 , n2850 );
and ( n2852 , n1755 , n2851 );
and ( n2853 , n1754 , n2851 );
or ( n2854 , n1756 , n2852 , n2853 );
and ( n2855 , n1752 , n2854 );
and ( n2856 , n1751 , n2854 );
or ( n2857 , n1753 , n2855 , n2856 );
and ( n2858 , n1749 , n2857 );
and ( n2859 , n1748 , n2857 );
or ( n2860 , n1750 , n2858 , n2859 );
and ( n2861 , n1746 , n2860 );
and ( n2862 , n1745 , n2860 );
or ( n2863 , n1747 , n2861 , n2862 );
and ( n2864 , n1743 , n2863 );
and ( n2865 , n1742 , n2863 );
or ( n2866 , n1744 , n2864 , n2865 );
and ( n2867 , n1740 , n2866 );
and ( n2868 , n1739 , n2866 );
or ( n2869 , n1741 , n2867 , n2868 );
and ( n2870 , n1737 , n2869 );
and ( n2871 , n1736 , n2869 );
or ( n2872 , n1738 , n2870 , n2871 );
and ( n2873 , n1734 , n2872 );
and ( n2874 , n1733 , n2872 );
or ( n2875 , n1735 , n2873 , n2874 );
and ( n2876 , n1731 , n2875 );
and ( n2877 , n1730 , n2875 );
or ( n2878 , n1732 , n2876 , n2877 );
and ( n2879 , n1728 , n2878 );
and ( n2880 , n1727 , n2878 );
or ( n2881 , n1729 , n2879 , n2880 );
and ( n2882 , n1725 , n2881 );
and ( n2883 , n1724 , n2881 );
or ( n2884 , n1726 , n2882 , n2883 );
and ( n2885 , n1722 , n2884 );
and ( n2886 , n1721 , n2884 );
or ( n2887 , n1723 , n2885 , n2886 );
and ( n2888 , n1719 , n2887 );
and ( n2889 , n1718 , n2887 );
or ( n2890 , n1720 , n2888 , n2889 );
and ( n2891 , n1716 , n2890 );
and ( n2892 , n1715 , n2890 );
or ( n2893 , n1717 , n2891 , n2892 );
and ( n2894 , n1713 , n2893 );
and ( n2895 , n1712 , n2893 );
or ( n2896 , n1714 , n2894 , n2895 );
and ( n2897 , n1710 , n2896 );
and ( n2898 , n1709 , n2896 );
or ( n2899 , n1711 , n2897 , n2898 );
and ( n2900 , n1707 , n2899 );
and ( n2901 , n1706 , n2899 );
or ( n2902 , n1708 , n2900 , n2901 );
and ( n2903 , n1704 , n2902 );
and ( n2904 , n1703 , n2902 );
or ( n2905 , n1705 , n2903 , n2904 );
and ( n2906 , n1701 , n2905 );
and ( n2907 , n1700 , n2905 );
or ( n2908 , n1702 , n2906 , n2907 );
and ( n2909 , n1698 , n2908 );
and ( n2910 , n1697 , n2908 );
or ( n2911 , n1699 , n2909 , n2910 );
and ( n2912 , n1695 , n2911 );
and ( n2913 , n1694 , n2911 );
or ( n2914 , n1696 , n2912 , n2913 );
and ( n2915 , n1692 , n2914 );
and ( n2916 , n1691 , n2914 );
or ( n2917 , n1693 , n2915 , n2916 );
and ( n2918 , n1689 , n2917 );
and ( n2919 , n1688 , n2917 );
or ( n2920 , n1690 , n2918 , n2919 );
and ( n2921 , n1686 , n2920 );
and ( n2922 , n1685 , n2920 );
or ( n2923 , n1687 , n2921 , n2922 );
and ( n2924 , n1683 , n2923 );
and ( n2925 , n1682 , n2923 );
or ( n2926 , n1684 , n2924 , n2925 );
and ( n2927 , n1680 , n2926 );
and ( n2928 , n1679 , n2926 );
or ( n2929 , n1681 , n2927 , n2928 );
and ( n2930 , n1677 , n2929 );
and ( n2931 , n1676 , n2929 );
or ( n2932 , n1678 , n2930 , n2931 );
and ( n2933 , n1674 , n2932 );
and ( n2934 , n1673 , n2932 );
or ( n2935 , n1675 , n2933 , n2934 );
and ( n2936 , n1671 , n2935 );
and ( n2937 , n1670 , n2935 );
or ( n2938 , n1672 , n2936 , n2937 );
and ( n2939 , n1668 , n2938 );
and ( n2940 , n1667 , n2938 );
or ( n2941 , n1669 , n2939 , n2940 );
and ( n2942 , n1665 , n2941 );
and ( n2943 , n1664 , n2941 );
or ( n2944 , n1666 , n2942 , n2943 );
and ( n2945 , n1662 , n2944 );
and ( n2946 , n1661 , n2944 );
or ( n2947 , n1663 , n2945 , n2946 );
and ( n2948 , n1659 , n2947 );
and ( n2949 , n1658 , n2947 );
or ( n2950 , n1660 , n2948 , n2949 );
and ( n2951 , n1656 , n2950 );
and ( n2952 , n1655 , n2950 );
or ( n2953 , n1657 , n2951 , n2952 );
and ( n2954 , n1653 , n2953 );
and ( n2955 , n1652 , n2953 );
or ( n2956 , n1654 , n2954 , n2955 );
and ( n2957 , n1650 , n2956 );
and ( n2958 , n1649 , n2956 );
or ( n2959 , n1651 , n2957 , n2958 );
and ( n2960 , n1647 , n2959 );
and ( n2961 , n1646 , n2959 );
or ( n2962 , n1648 , n2960 , n2961 );
and ( n2963 , n1644 , n2962 );
and ( n2964 , n1643 , n2962 );
or ( n2965 , n1645 , n2963 , n2964 );
and ( n2966 , n1641 , n2965 );
and ( n2967 , n1640 , n2965 );
or ( n2968 , n1642 , n2966 , n2967 );
and ( n2969 , n1638 , n2968 );
and ( n2970 , n1637 , n2968 );
or ( n2971 , n1639 , n2969 , n2970 );
and ( n2972 , n1635 , n2971 );
and ( n2973 , n1634 , n2971 );
or ( n2974 , n1636 , n2972 , n2973 );
and ( n2975 , n1632 , n2974 );
and ( n2976 , n1631 , n2974 );
or ( n2977 , n1633 , n2975 , n2976 );
and ( n2978 , n1629 , n2977 );
and ( n2979 , n1628 , n2977 );
or ( n2980 , n1630 , n2978 , n2979 );
and ( n2981 , n1626 , n2980 );
and ( n2982 , n1625 , n2980 );
or ( n2983 , n1627 , n2981 , n2982 );
and ( n2984 , n1623 , n2983 );
and ( n2985 , n1622 , n2983 );
or ( n2986 , n1624 , n2984 , n2985 );
and ( n2987 , n1620 , n2986 );
and ( n2988 , n1619 , n2986 );
or ( n2989 , n1621 , n2987 , n2988 );
and ( n2990 , n1617 , n2989 );
and ( n2991 , n1616 , n2989 );
or ( n2992 , n1618 , n2990 , n2991 );
and ( n2993 , n1614 , n2992 );
and ( n2994 , n1613 , n2992 );
or ( n2995 , n1615 , n2993 , n2994 );
and ( n2996 , n1611 , n2995 );
and ( n2997 , n1610 , n2995 );
or ( n2998 , n1612 , n2996 , n2997 );
and ( n2999 , n1608 , n2998 );
and ( n3000 , n1607 , n2998 );
or ( n3001 , n1609 , n2999 , n3000 );
and ( n3002 , n1605 , n3001 );
and ( n3003 , n1604 , n3001 );
or ( n3004 , n1606 , n3002 , n3003 );
and ( n3005 , n1602 , n3004 );
and ( n3006 , n1601 , n3004 );
or ( n3007 , n1603 , n3005 , n3006 );
and ( n3008 , n1599 , n3007 );
and ( n3009 , n1598 , n3007 );
or ( n3010 , n1600 , n3008 , n3009 );
and ( n3011 , n1596 , n3010 );
and ( n3012 , n1595 , n3010 );
or ( n3013 , n1597 , n3011 , n3012 );
and ( n3014 , n1593 , n3013 );
and ( n3015 , n1592 , n3013 );
or ( n3016 , n1594 , n3014 , n3015 );
and ( n3017 , n1590 , n3016 );
and ( n3018 , n1589 , n3016 );
or ( n3019 , n1591 , n3017 , n3018 );
and ( n3020 , n1587 , n3019 );
and ( n3021 , n1586 , n3019 );
or ( n3022 , n1588 , n3020 , n3021 );
and ( n3023 , n1584 , n3022 );
and ( n3024 , n1583 , n3022 );
or ( n3025 , n1585 , n3023 , n3024 );
and ( n3026 , n1581 , n3025 );
and ( n3027 , n1580 , n3025 );
or ( n3028 , n1582 , n3026 , n3027 );
and ( n3029 , n1578 , n3028 );
and ( n3030 , n1577 , n3028 );
or ( n3031 , n1579 , n3029 , n3030 );
and ( n3032 , n1575 , n3031 );
and ( n3033 , n1574 , n3031 );
or ( n3034 , n1576 , n3032 , n3033 );
and ( n3035 , n1572 , n3034 );
and ( n3036 , n1571 , n3034 );
or ( n3037 , n1573 , n3035 , n3036 );
and ( n3038 , n1569 , n3037 );
and ( n3039 , n1568 , n3037 );
or ( n3040 , n1570 , n3038 , n3039 );
and ( n3041 , n1566 , n3040 );
and ( n3042 , n1565 , n3040 );
or ( n3043 , n1567 , n3041 , n3042 );
and ( n3044 , n1563 , n3043 );
and ( n3045 , n1562 , n3043 );
or ( n3046 , n1564 , n3044 , n3045 );
and ( n3047 , n1560 , n3046 );
and ( n3048 , n1559 , n3046 );
or ( n3049 , n1561 , n3047 , n3048 );
and ( n3050 , n1557 , n3049 );
and ( n3051 , n1556 , n3049 );
or ( n3052 , n1558 , n3050 , n3051 );
and ( n3053 , n1554 , n3052 );
and ( n3054 , n1553 , n3052 );
or ( n3055 , n1555 , n3053 , n3054 );
and ( n3056 , n1551 , n3055 );
and ( n3057 , n1550 , n3055 );
or ( n3058 , n1552 , n3056 , n3057 );
and ( n3059 , n1548 , n3058 );
and ( n3060 , n1547 , n3058 );
or ( n3061 , n1549 , n3059 , n3060 );
and ( n3062 , n1545 , n3061 );
and ( n3063 , n1544 , n3061 );
or ( n3064 , n1546 , n3062 , n3063 );
and ( n3065 , n1542 , n3064 );
and ( n3066 , n1541 , n3064 );
or ( n3067 , n1543 , n3065 , n3066 );
xor ( n3068 , n1540 , n3067 );
buf ( n3069 , n3068 );
xor ( n3070 , n1541 , n1542 );
xor ( n3071 , n3070 , n3064 );
buf ( n3072 , n3071 );
xor ( n3073 , n3069 , n3072 );
xor ( n3074 , n1544 , n1545 );
xor ( n3075 , n3074 , n3061 );
buf ( n3076 , n3075 );
xor ( n3077 , n1547 , n1548 );
xor ( n3078 , n3077 , n3058 );
buf ( n3079 , n3078 );
xor ( n3080 , n3076 , n3079 );
xor ( n3081 , n3073 , n3080 );
xor ( n3082 , n1550 , n1551 );
xor ( n3083 , n3082 , n3055 );
buf ( n3084 , n3083 );
xor ( n3085 , n1553 , n1554 );
xor ( n3086 , n3085 , n3052 );
buf ( n3087 , n3086 );
xor ( n3088 , n3084 , n3087 );
xor ( n3089 , n1556 , n1557 );
xor ( n3090 , n3089 , n3049 );
buf ( n3091 , n3090 );
xor ( n3092 , n1559 , n1560 );
xor ( n3093 , n3092 , n3046 );
buf ( n3094 , n3093 );
xor ( n3095 , n3091 , n3094 );
xor ( n3096 , n3088 , n3095 );
xor ( n3097 , n3081 , n3096 );
xor ( n3098 , n1562 , n1563 );
xor ( n3099 , n3098 , n3043 );
buf ( n3100 , n3099 );
xor ( n3101 , n1565 , n1566 );
xor ( n3102 , n3101 , n3040 );
buf ( n3103 , n3102 );
xor ( n3104 , n3100 , n3103 );
xor ( n3105 , n1568 , n1569 );
xor ( n3106 , n3105 , n3037 );
buf ( n3107 , n3106 );
xor ( n3108 , n1571 , n1572 );
xor ( n3109 , n3108 , n3034 );
buf ( n3110 , n3109 );
xor ( n3111 , n3107 , n3110 );
xor ( n3112 , n3104 , n3111 );
xor ( n3113 , n1574 , n1575 );
xor ( n3114 , n3113 , n3031 );
buf ( n3115 , n3114 );
xor ( n3116 , n1577 , n1578 );
xor ( n3117 , n3116 , n3028 );
buf ( n3118 , n3117 );
xor ( n3119 , n3115 , n3118 );
xor ( n3120 , n1580 , n1581 );
xor ( n3121 , n3120 , n3025 );
buf ( n3122 , n3121 );
xor ( n3123 , n1583 , n1584 );
xor ( n3124 , n3123 , n3022 );
buf ( n3125 , n3124 );
xor ( n3126 , n3122 , n3125 );
xor ( n3127 , n3119 , n3126 );
xor ( n3128 , n3112 , n3127 );
xor ( n3129 , n3097 , n3128 );
xor ( n3130 , n1586 , n1587 );
xor ( n3131 , n3130 , n3019 );
buf ( n3132 , n3131 );
xor ( n3133 , n1589 , n1590 );
xor ( n3134 , n3133 , n3016 );
buf ( n3135 , n3134 );
xor ( n3136 , n3132 , n3135 );
xor ( n3137 , n1592 , n1593 );
xor ( n3138 , n3137 , n3013 );
buf ( n3139 , n3138 );
xor ( n3140 , n1595 , n1596 );
xor ( n3141 , n3140 , n3010 );
buf ( n3142 , n3141 );
xor ( n3143 , n3139 , n3142 );
xor ( n3144 , n3136 , n3143 );
xor ( n3145 , n1598 , n1599 );
xor ( n3146 , n3145 , n3007 );
buf ( n3147 , n3146 );
xor ( n3148 , n1601 , n1602 );
xor ( n3149 , n3148 , n3004 );
buf ( n3150 , n3149 );
xor ( n3151 , n3147 , n3150 );
xor ( n3152 , n1604 , n1605 );
xor ( n3153 , n3152 , n3001 );
buf ( n3154 , n3153 );
xor ( n3155 , n1607 , n1608 );
xor ( n3156 , n3155 , n2998 );
buf ( n3157 , n3156 );
xor ( n3158 , n3154 , n3157 );
xor ( n3159 , n3151 , n3158 );
xor ( n3160 , n3144 , n3159 );
xor ( n3161 , n1610 , n1611 );
xor ( n3162 , n3161 , n2995 );
buf ( n3163 , n3162 );
xor ( n3164 , n1613 , n1614 );
xor ( n3165 , n3164 , n2992 );
buf ( n3166 , n3165 );
xor ( n3167 , n3163 , n3166 );
xor ( n3168 , n1616 , n1617 );
xor ( n3169 , n3168 , n2989 );
buf ( n3170 , n3169 );
xor ( n3171 , n1619 , n1620 );
xor ( n3172 , n3171 , n2986 );
buf ( n3173 , n3172 );
xor ( n3174 , n3170 , n3173 );
xor ( n3175 , n3167 , n3174 );
xor ( n3176 , n1622 , n1623 );
xor ( n3177 , n3176 , n2983 );
buf ( n3178 , n3177 );
xor ( n3179 , n1625 , n1626 );
xor ( n3180 , n3179 , n2980 );
buf ( n3181 , n3180 );
xor ( n3182 , n3178 , n3181 );
xor ( n3183 , n1628 , n1629 );
xor ( n3184 , n3183 , n2977 );
buf ( n3185 , n3184 );
xor ( n3186 , n1631 , n1632 );
xor ( n3187 , n3186 , n2974 );
buf ( n3188 , n3187 );
xor ( n3189 , n3185 , n3188 );
xor ( n3190 , n3182 , n3189 );
xor ( n3191 , n3175 , n3190 );
xor ( n3192 , n3160 , n3191 );
xor ( n3193 , n3129 , n3192 );
xor ( n3194 , n1634 , n1635 );
xor ( n3195 , n3194 , n2971 );
buf ( n3196 , n3195 );
xor ( n3197 , n1637 , n1638 );
xor ( n3198 , n3197 , n2968 );
buf ( n3199 , n3198 );
xor ( n3200 , n3196 , n3199 );
xor ( n3201 , n1640 , n1641 );
xor ( n3202 , n3201 , n2965 );
buf ( n3203 , n3202 );
xor ( n3204 , n1643 , n1644 );
xor ( n3205 , n3204 , n2962 );
buf ( n3206 , n3205 );
xor ( n3207 , n3203 , n3206 );
xor ( n3208 , n3200 , n3207 );
xor ( n3209 , n1646 , n1647 );
xor ( n3210 , n3209 , n2959 );
buf ( n3211 , n3210 );
xor ( n3212 , n1649 , n1650 );
xor ( n3213 , n3212 , n2956 );
buf ( n3214 , n3213 );
xor ( n3215 , n3211 , n3214 );
xor ( n3216 , n1652 , n1653 );
xor ( n3217 , n3216 , n2953 );
buf ( n3218 , n3217 );
xor ( n3219 , n1655 , n1656 );
xor ( n3220 , n3219 , n2950 );
buf ( n3221 , n3220 );
xor ( n3222 , n3218 , n3221 );
xor ( n3223 , n3215 , n3222 );
xor ( n3224 , n3208 , n3223 );
xor ( n3225 , n1658 , n1659 );
xor ( n3226 , n3225 , n2947 );
buf ( n3227 , n3226 );
xor ( n3228 , n1661 , n1662 );
xor ( n3229 , n3228 , n2944 );
buf ( n3230 , n3229 );
xor ( n3231 , n3227 , n3230 );
xor ( n3232 , n1664 , n1665 );
xor ( n3233 , n3232 , n2941 );
buf ( n3234 , n3233 );
xor ( n3235 , n1667 , n1668 );
xor ( n3236 , n3235 , n2938 );
buf ( n3237 , n3236 );
xor ( n3238 , n3234 , n3237 );
xor ( n3239 , n3231 , n3238 );
xor ( n3240 , n1670 , n1671 );
xor ( n3241 , n3240 , n2935 );
buf ( n3242 , n3241 );
xor ( n3243 , n1673 , n1674 );
xor ( n3244 , n3243 , n2932 );
buf ( n3245 , n3244 );
xor ( n3246 , n3242 , n3245 );
xor ( n3247 , n1676 , n1677 );
xor ( n3248 , n3247 , n2929 );
buf ( n3249 , n3248 );
xor ( n3250 , n1679 , n1680 );
xor ( n3251 , n3250 , n2926 );
buf ( n3252 , n3251 );
xor ( n3253 , n3249 , n3252 );
xor ( n3254 , n3246 , n3253 );
xor ( n3255 , n3239 , n3254 );
xor ( n3256 , n3224 , n3255 );
xor ( n3257 , n1682 , n1683 );
xor ( n3258 , n3257 , n2923 );
buf ( n3259 , n3258 );
xor ( n3260 , n1685 , n1686 );
xor ( n3261 , n3260 , n2920 );
buf ( n3262 , n3261 );
xor ( n3263 , n3259 , n3262 );
xor ( n3264 , n1688 , n1689 );
xor ( n3265 , n3264 , n2917 );
buf ( n3266 , n3265 );
xor ( n3267 , n1691 , n1692 );
xor ( n3268 , n3267 , n2914 );
buf ( n3269 , n3268 );
xor ( n3270 , n3266 , n3269 );
xor ( n3271 , n3263 , n3270 );
xor ( n3272 , n1694 , n1695 );
xor ( n3273 , n3272 , n2911 );
buf ( n3274 , n3273 );
xor ( n3275 , n1697 , n1698 );
xor ( n3276 , n3275 , n2908 );
buf ( n3277 , n3276 );
xor ( n3278 , n3274 , n3277 );
xor ( n3279 , n1700 , n1701 );
xor ( n3280 , n3279 , n2905 );
buf ( n3281 , n3280 );
xor ( n3282 , n1703 , n1704 );
xor ( n3283 , n3282 , n2902 );
buf ( n3284 , n3283 );
xor ( n3285 , n3281 , n3284 );
xor ( n3286 , n3278 , n3285 );
xor ( n3287 , n3271 , n3286 );
xor ( n3288 , n1706 , n1707 );
xor ( n3289 , n3288 , n2899 );
buf ( n3290 , n3289 );
xor ( n3291 , n1709 , n1710 );
xor ( n3292 , n3291 , n2896 );
buf ( n3293 , n3292 );
xor ( n3294 , n3290 , n3293 );
xor ( n3295 , n1712 , n1713 );
xor ( n3296 , n3295 , n2893 );
buf ( n3297 , n3296 );
xor ( n3298 , n1715 , n1716 );
xor ( n3299 , n3298 , n2890 );
buf ( n3300 , n3299 );
xor ( n3301 , n3297 , n3300 );
xor ( n3302 , n3294 , n3301 );
xor ( n3303 , n1718 , n1719 );
xor ( n3304 , n3303 , n2887 );
buf ( n3305 , n3304 );
xor ( n3306 , n1721 , n1722 );
xor ( n3307 , n3306 , n2884 );
buf ( n3308 , n3307 );
xor ( n3309 , n3305 , n3308 );
xor ( n3310 , n1724 , n1725 );
xor ( n3311 , n3310 , n2881 );
buf ( n3312 , n3311 );
xor ( n3313 , n1727 , n1728 );
xor ( n3314 , n3313 , n2878 );
buf ( n3315 , n3314 );
xor ( n3316 , n3312 , n3315 );
xor ( n3317 , n3309 , n3316 );
xor ( n3318 , n3302 , n3317 );
xor ( n3319 , n3287 , n3318 );
xor ( n3320 , n3256 , n3319 );
xor ( n3321 , n3193 , n3320 );
xor ( n3322 , n1730 , n1731 );
xor ( n3323 , n3322 , n2875 );
buf ( n3324 , n3323 );
xor ( n3325 , n1733 , n1734 );
xor ( n3326 , n3325 , n2872 );
buf ( n3327 , n3326 );
xor ( n3328 , n3324 , n3327 );
xor ( n3329 , n1736 , n1737 );
xor ( n3330 , n3329 , n2869 );
buf ( n3331 , n3330 );
xor ( n3332 , n1739 , n1740 );
xor ( n3333 , n3332 , n2866 );
buf ( n3334 , n3333 );
xor ( n3335 , n3331 , n3334 );
xor ( n3336 , n3328 , n3335 );
xor ( n3337 , n1742 , n1743 );
xor ( n3338 , n3337 , n2863 );
buf ( n3339 , n3338 );
xor ( n3340 , n1745 , n1746 );
xor ( n3341 , n3340 , n2860 );
buf ( n3342 , n3341 );
xor ( n3343 , n3339 , n3342 );
xor ( n3344 , n1748 , n1749 );
xor ( n3345 , n3344 , n2857 );
buf ( n3346 , n3345 );
xor ( n3347 , n1751 , n1752 );
xor ( n3348 , n3347 , n2854 );
buf ( n3349 , n3348 );
xor ( n3350 , n3346 , n3349 );
xor ( n3351 , n3343 , n3350 );
xor ( n3352 , n3336 , n3351 );
xor ( n3353 , n1754 , n1755 );
xor ( n3354 , n3353 , n2851 );
buf ( n3355 , n3354 );
xor ( n3356 , n1757 , n1758 );
xor ( n3357 , n3356 , n2848 );
buf ( n3358 , n3357 );
xor ( n3359 , n3355 , n3358 );
xor ( n3360 , n1760 , n1761 );
xor ( n3361 , n3360 , n2845 );
buf ( n3362 , n3361 );
xor ( n3363 , n1763 , n1764 );
xor ( n3364 , n3363 , n2842 );
buf ( n3365 , n3364 );
xor ( n3366 , n3362 , n3365 );
xor ( n3367 , n3359 , n3366 );
xor ( n3368 , n1766 , n1767 );
xor ( n3369 , n3368 , n2839 );
buf ( n3370 , n3369 );
xor ( n3371 , n1769 , n1770 );
xor ( n3372 , n3371 , n2836 );
buf ( n3373 , n3372 );
xor ( n3374 , n3370 , n3373 );
xor ( n3375 , n1772 , n1773 );
xor ( n3376 , n3375 , n2833 );
buf ( n3377 , n3376 );
xor ( n3378 , n1775 , n1776 );
xor ( n3379 , n3378 , n2830 );
buf ( n3380 , n3379 );
xor ( n3381 , n3377 , n3380 );
xor ( n3382 , n3374 , n3381 );
xor ( n3383 , n3367 , n3382 );
xor ( n3384 , n3352 , n3383 );
xor ( n3385 , n1778 , n1779 );
xor ( n3386 , n3385 , n2827 );
buf ( n3387 , n3386 );
xor ( n3388 , n1781 , n1782 );
xor ( n3389 , n3388 , n2824 );
buf ( n3390 , n3389 );
xor ( n3391 , n3387 , n3390 );
xor ( n3392 , n1784 , n1785 );
xor ( n3393 , n3392 , n2821 );
buf ( n3394 , n3393 );
xor ( n3395 , n1787 , n1788 );
xor ( n3396 , n3395 , n2818 );
buf ( n3397 , n3396 );
xor ( n3398 , n3394 , n3397 );
xor ( n3399 , n3391 , n3398 );
xor ( n3400 , n1790 , n1791 );
xor ( n3401 , n3400 , n2815 );
buf ( n3402 , n3401 );
xor ( n3403 , n1793 , n1794 );
xor ( n3404 , n3403 , n2812 );
buf ( n3405 , n3404 );
xor ( n3406 , n3402 , n3405 );
xor ( n3407 , n1796 , n1797 );
xor ( n3408 , n3407 , n2809 );
buf ( n3409 , n3408 );
xor ( n3410 , n1799 , n1800 );
xor ( n3411 , n3410 , n2806 );
buf ( n3412 , n3411 );
xor ( n3413 , n3409 , n3412 );
xor ( n3414 , n3406 , n3413 );
xor ( n3415 , n3399 , n3414 );
xor ( n3416 , n1802 , n1803 );
xor ( n3417 , n3416 , n2803 );
buf ( n3418 , n3417 );
xor ( n3419 , n1805 , n1806 );
xor ( n3420 , n3419 , n2800 );
buf ( n3421 , n3420 );
xor ( n3422 , n3418 , n3421 );
xor ( n3423 , n1808 , n1809 );
xor ( n3424 , n3423 , n2797 );
buf ( n3425 , n3424 );
xor ( n3426 , n1811 , n1812 );
xor ( n3427 , n3426 , n2794 );
buf ( n3428 , n3427 );
xor ( n3429 , n3425 , n3428 );
xor ( n3430 , n3422 , n3429 );
xor ( n3431 , n1814 , n1815 );
xor ( n3432 , n3431 , n2791 );
buf ( n3433 , n3432 );
xor ( n3434 , n1817 , n1818 );
xor ( n3435 , n3434 , n2788 );
buf ( n3436 , n3435 );
xor ( n3437 , n3433 , n3436 );
xor ( n3438 , n1820 , n1821 );
xor ( n3439 , n3438 , n2785 );
buf ( n3440 , n3439 );
xor ( n3441 , n1823 , n1824 );
xor ( n3442 , n3441 , n2782 );
buf ( n3443 , n3442 );
xor ( n3444 , n3440 , n3443 );
xor ( n3445 , n3437 , n3444 );
xor ( n3446 , n3430 , n3445 );
xor ( n3447 , n3415 , n3446 );
xor ( n3448 , n3384 , n3447 );
xor ( n3449 , n1826 , n1827 );
xor ( n3450 , n3449 , n2779 );
buf ( n3451 , n3450 );
xor ( n3452 , n1829 , n1830 );
xor ( n3453 , n3452 , n2776 );
buf ( n3454 , n3453 );
xor ( n3455 , n3451 , n3454 );
xor ( n3456 , n1832 , n1833 );
xor ( n3457 , n3456 , n2773 );
buf ( n3458 , n3457 );
xor ( n3459 , n1835 , n1836 );
xor ( n3460 , n3459 , n2770 );
buf ( n3461 , n3460 );
xor ( n3462 , n3458 , n3461 );
xor ( n3463 , n3455 , n3462 );
xor ( n3464 , n1838 , n1839 );
xor ( n3465 , n3464 , n2767 );
buf ( n3466 , n3465 );
xor ( n3467 , n1841 , n1842 );
xor ( n3468 , n3467 , n2764 );
buf ( n3469 , n3468 );
xor ( n3470 , n3466 , n3469 );
xor ( n3471 , n1844 , n1845 );
xor ( n3472 , n3471 , n2761 );
buf ( n3473 , n3472 );
xor ( n3474 , n1847 , n1848 );
xor ( n3475 , n3474 , n2758 );
buf ( n3476 , n3475 );
xor ( n3477 , n3473 , n3476 );
xor ( n3478 , n3470 , n3477 );
xor ( n3479 , n3463 , n3478 );
xor ( n3480 , n1850 , n1851 );
xor ( n3481 , n3480 , n2755 );
buf ( n3482 , n3481 );
xor ( n3483 , n1853 , n1854 );
xor ( n3484 , n3483 , n2752 );
buf ( n3485 , n3484 );
xor ( n3486 , n3482 , n3485 );
xor ( n3487 , n1856 , n1857 );
xor ( n3488 , n3487 , n2749 );
buf ( n3489 , n3488 );
xor ( n3490 , n1859 , n1860 );
xor ( n3491 , n3490 , n2746 );
buf ( n3492 , n3491 );
xor ( n3493 , n3489 , n3492 );
xor ( n3494 , n3486 , n3493 );
xor ( n3495 , n1862 , n1863 );
xor ( n3496 , n3495 , n2743 );
buf ( n3497 , n3496 );
xor ( n3498 , n1865 , n1866 );
xor ( n3499 , n3498 , n2740 );
buf ( n3500 , n3499 );
xor ( n3501 , n3497 , n3500 );
xor ( n3502 , n1868 , n1869 );
xor ( n3503 , n3502 , n2737 );
buf ( n3504 , n3503 );
xor ( n3505 , n1871 , n1872 );
xor ( n3506 , n3505 , n2734 );
buf ( n3507 , n3506 );
xor ( n3508 , n3504 , n3507 );
xor ( n3509 , n3501 , n3508 );
xor ( n3510 , n3494 , n3509 );
xor ( n3511 , n3479 , n3510 );
xor ( n3512 , n1874 , n1875 );
xor ( n3513 , n3512 , n2731 );
buf ( n3514 , n3513 );
xor ( n3515 , n1877 , n1878 );
xor ( n3516 , n3515 , n2728 );
buf ( n3517 , n3516 );
xor ( n3518 , n3514 , n3517 );
xor ( n3519 , n1880 , n1881 );
xor ( n3520 , n3519 , n2725 );
buf ( n3521 , n3520 );
xor ( n3522 , n1883 , n1884 );
xor ( n3523 , n3522 , n2722 );
buf ( n3524 , n3523 );
xor ( n3525 , n3521 , n3524 );
xor ( n3526 , n3518 , n3525 );
xor ( n3527 , n1886 , n1887 );
xor ( n3528 , n3527 , n2719 );
buf ( n3529 , n3528 );
xor ( n3530 , n1889 , n1890 );
xor ( n3531 , n3530 , n2716 );
buf ( n3532 , n3531 );
xor ( n3533 , n3529 , n3532 );
xor ( n3534 , n1892 , n1893 );
xor ( n3535 , n3534 , n2713 );
buf ( n3536 , n3535 );
xor ( n3537 , n1895 , n1896 );
xor ( n3538 , n3537 , n2710 );
buf ( n3539 , n3538 );
xor ( n3540 , n3536 , n3539 );
xor ( n3541 , n3533 , n3540 );
xor ( n3542 , n3526 , n3541 );
xor ( n3543 , n1898 , n1899 );
xor ( n3544 , n3543 , n2707 );
buf ( n3545 , n3544 );
xor ( n3546 , n1901 , n1902 );
xor ( n3547 , n3546 , n2704 );
buf ( n3548 , n3547 );
xor ( n3549 , n3545 , n3548 );
xor ( n3550 , n1904 , n1905 );
xor ( n3551 , n3550 , n2701 );
buf ( n3552 , n3551 );
xor ( n3553 , n1907 , n1908 );
xor ( n3554 , n3553 , n2698 );
buf ( n3555 , n3554 );
xor ( n3556 , n3552 , n3555 );
xor ( n3557 , n3549 , n3556 );
xor ( n3558 , n1910 , n1911 );
xor ( n3559 , n3558 , n2695 );
buf ( n3560 , n3559 );
xor ( n3561 , n1913 , n1914 );
xor ( n3562 , n3561 , n2692 );
buf ( n3563 , n3562 );
xor ( n3564 , n3560 , n3563 );
xor ( n3565 , n1916 , n1917 );
xor ( n3566 , n3565 , n2689 );
buf ( n3567 , n3566 );
xor ( n3568 , n1919 , n1920 );
xor ( n3569 , n3568 , n2686 );
buf ( n3570 , n3569 );
xor ( n3571 , n3567 , n3570 );
xor ( n3572 , n3564 , n3571 );
xor ( n3573 , n3557 , n3572 );
xor ( n3574 , n3542 , n3573 );
xor ( n3575 , n3511 , n3574 );
xor ( n3576 , n3448 , n3575 );
xor ( n3577 , n3321 , n3576 );
xor ( n3578 , n1922 , n1923 );
xor ( n3579 , n3578 , n2683 );
buf ( n3580 , n3579 );
xor ( n3581 , n1925 , n1926 );
xor ( n3582 , n3581 , n2680 );
buf ( n3583 , n3582 );
xor ( n3584 , n3580 , n3583 );
xor ( n3585 , n1928 , n1929 );
xor ( n3586 , n3585 , n2677 );
buf ( n3587 , n3586 );
xor ( n3588 , n1931 , n1932 );
xor ( n3589 , n3588 , n2674 );
buf ( n3590 , n3589 );
xor ( n3591 , n3587 , n3590 );
xor ( n3592 , n3584 , n3591 );
xor ( n3593 , n1934 , n1935 );
xor ( n3594 , n3593 , n2671 );
buf ( n3595 , n3594 );
xor ( n3596 , n1937 , n1938 );
xor ( n3597 , n3596 , n2668 );
buf ( n3598 , n3597 );
xor ( n3599 , n3595 , n3598 );
xor ( n3600 , n1940 , n1941 );
xor ( n3601 , n3600 , n2665 );
buf ( n3602 , n3601 );
xor ( n3603 , n1943 , n1944 );
xor ( n3604 , n3603 , n2662 );
buf ( n3605 , n3604 );
xor ( n3606 , n3602 , n3605 );
xor ( n3607 , n3599 , n3606 );
xor ( n3608 , n3592 , n3607 );
xor ( n3609 , n1946 , n1947 );
xor ( n3610 , n3609 , n2659 );
buf ( n3611 , n3610 );
xor ( n3612 , n1949 , n1950 );
xor ( n3613 , n3612 , n2656 );
buf ( n3614 , n3613 );
xor ( n3615 , n3611 , n3614 );
xor ( n3616 , n1952 , n1953 );
xor ( n3617 , n3616 , n2653 );
buf ( n3618 , n3617 );
xor ( n3619 , n1955 , n1956 );
xor ( n3620 , n3619 , n2650 );
buf ( n3621 , n3620 );
xor ( n3622 , n3618 , n3621 );
xor ( n3623 , n3615 , n3622 );
xor ( n3624 , n1958 , n1959 );
xor ( n3625 , n3624 , n2647 );
buf ( n3626 , n3625 );
xor ( n3627 , n1961 , n1962 );
xor ( n3628 , n3627 , n2644 );
buf ( n3629 , n3628 );
xor ( n3630 , n3626 , n3629 );
xor ( n3631 , n1964 , n1965 );
xor ( n3632 , n3631 , n2641 );
buf ( n3633 , n3632 );
xor ( n3634 , n1967 , n1968 );
xor ( n3635 , n3634 , n2638 );
buf ( n3636 , n3635 );
xor ( n3637 , n3633 , n3636 );
xor ( n3638 , n3630 , n3637 );
xor ( n3639 , n3623 , n3638 );
xor ( n3640 , n3608 , n3639 );
xor ( n3641 , n1970 , n1971 );
xor ( n3642 , n3641 , n2635 );
buf ( n3643 , n3642 );
xor ( n3644 , n1973 , n1974 );
xor ( n3645 , n3644 , n2632 );
buf ( n3646 , n3645 );
xor ( n3647 , n3643 , n3646 );
xor ( n3648 , n1976 , n1977 );
xor ( n3649 , n3648 , n2629 );
buf ( n3650 , n3649 );
xor ( n3651 , n1979 , n1980 );
xor ( n3652 , n3651 , n2626 );
buf ( n3653 , n3652 );
xor ( n3654 , n3650 , n3653 );
xor ( n3655 , n3647 , n3654 );
xor ( n3656 , n1982 , n1983 );
xor ( n3657 , n3656 , n2623 );
buf ( n3658 , n3657 );
xor ( n3659 , n1985 , n1986 );
xor ( n3660 , n3659 , n2620 );
buf ( n3661 , n3660 );
xor ( n3662 , n3658 , n3661 );
xor ( n3663 , n1988 , n1989 );
xor ( n3664 , n3663 , n2617 );
buf ( n3665 , n3664 );
xor ( n3666 , n1991 , n1992 );
xor ( n3667 , n3666 , n2614 );
buf ( n3668 , n3667 );
xor ( n3669 , n3665 , n3668 );
xor ( n3670 , n3662 , n3669 );
xor ( n3671 , n3655 , n3670 );
xor ( n3672 , n1994 , n1995 );
xor ( n3673 , n3672 , n2611 );
buf ( n3674 , n3673 );
xor ( n3675 , n1997 , n1998 );
xor ( n3676 , n3675 , n2608 );
buf ( n3677 , n3676 );
xor ( n3678 , n3674 , n3677 );
xor ( n3679 , n2000 , n2001 );
xor ( n3680 , n3679 , n2605 );
buf ( n3681 , n3680 );
xor ( n3682 , n2003 , n2004 );
xor ( n3683 , n3682 , n2602 );
buf ( n3684 , n3683 );
xor ( n3685 , n3681 , n3684 );
xor ( n3686 , n3678 , n3685 );
xor ( n3687 , n2006 , n2007 );
xor ( n3688 , n3687 , n2599 );
buf ( n3689 , n3688 );
xor ( n3690 , n2009 , n2010 );
xor ( n3691 , n3690 , n2596 );
buf ( n3692 , n3691 );
xor ( n3693 , n3689 , n3692 );
xor ( n3694 , n2012 , n2013 );
xor ( n3695 , n3694 , n2593 );
buf ( n3696 , n3695 );
xor ( n3697 , n2015 , n2016 );
xor ( n3698 , n3697 , n2590 );
buf ( n3699 , n3698 );
xor ( n3700 , n3696 , n3699 );
xor ( n3701 , n3693 , n3700 );
xor ( n3702 , n3686 , n3701 );
xor ( n3703 , n3671 , n3702 );
xor ( n3704 , n3640 , n3703 );
xor ( n3705 , n2018 , n2019 );
xor ( n3706 , n3705 , n2587 );
buf ( n3707 , n3706 );
xor ( n3708 , n2021 , n2022 );
xor ( n3709 , n3708 , n2584 );
buf ( n3710 , n3709 );
xor ( n3711 , n3707 , n3710 );
xor ( n3712 , n2024 , n2025 );
xor ( n3713 , n3712 , n2581 );
buf ( n3714 , n3713 );
xor ( n3715 , n2027 , n2028 );
xor ( n3716 , n3715 , n2578 );
buf ( n3717 , n3716 );
xor ( n3718 , n3714 , n3717 );
xor ( n3719 , n3711 , n3718 );
xor ( n3720 , n2030 , n2031 );
xor ( n3721 , n3720 , n2575 );
buf ( n3722 , n3721 );
xor ( n3723 , n2033 , n2034 );
xor ( n3724 , n3723 , n2572 );
buf ( n3725 , n3724 );
xor ( n3726 , n3722 , n3725 );
xor ( n3727 , n2036 , n2037 );
xor ( n3728 , n3727 , n2569 );
buf ( n3729 , n3728 );
xor ( n3730 , n2039 , n2040 );
xor ( n3731 , n3730 , n2566 );
buf ( n3732 , n3731 );
xor ( n3733 , n3729 , n3732 );
xor ( n3734 , n3726 , n3733 );
xor ( n3735 , n3719 , n3734 );
xor ( n3736 , n2042 , n2043 );
xor ( n3737 , n3736 , n2563 );
buf ( n3738 , n3737 );
xor ( n3739 , n2045 , n2046 );
xor ( n3740 , n3739 , n2560 );
buf ( n3741 , n3740 );
xor ( n3742 , n3738 , n3741 );
xor ( n3743 , n2048 , n2049 );
xor ( n3744 , n3743 , n2557 );
buf ( n3745 , n3744 );
xor ( n3746 , n2051 , n2052 );
xor ( n3747 , n3746 , n2554 );
buf ( n3748 , n3747 );
xor ( n3749 , n3745 , n3748 );
xor ( n3750 , n3742 , n3749 );
xor ( n3751 , n2054 , n2055 );
xor ( n3752 , n3751 , n2551 );
buf ( n3753 , n3752 );
xor ( n3754 , n2057 , n2058 );
xor ( n3755 , n3754 , n2548 );
buf ( n3756 , n3755 );
xor ( n3757 , n3753 , n3756 );
xor ( n3758 , n2060 , n2061 );
xor ( n3759 , n3758 , n2545 );
buf ( n3760 , n3759 );
xor ( n3761 , n2063 , n2064 );
xor ( n3762 , n3761 , n2542 );
buf ( n3763 , n3762 );
xor ( n3764 , n3760 , n3763 );
xor ( n3765 , n3757 , n3764 );
xor ( n3766 , n3750 , n3765 );
xor ( n3767 , n3735 , n3766 );
xor ( n3768 , n2066 , n2067 );
xor ( n3769 , n3768 , n2539 );
buf ( n3770 , n3769 );
xor ( n3771 , n2069 , n2070 );
xor ( n3772 , n3771 , n2536 );
buf ( n3773 , n3772 );
xor ( n3774 , n3770 , n3773 );
xor ( n3775 , n2072 , n2073 );
xor ( n3776 , n3775 , n2533 );
buf ( n3777 , n3776 );
xor ( n3778 , n2075 , n2076 );
xor ( n3779 , n3778 , n2530 );
buf ( n3780 , n3779 );
xor ( n3781 , n3777 , n3780 );
xor ( n3782 , n3774 , n3781 );
xor ( n3783 , n2078 , n2079 );
xor ( n3784 , n3783 , n2527 );
buf ( n3785 , n3784 );
xor ( n3786 , n2081 , n2082 );
xor ( n3787 , n3786 , n2524 );
buf ( n3788 , n3787 );
xor ( n3789 , n3785 , n3788 );
xor ( n3790 , n2084 , n2085 );
xor ( n3791 , n3790 , n2521 );
buf ( n3792 , n3791 );
xor ( n3793 , n2087 , n2088 );
xor ( n3794 , n3793 , n2518 );
buf ( n3795 , n3794 );
xor ( n3796 , n3792 , n3795 );
xor ( n3797 , n3789 , n3796 );
xor ( n3798 , n3782 , n3797 );
xor ( n3799 , n2090 , n2091 );
xor ( n3800 , n3799 , n2515 );
buf ( n3801 , n3800 );
xor ( n3802 , n2093 , n2094 );
xor ( n3803 , n3802 , n2512 );
buf ( n3804 , n3803 );
xor ( n3805 , n3801 , n3804 );
xor ( n3806 , n2096 , n2097 );
xor ( n3807 , n3806 , n2509 );
buf ( n3808 , n3807 );
xor ( n3809 , n2099 , n2100 );
xor ( n3810 , n3809 , n2506 );
buf ( n3811 , n3810 );
xor ( n3812 , n3808 , n3811 );
xor ( n3813 , n3805 , n3812 );
xor ( n3814 , n2102 , n2103 );
xor ( n3815 , n3814 , n2503 );
buf ( n3816 , n3815 );
xor ( n3817 , n2105 , n2106 );
xor ( n3818 , n3817 , n2500 );
buf ( n3819 , n3818 );
xor ( n3820 , n3816 , n3819 );
xor ( n3821 , n2108 , n2109 );
xor ( n3822 , n3821 , n2497 );
buf ( n3823 , n3822 );
xor ( n3824 , n2111 , n2112 );
xor ( n3825 , n3824 , n2494 );
buf ( n3826 , n3825 );
xor ( n3827 , n3823 , n3826 );
xor ( n3828 , n3820 , n3827 );
xor ( n3829 , n3813 , n3828 );
xor ( n3830 , n3798 , n3829 );
xor ( n3831 , n3767 , n3830 );
xor ( n3832 , n3704 , n3831 );
xor ( n3833 , n2114 , n2115 );
xor ( n3834 , n3833 , n2491 );
buf ( n3835 , n3834 );
xor ( n3836 , n2117 , n2118 );
xor ( n3837 , n3836 , n2488 );
buf ( n3838 , n3837 );
xor ( n3839 , n3835 , n3838 );
xor ( n3840 , n2120 , n2121 );
xor ( n3841 , n3840 , n2485 );
buf ( n3842 , n3841 );
xor ( n3843 , n2123 , n2124 );
xor ( n3844 , n3843 , n2482 );
buf ( n3845 , n3844 );
xor ( n3846 , n3842 , n3845 );
xor ( n3847 , n3839 , n3846 );
xor ( n3848 , n2126 , n2127 );
xor ( n3849 , n3848 , n2479 );
buf ( n3850 , n3849 );
xor ( n3851 , n2129 , n2130 );
xor ( n3852 , n3851 , n2476 );
buf ( n3853 , n3852 );
xor ( n3854 , n3850 , n3853 );
xor ( n3855 , n2132 , n2133 );
xor ( n3856 , n3855 , n2473 );
buf ( n3857 , n3856 );
xor ( n3858 , n2135 , n2136 );
xor ( n3859 , n3858 , n2470 );
buf ( n3860 , n3859 );
xor ( n3861 , n3857 , n3860 );
xor ( n3862 , n3854 , n3861 );
xor ( n3863 , n3847 , n3862 );
xor ( n3864 , n2138 , n2139 );
xor ( n3865 , n3864 , n2467 );
buf ( n3866 , n3865 );
xor ( n3867 , n2141 , n2142 );
xor ( n3868 , n3867 , n2464 );
buf ( n3869 , n3868 );
xor ( n3870 , n3866 , n3869 );
xor ( n3871 , n2144 , n2145 );
xor ( n3872 , n3871 , n2461 );
buf ( n3873 , n3872 );
xor ( n3874 , n2147 , n2148 );
xor ( n3875 , n3874 , n2458 );
buf ( n3876 , n3875 );
xor ( n3877 , n3873 , n3876 );
xor ( n3878 , n3870 , n3877 );
xor ( n3879 , n2150 , n2151 );
xor ( n3880 , n3879 , n2455 );
buf ( n3881 , n3880 );
xor ( n3882 , n2153 , n2154 );
xor ( n3883 , n3882 , n2452 );
buf ( n3884 , n3883 );
xor ( n3885 , n3881 , n3884 );
xor ( n3886 , n2156 , n2157 );
xor ( n3887 , n3886 , n2449 );
buf ( n3888 , n3887 );
xor ( n3889 , n2159 , n2160 );
xor ( n3890 , n3889 , n2446 );
buf ( n3891 , n3890 );
xor ( n3892 , n3888 , n3891 );
xor ( n3893 , n3885 , n3892 );
xor ( n3894 , n3878 , n3893 );
xor ( n3895 , n3863 , n3894 );
xor ( n3896 , n2162 , n2163 );
xor ( n3897 , n3896 , n2443 );
buf ( n3898 , n3897 );
xor ( n3899 , n2165 , n2166 );
xor ( n3900 , n3899 , n2440 );
buf ( n3901 , n3900 );
xor ( n3902 , n3898 , n3901 );
xor ( n3903 , n2168 , n2169 );
xor ( n3904 , n3903 , n2437 );
buf ( n3905 , n3904 );
xor ( n3906 , n2171 , n2172 );
xor ( n3907 , n3906 , n2434 );
buf ( n3908 , n3907 );
xor ( n3909 , n3905 , n3908 );
xor ( n3910 , n3902 , n3909 );
xor ( n3911 , n2174 , n2175 );
xor ( n3912 , n3911 , n2431 );
buf ( n3913 , n3912 );
xor ( n3914 , n2177 , n2178 );
xor ( n3915 , n3914 , n2428 );
buf ( n3916 , n3915 );
xor ( n3917 , n3913 , n3916 );
xor ( n3918 , n2180 , n2181 );
xor ( n3919 , n3918 , n2425 );
buf ( n3920 , n3919 );
xor ( n3921 , n2183 , n2184 );
xor ( n3922 , n3921 , n2422 );
buf ( n3923 , n3922 );
xor ( n3924 , n3920 , n3923 );
xor ( n3925 , n3917 , n3924 );
xor ( n3926 , n3910 , n3925 );
xor ( n3927 , n2186 , n2187 );
xor ( n3928 , n3927 , n2419 );
buf ( n3929 , n3928 );
xor ( n3930 , n2189 , n2190 );
xor ( n3931 , n3930 , n2416 );
buf ( n3932 , n3931 );
xor ( n3933 , n3929 , n3932 );
xor ( n3934 , n2192 , n2193 );
xor ( n3935 , n3934 , n2413 );
buf ( n3936 , n3935 );
xor ( n3937 , n2195 , n2196 );
xor ( n3938 , n3937 , n2410 );
buf ( n3939 , n3938 );
xor ( n3940 , n3936 , n3939 );
xor ( n3941 , n3933 , n3940 );
xor ( n3942 , n2198 , n2199 );
xor ( n3943 , n3942 , n2407 );
buf ( n3944 , n3943 );
xor ( n3945 , n2201 , n2202 );
xor ( n3946 , n3945 , n2404 );
buf ( n3947 , n3946 );
xor ( n3948 , n3944 , n3947 );
xor ( n3949 , n2204 , n2205 );
xor ( n3950 , n3949 , n2401 );
buf ( n3951 , n3950 );
xor ( n3952 , n2207 , n2208 );
xor ( n3953 , n3952 , n2398 );
buf ( n3954 , n3953 );
xor ( n3955 , n3951 , n3954 );
xor ( n3956 , n3948 , n3955 );
xor ( n3957 , n3941 , n3956 );
xor ( n3958 , n3926 , n3957 );
xor ( n3959 , n3895 , n3958 );
xor ( n3960 , n2210 , n2211 );
xor ( n3961 , n3960 , n2395 );
buf ( n3962 , n3961 );
xor ( n3963 , n2213 , n2214 );
xor ( n3964 , n3963 , n2392 );
buf ( n3965 , n3964 );
xor ( n3966 , n3962 , n3965 );
xor ( n3967 , n2216 , n2217 );
xor ( n3968 , n3967 , n2389 );
buf ( n3969 , n3968 );
xor ( n3970 , n2219 , n2220 );
xor ( n3971 , n3970 , n2386 );
buf ( n3972 , n3971 );
xor ( n3973 , n3969 , n3972 );
xor ( n3974 , n3966 , n3973 );
xor ( n3975 , n2222 , n2223 );
xor ( n3976 , n3975 , n2383 );
buf ( n3977 , n3976 );
xor ( n3978 , n2225 , n2226 );
xor ( n3979 , n3978 , n2380 );
buf ( n3980 , n3979 );
xor ( n3981 , n3977 , n3980 );
xor ( n3982 , n2228 , n2229 );
xor ( n3983 , n3982 , n2377 );
buf ( n3984 , n3983 );
xor ( n3985 , n2231 , n2232 );
xor ( n3986 , n3985 , n2374 );
buf ( n3987 , n3986 );
xor ( n3988 , n3984 , n3987 );
xor ( n3989 , n3981 , n3988 );
xor ( n3990 , n3974 , n3989 );
xor ( n3991 , n2234 , n2235 );
xor ( n3992 , n3991 , n2371 );
buf ( n3993 , n3992 );
xor ( n3994 , n2237 , n2238 );
xor ( n3995 , n3994 , n2368 );
buf ( n3996 , n3995 );
xor ( n3997 , n3993 , n3996 );
xor ( n3998 , n2240 , n2241 );
xor ( n3999 , n3998 , n2365 );
buf ( n4000 , n3999 );
xor ( n4001 , n2243 , n2244 );
xor ( n4002 , n4001 , n2362 );
buf ( n4003 , n4002 );
xor ( n4004 , n4000 , n4003 );
xor ( n4005 , n3997 , n4004 );
xor ( n4006 , n2246 , n2247 );
xor ( n4007 , n4006 , n2359 );
buf ( n4008 , n4007 );
xor ( n4009 , n2249 , n2250 );
xor ( n4010 , n4009 , n2356 );
buf ( n4011 , n4010 );
xor ( n4012 , n4008 , n4011 );
xor ( n4013 , n2252 , n2253 );
xor ( n4014 , n4013 , n2353 );
buf ( n4015 , n4014 );
xor ( n4016 , n2255 , n2256 );
xor ( n4017 , n4016 , n2350 );
buf ( n4018 , n4017 );
xor ( n4019 , n4015 , n4018 );
xor ( n4020 , n4012 , n4019 );
xor ( n4021 , n4005 , n4020 );
xor ( n4022 , n3990 , n4021 );
xor ( n4023 , n2258 , n2259 );
xor ( n4024 , n4023 , n2347 );
buf ( n4025 , n4024 );
xor ( n4026 , n2261 , n2262 );
xor ( n4027 , n4026 , n2344 );
buf ( n4028 , n4027 );
xor ( n4029 , n4025 , n4028 );
xor ( n4030 , n2264 , n2265 );
xor ( n4031 , n4030 , n2341 );
buf ( n4032 , n4031 );
xor ( n4033 , n2267 , n2268 );
xor ( n4034 , n4033 , n2338 );
buf ( n4035 , n4034 );
xor ( n4036 , n4032 , n4035 );
xor ( n4037 , n4029 , n4036 );
xor ( n4038 , n2270 , n2271 );
xor ( n4039 , n4038 , n2335 );
buf ( n4040 , n4039 );
xor ( n4041 , n2273 , n2274 );
xor ( n4042 , n4041 , n2332 );
buf ( n4043 , n4042 );
xor ( n4044 , n4040 , n4043 );
xor ( n4045 , n2276 , n2277 );
xor ( n4046 , n4045 , n2329 );
buf ( n4047 , n4046 );
xor ( n4048 , n2279 , n2280 );
xor ( n4049 , n4048 , n2326 );
buf ( n4050 , n4049 );
xor ( n4051 , n4047 , n4050 );
xor ( n4052 , n4044 , n4051 );
xor ( n4053 , n4037 , n4052 );
xor ( n4054 , n2282 , n2283 );
xor ( n4055 , n4054 , n2323 );
buf ( n4056 , n4055 );
xor ( n4057 , n2285 , n2286 );
xor ( n4058 , n4057 , n2320 );
buf ( n4059 , n4058 );
xor ( n4060 , n4056 , n4059 );
xor ( n4061 , n2288 , n2289 );
xor ( n4062 , n4061 , n2317 );
buf ( n4063 , n4062 );
xor ( n4064 , n2291 , n2292 );
xor ( n4065 , n4064 , n2314 );
buf ( n4066 , n4065 );
xor ( n4067 , n4063 , n4066 );
xor ( n4068 , n4060 , n4067 );
xor ( n4069 , n2294 , n2295 );
xor ( n4070 , n4069 , n2311 );
buf ( n4071 , n4070 );
xor ( n4072 , n2297 , n2298 );
xor ( n4073 , n4072 , n2308 );
buf ( n4074 , n4073 );
xor ( n4075 , n4071 , n4074 );
xor ( n4076 , n2300 , n2301 );
xor ( n4077 , n4076 , n2305 );
buf ( n4078 , n4077 );
xor ( n4079 , n2303 , n2304 );
buf ( n4080 , n4079 );
xor ( n4081 , n4078 , n4080 );
xor ( n4082 , n4075 , n4081 );
xor ( n4083 , n4068 , n4082 );
xor ( n4084 , n4053 , n4083 );
xor ( n4085 , n4022 , n4084 );
xor ( n4086 , n3959 , n4085 );
xor ( n4087 , n3832 , n4086 );
xor ( n4088 , n3577 , n4087 );
buf ( n4089 , n4088 );
buf ( n4090 , n4089 );
endmodule

