//
// Conformal-LEC Version 15.20-d227 ( 10-Mar-2016) ( 64 bit executable)
//
module top ( n0 , n1 , n2 , n3 , n4 , n6 , n7 , n9 , n12 , n13 ,  n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 );
input n0 , n1 , n2 , n3 , n4 , n6 , n7 , n9 , n12 , n13 ,  n15 ;
output n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;

wire n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , 
     n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , 
     n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , 
     n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , 
     n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , 
     n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , 
     n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , 
     n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , 
     n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , 
     n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , 
     n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , 
     n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , 
     n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , 
     n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , 
     n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , 
     n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , 
     n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , 
     n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , 
     n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , 
     n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , 
     n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , 
     n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , 
     n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , 
     n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , 
     n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , 
     n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , 
     n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , 
     n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , 
     n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , 
     n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , 
     n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , 
     n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , 
     n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , 
     n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , 
     n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , 
     n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , 
     n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , 
     n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , 
     n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , 
     n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , 
     n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , 
     n473 , n474 , n475 , n476 ;
buf ( n29 , n428 );
buf ( n23 , n431 );
buf ( n31 , n434 );
buf ( n19 , n437 );
buf ( n16 , n440 );
buf ( n18 , n443 );
buf ( n17 , n446 );
buf ( n25 , n449 );
buf ( n22 , n452 );
buf ( n27 , n455 );
buf ( n28 , n458 );
buf ( n30 , n462 );
buf ( n20 , n466 );
buf ( n26 , n470 );
buf ( n21 , n473 );
buf ( n24 , n476 );
buf ( n66 , n13 );
buf ( n67 , n9 );
buf ( n68 , n3 );
buf ( n69 , n15 );
buf ( n70 , n7 );
buf ( n71 , n2 );
buf ( n72 , n1 );
buf ( n73 , n6 );
buf ( n74 , n4 );
buf ( n75 , n0 );
buf ( n76 , n12 );
buf ( n77 , n67 );
buf ( n78 , n70 );
and ( n79 , n77 , n78 );
buf ( n80 , n69 );
not ( n81 , n80 );
not ( n82 , n78 );
and ( n83 , n82 , n80 );
nor ( n84 , n81 , n83 );
buf ( n85 , n68 );
buf ( n86 , n71 );
and ( n87 , n85 , n86 );
and ( n88 , n84 , n87 );
buf ( n89 , n67 );
buf ( n90 , n72 );
and ( n91 , n89 , n90 );
and ( n92 , n87 , n91 );
and ( n93 , n84 , n91 );
or ( n94 , n88 , n92 , n93 );
not ( n95 , n85 );
and ( n96 , n82 , n85 );
nor ( n97 , n95 , n96 );
and ( n98 , n94 , n97 );
and ( n99 , n89 , n86 );
and ( n100 , n97 , n99 );
and ( n101 , n94 , n99 );
or ( n102 , n98 , n100 , n101 );
not ( n103 , n89 );
and ( n104 , n82 , n89 );
nor ( n105 , n103 , n104 );
and ( n106 , n102 , n105 );
not ( n107 , n77 );
and ( n108 , n107 , n86 );
not ( n109 , n86 );
nor ( n110 , n108 , n109 );
and ( n111 , n105 , n110 );
and ( n112 , n102 , n110 );
or ( n113 , n106 , n111 , n112 );
and ( n114 , n79 , n113 );
xor ( n115 , n79 , n113 );
xor ( n116 , n102 , n105 );
xor ( n117 , n116 , n110 );
buf ( n118 , n69 );
not ( n119 , n118 );
and ( n120 , n82 , n118 );
nor ( n121 , n119 , n120 );
and ( n122 , n80 , n86 );
and ( n123 , n121 , n122 );
buf ( n124 , n74 );
and ( n125 , n107 , n124 );
not ( n126 , n124 );
nor ( n127 , n125 , n126 );
and ( n128 , n122 , n127 );
and ( n129 , n121 , n127 );
or ( n130 , n123 , n128 , n129 );
and ( n131 , n80 , n90 );
buf ( n132 , n73 );
and ( n133 , n85 , n132 );
and ( n134 , n131 , n133 );
and ( n135 , n89 , n124 );
and ( n136 , n133 , n135 );
and ( n137 , n131 , n135 );
or ( n138 , n134 , n136 , n137 );
and ( n139 , n85 , n90 );
and ( n140 , n138 , n139 );
and ( n141 , n89 , n132 );
and ( n142 , n139 , n141 );
and ( n143 , n138 , n141 );
or ( n144 , n140 , n142 , n143 );
and ( n145 , n130 , n144 );
xor ( n146 , n84 , n87 );
xor ( n147 , n146 , n91 );
and ( n148 , n144 , n147 );
and ( n149 , n130 , n147 );
or ( n150 , n145 , n148 , n149 );
and ( n151 , n107 , n90 );
not ( n152 , n90 );
nor ( n153 , n151 , n152 );
and ( n154 , n150 , n153 );
xor ( n155 , n94 , n97 );
xor ( n156 , n155 , n99 );
and ( n157 , n153 , n156 );
and ( n158 , n150 , n156 );
or ( n159 , n154 , n157 , n158 );
and ( n160 , n117 , n159 );
xor ( n161 , n117 , n159 );
xor ( n162 , n150 , n153 );
xor ( n163 , n162 , n156 );
and ( n164 , n80 , n132 );
and ( n165 , n85 , n124 );
and ( n166 , n164 , n165 );
buf ( n167 , n75 );
and ( n168 , n89 , n167 );
and ( n169 , n165 , n168 );
and ( n170 , n164 , n168 );
or ( n171 , n166 , n169 , n170 );
buf ( n172 , n86 );
and ( n173 , n118 , n90 );
and ( n174 , n172 , n173 );
and ( n175 , n171 , n174 );
xor ( n176 , n131 , n133 );
xor ( n177 , n176 , n135 );
and ( n178 , n174 , n177 );
and ( n179 , n171 , n177 );
or ( n180 , n175 , n178 , n179 );
xor ( n181 , n121 , n122 );
xor ( n182 , n181 , n127 );
and ( n183 , n180 , n182 );
xor ( n184 , n138 , n139 );
xor ( n185 , n184 , n141 );
and ( n186 , n182 , n185 );
and ( n187 , n180 , n185 );
or ( n188 , n183 , n186 , n187 );
and ( n189 , n107 , n132 );
not ( n190 , n132 );
nor ( n191 , n189 , n190 );
and ( n192 , n188 , n191 );
xor ( n193 , n130 , n144 );
xor ( n194 , n193 , n147 );
and ( n195 , n191 , n194 );
and ( n196 , n188 , n194 );
or ( n197 , n192 , n195 , n196 );
and ( n198 , n163 , n197 );
xor ( n199 , n163 , n197 );
xor ( n200 , n188 , n191 );
xor ( n201 , n200 , n194 );
buf ( n202 , n82 );
not ( n203 , n202 );
and ( n204 , n118 , n86 );
and ( n205 , n203 , n204 );
and ( n206 , n107 , n167 );
not ( n207 , n167 );
nor ( n208 , n206 , n207 );
and ( n209 , n204 , n208 );
and ( n210 , n203 , n208 );
or ( n211 , n205 , n209 , n210 );
and ( n212 , n80 , n124 );
and ( n213 , n85 , n167 );
and ( n214 , n212 , n213 );
buf ( n215 , n76 );
and ( n216 , n89 , n215 );
and ( n217 , n213 , n216 );
and ( n218 , n212 , n216 );
or ( n219 , n214 , n217 , n218 );
xor ( n220 , n164 , n165 );
xor ( n221 , n220 , n168 );
and ( n222 , n219 , n221 );
xor ( n223 , n172 , n173 );
and ( n224 , n221 , n223 );
and ( n225 , n219 , n223 );
or ( n226 , n222 , n224 , n225 );
xor ( n227 , n203 , n204 );
xor ( n228 , n227 , n208 );
and ( n229 , n226 , n228 );
xor ( n230 , n171 , n174 );
xor ( n231 , n230 , n177 );
and ( n232 , n228 , n231 );
and ( n233 , n226 , n231 );
or ( n234 , n229 , n232 , n233 );
and ( n235 , n211 , n234 );
xor ( n236 , n180 , n182 );
xor ( n237 , n236 , n185 );
and ( n238 , n234 , n237 );
and ( n239 , n211 , n237 );
or ( n240 , n235 , n238 , n239 );
and ( n241 , n201 , n240 );
xor ( n242 , n201 , n240 );
xor ( n243 , n211 , n234 );
xor ( n244 , n243 , n237 );
buf ( n245 , n90 );
and ( n246 , n118 , n132 );
and ( n247 , n245 , n246 );
buf ( n248 , n247 );
and ( n249 , n107 , n215 );
not ( n250 , n215 );
nor ( n251 , n249 , n250 );
and ( n252 , n248 , n251 );
buf ( n253 , n252 );
and ( n254 , n80 , n167 );
and ( n255 , n85 , n215 );
and ( n256 , n254 , n255 );
not ( n257 , n73 );
buf ( n258 , n257 );
and ( n259 , n89 , n258 );
and ( n260 , n255 , n259 );
and ( n261 , n254 , n259 );
or ( n262 , n256 , n260 , n261 );
buf ( n263 , n245 );
xor ( n264 , n263 , n246 );
and ( n265 , n262 , n264 );
xor ( n266 , n212 , n213 );
xor ( n267 , n266 , n216 );
and ( n268 , n264 , n267 );
and ( n269 , n262 , n267 );
or ( n270 , n265 , n268 , n269 );
buf ( n271 , n248 );
xor ( n272 , n271 , n251 );
and ( n273 , n270 , n272 );
xor ( n274 , n219 , n221 );
xor ( n275 , n274 , n223 );
and ( n276 , n272 , n275 );
and ( n277 , n270 , n275 );
or ( n278 , n273 , n276 , n277 );
and ( n279 , n253 , n278 );
xor ( n280 , n226 , n228 );
xor ( n281 , n280 , n231 );
and ( n282 , n278 , n281 );
and ( n283 , n253 , n281 );
or ( n284 , n279 , n282 , n283 );
and ( n285 , n244 , n284 );
xor ( n286 , n244 , n284 );
xor ( n287 , n253 , n278 );
xor ( n288 , n287 , n281 );
buf ( n289 , n66 );
not ( n290 , n289 );
and ( n291 , n82 , n289 );
nor ( n292 , n290 , n291 );
and ( n293 , n107 , n258 );
not ( n294 , n258 );
nor ( n295 , n293 , n294 );
and ( n296 , n292 , n295 );
and ( n297 , n80 , n215 );
and ( n298 , n85 , n258 );
and ( n299 , n297 , n298 );
and ( n300 , n118 , n124 );
and ( n301 , n299 , n300 );
xor ( n302 , n254 , n255 );
xor ( n303 , n302 , n259 );
and ( n304 , n300 , n303 );
and ( n305 , n299 , n303 );
or ( n306 , n301 , n304 , n305 );
xor ( n307 , n262 , n264 );
xor ( n308 , n307 , n267 );
and ( n309 , n306 , n308 );
xor ( n310 , n292 , n295 );
and ( n311 , n308 , n310 );
and ( n312 , n306 , n310 );
or ( n313 , n309 , n311 , n312 );
and ( n314 , n296 , n313 );
xor ( n315 , n270 , n272 );
xor ( n316 , n315 , n275 );
and ( n317 , n313 , n316 );
and ( n318 , n296 , n316 );
or ( n319 , n314 , n317 , n318 );
and ( n320 , n288 , n319 );
xor ( n321 , n288 , n319 );
xor ( n322 , n296 , n313 );
xor ( n323 , n322 , n316 );
and ( n324 , n289 , n86 );
buf ( n325 , n132 );
and ( n326 , n324 , n325 );
buf ( n327 , n326 );
buf ( n328 , n167 );
and ( n329 , n118 , n215 );
and ( n330 , n328 , n329 );
and ( n331 , n80 , n258 );
and ( n332 , n329 , n331 );
and ( n333 , n328 , n331 );
or ( n334 , n330 , n332 , n333 );
and ( n335 , n118 , n167 );
and ( n336 , n334 , n335 );
xor ( n337 , n297 , n298 );
and ( n338 , n335 , n337 );
and ( n339 , n334 , n337 );
or ( n340 , n336 , n338 , n339 );
buf ( n341 , n324 );
xor ( n342 , n341 , n325 );
and ( n343 , n340 , n342 );
xor ( n344 , n299 , n300 );
xor ( n345 , n344 , n303 );
and ( n346 , n342 , n345 );
and ( n347 , n340 , n345 );
or ( n348 , n343 , n346 , n347 );
and ( n349 , n327 , n348 );
xor ( n350 , n306 , n308 );
xor ( n351 , n350 , n310 );
and ( n352 , n348 , n351 );
and ( n353 , n327 , n351 );
or ( n354 , n349 , n352 , n353 );
and ( n355 , n323 , n354 );
xor ( n356 , n323 , n354 );
xor ( n357 , n327 , n348 );
xor ( n358 , n357 , n351 );
buf ( n359 , n215 );
and ( n360 , n118 , n258 );
and ( n361 , n359 , n360 );
buf ( n362 , n361 );
xor ( n363 , n328 , n329 );
xor ( n364 , n363 , n331 );
and ( n365 , n362 , n364 );
buf ( n366 , n365 );
buf ( n367 , n124 );
and ( n368 , n366 , n367 );
xor ( n369 , n334 , n335 );
xor ( n370 , n369 , n337 );
and ( n371 , n367 , n370 );
and ( n372 , n366 , n370 );
or ( n373 , n368 , n371 , n372 );
xor ( n374 , n340 , n342 );
xor ( n375 , n374 , n345 );
and ( n376 , n373 , n375 );
buf ( n377 , n376 );
and ( n378 , n358 , n377 );
xor ( n379 , n358 , n377 );
buf ( n380 , n373 );
xor ( n381 , n380 , n375 );
and ( n382 , n289 , n167 );
buf ( n383 , n258 );
and ( n384 , n382 , n383 );
buf ( n385 , n384 );
and ( n386 , n289 , n124 );
and ( n387 , n385 , n386 );
buf ( n388 , n359 );
xor ( n389 , n388 , n360 );
and ( n390 , n386 , n389 );
and ( n391 , n385 , n389 );
or ( n392 , n387 , n390 , n391 );
and ( n393 , n289 , n132 );
and ( n394 , n392 , n393 );
buf ( n395 , n362 );
xor ( n396 , n395 , n364 );
and ( n397 , n393 , n396 );
and ( n398 , n392 , n396 );
or ( n399 , n394 , n397 , n398 );
xor ( n400 , n367 , n366 );
xor ( n401 , n400 , n370 );
and ( n402 , n399 , n401 );
and ( n403 , n381 , n402 );
xor ( n404 , n381 , n402 );
and ( n405 , n289 , n90 );
xor ( n406 , n399 , n401 );
and ( n407 , n405 , n406 );
buf ( n408 , n407 );
and ( n409 , n404 , n408 );
or ( n410 , n403 , n409 );
and ( n411 , n379 , n410 );
or ( n412 , n378 , n411 );
and ( n413 , n356 , n412 );
or ( n414 , n355 , n413 );
and ( n415 , n321 , n414 );
or ( n416 , n320 , n415 );
and ( n417 , n286 , n416 );
or ( n418 , n285 , n417 );
and ( n419 , n242 , n418 );
or ( n420 , n241 , n419 );
and ( n421 , n199 , n420 );
or ( n422 , n198 , n421 );
and ( n423 , n161 , n422 );
or ( n424 , n160 , n423 );
and ( n425 , n115 , n424 );
or ( n426 , n114 , n425 );
buf ( n427 , n426 );
buf ( n428 , n427 );
xor ( n429 , n115 , n424 );
buf ( n430 , n429 );
buf ( n431 , n430 );
xor ( n432 , n161 , n422 );
buf ( n433 , n432 );
buf ( n434 , n433 );
xor ( n435 , n199 , n420 );
buf ( n436 , n435 );
buf ( n437 , n436 );
xor ( n438 , n242 , n418 );
buf ( n439 , n438 );
buf ( n440 , n439 );
xor ( n441 , n286 , n416 );
buf ( n442 , n441 );
buf ( n443 , n442 );
xor ( n444 , n321 , n414 );
buf ( n445 , n444 );
buf ( n446 , n445 );
xor ( n447 , n356 , n412 );
buf ( n448 , n447 );
buf ( n449 , n448 );
xor ( n450 , n379 , n410 );
buf ( n451 , n450 );
buf ( n452 , n451 );
xor ( n453 , n408 , n404 );
buf ( n454 , n453 );
buf ( n455 , n454 );
xor ( n456 , n405 , n406 );
buf ( n457 , n456 );
buf ( n458 , n457 );
xor ( n459 , n393 , n392 );
xor ( n460 , n459 , n396 );
buf ( n461 , n460 );
buf ( n462 , n461 );
xor ( n463 , n385 , n386 );
xor ( n464 , n463 , n389 );
buf ( n465 , n464 );
buf ( n466 , n465 );
buf ( n467 , n382 );
xor ( n468 , n467 , n383 );
buf ( n469 , n468 );
buf ( n470 , n469 );
and ( n471 , n289 , n215 );
buf ( n472 , n471 );
buf ( n473 , n472 );
and ( n474 , n289 , n258 );
buf ( n475 , n474 );
buf ( n476 , n475 );
endmodule

