//
// Conformal-LEC Version 15.20-d227 ( 10-Mar-2016) ( 64 bit executable)
//
module top ( n0 , n1 , n2 , n3 , n4 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 );
input n0 , n1 , n2 , n3 , n4 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 ;
output n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 ;

wire n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , 
     n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , 
     n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , 
     n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , 
     n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
     n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
     n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , 
     n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , 
     n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , 
     n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , 
     n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , 
     n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , 
     n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , 
     n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , 
     n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , 
     n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , 
     n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , 
     n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , 
     n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
     n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
     n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
     n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
     n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , 
     n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , 
     n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , 
     n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , 
     n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , 
     n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , 
     n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , 
     n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , 
     n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , 
     n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , 
     n437 , n438 , n439 , n440 , n441 ;
buf ( n53 , n382 );
buf ( n43 , n386 );
buf ( n58 , n390 );
buf ( n56 , n394 );
buf ( n52 , n398 );
buf ( n51 , n402 );
buf ( n44 , n406 );
buf ( n50 , n410 );
buf ( n45 , n414 );
buf ( n47 , n418 );
buf ( n49 , n422 );
buf ( n55 , n426 );
buf ( n57 , n430 );
buf ( n48 , n434 );
buf ( n54 , n438 );
buf ( n46 , n441 );
buf ( n120 , n4 );
buf ( n121 , n25 );
buf ( n122 , n40 );
buf ( n123 , n24 );
buf ( n124 , n3 );
buf ( n125 , n38 );
buf ( n126 , n9 );
buf ( n127 , n39 );
buf ( n128 , n33 );
buf ( n129 , n14 );
buf ( n130 , n17 );
buf ( n131 , n2 );
buf ( n132 , n15 );
buf ( n133 , n10 );
buf ( n134 , n37 );
buf ( n135 , n32 );
buf ( n136 , n31 );
buf ( n137 , n19 );
buf ( n138 , n8 );
buf ( n139 , n7 );
buf ( n140 , n18 );
buf ( n141 , n21 );
buf ( n142 , n12 );
buf ( n143 , n23 );
buf ( n144 , n34 );
buf ( n145 , n36 );
buf ( n146 , n1 );
buf ( n147 , n42 );
buf ( n148 , n11 );
buf ( n149 , n30 );
buf ( n150 , n20 );
buf ( n151 , n35 );
buf ( n152 , n26 );
buf ( n153 , n13 );
buf ( n154 , n16 );
buf ( n155 , n0 );
buf ( n156 , n41 );
buf ( n157 , n28 );
buf ( n158 , n22 );
buf ( n159 , n27 );
buf ( n160 , n29 );
buf ( n161 , n6 );
buf ( n162 , n120 );
buf ( n163 , n121 );
buf ( n164 , n122 );
buf ( n165 , n123 );
buf ( n166 , n152 );
and ( n167 , n165 , n166 );
buf ( n168 , n124 );
buf ( n169 , n153 );
and ( n170 , n168 , n169 );
buf ( n171 , n125 );
buf ( n172 , n154 );
and ( n173 , n171 , n172 );
buf ( n174 , n126 );
buf ( n175 , n155 );
and ( n176 , n174 , n175 );
buf ( n177 , n127 );
buf ( n178 , n156 );
and ( n179 , n177 , n178 );
buf ( n180 , n128 );
buf ( n181 , n157 );
and ( n182 , n180 , n181 );
buf ( n183 , n129 );
buf ( n184 , n158 );
and ( n185 , n183 , n184 );
buf ( n186 , n130 );
buf ( n187 , n159 );
and ( n188 , n186 , n187 );
buf ( n189 , n131 );
buf ( n190 , n160 );
and ( n191 , n189 , n190 );
buf ( n192 , n132 );
buf ( n193 , n161 );
and ( n194 , n192 , n193 );
buf ( n195 , n133 );
buf ( n196 , n134 );
buf ( n197 , n135 );
or ( n198 , n196 , n197 );
or ( n199 , n195 , n198 );
and ( n200 , n193 , n199 );
and ( n201 , n192 , n199 );
or ( n202 , n194 , n200 , n201 );
and ( n203 , n190 , n202 );
and ( n204 , n189 , n202 );
or ( n205 , n191 , n203 , n204 );
and ( n206 , n187 , n205 );
and ( n207 , n186 , n205 );
or ( n208 , n188 , n206 , n207 );
and ( n209 , n184 , n208 );
and ( n210 , n183 , n208 );
or ( n211 , n185 , n209 , n210 );
and ( n212 , n181 , n211 );
and ( n213 , n180 , n211 );
or ( n214 , n182 , n212 , n213 );
and ( n215 , n178 , n214 );
and ( n216 , n177 , n214 );
or ( n217 , n179 , n215 , n216 );
and ( n218 , n175 , n217 );
and ( n219 , n174 , n217 );
or ( n220 , n176 , n218 , n219 );
and ( n221 , n172 , n220 );
and ( n222 , n171 , n220 );
or ( n223 , n173 , n221 , n222 );
and ( n224 , n169 , n223 );
and ( n225 , n168 , n223 );
or ( n226 , n170 , n224 , n225 );
and ( n227 , n166 , n226 );
and ( n228 , n165 , n226 );
or ( n229 , n167 , n227 , n228 );
and ( n230 , n164 , n229 );
and ( n231 , n163 , n230 );
xor ( n232 , n162 , n231 );
buf ( n233 , n232 );
buf ( n234 , n233 );
buf ( n235 , n136 );
not ( n236 , n235 );
xor ( n237 , n234 , n236 );
xor ( n238 , n163 , n230 );
buf ( n239 , n238 );
buf ( n240 , n239 );
buf ( n241 , n137 );
not ( n242 , n241 );
and ( n243 , n240 , n242 );
xor ( n244 , n164 , n229 );
buf ( n245 , n244 );
buf ( n246 , n245 );
buf ( n247 , n138 );
not ( n248 , n247 );
and ( n249 , n246 , n248 );
xor ( n250 , n165 , n166 );
xor ( n251 , n250 , n226 );
buf ( n252 , n251 );
buf ( n253 , n252 );
buf ( n254 , n139 );
not ( n255 , n254 );
and ( n256 , n253 , n255 );
xor ( n257 , n168 , n169 );
xor ( n258 , n257 , n223 );
buf ( n259 , n258 );
buf ( n260 , n259 );
buf ( n261 , n140 );
not ( n262 , n261 );
and ( n263 , n260 , n262 );
xor ( n264 , n171 , n172 );
xor ( n265 , n264 , n220 );
buf ( n266 , n265 );
buf ( n267 , n266 );
buf ( n268 , n141 );
not ( n269 , n268 );
and ( n270 , n267 , n269 );
xor ( n271 , n174 , n175 );
xor ( n272 , n271 , n217 );
buf ( n273 , n272 );
buf ( n274 , n273 );
buf ( n275 , n142 );
not ( n276 , n275 );
and ( n277 , n274 , n276 );
xor ( n278 , n177 , n178 );
xor ( n279 , n278 , n214 );
buf ( n280 , n279 );
buf ( n281 , n280 );
buf ( n282 , n143 );
not ( n283 , n282 );
and ( n284 , n281 , n283 );
xor ( n285 , n180 , n181 );
xor ( n286 , n285 , n211 );
buf ( n287 , n286 );
buf ( n288 , n287 );
buf ( n289 , n144 );
not ( n290 , n289 );
and ( n291 , n288 , n290 );
xor ( n292 , n183 , n184 );
xor ( n293 , n292 , n208 );
buf ( n294 , n293 );
buf ( n295 , n294 );
buf ( n296 , n145 );
not ( n297 , n296 );
and ( n298 , n295 , n297 );
xor ( n299 , n186 , n187 );
xor ( n300 , n299 , n205 );
buf ( n301 , n300 );
buf ( n302 , n301 );
buf ( n303 , n146 );
not ( n304 , n303 );
and ( n305 , n302 , n304 );
xor ( n306 , n189 , n190 );
xor ( n307 , n306 , n202 );
buf ( n308 , n307 );
buf ( n309 , n308 );
buf ( n310 , n147 );
not ( n311 , n310 );
and ( n312 , n309 , n311 );
xor ( n313 , n192 , n193 );
xor ( n314 , n313 , n199 );
buf ( n315 , n314 );
buf ( n316 , n315 );
buf ( n317 , n148 );
not ( n318 , n317 );
and ( n319 , n316 , n318 );
xnor ( n320 , n195 , n198 );
buf ( n321 , n320 );
buf ( n322 , n321 );
buf ( n323 , n149 );
not ( n324 , n323 );
and ( n325 , n322 , n324 );
xnor ( n326 , n196 , n197 );
buf ( n327 , n326 );
buf ( n328 , n327 );
buf ( n329 , n150 );
not ( n330 , n329 );
and ( n331 , n328 , n330 );
not ( n332 , n197 );
buf ( n333 , n332 );
buf ( n334 , n333 );
buf ( n335 , n151 );
not ( n336 , n335 );
or ( n337 , n334 , n336 );
and ( n338 , n330 , n337 );
and ( n339 , n328 , n337 );
or ( n340 , n331 , n338 , n339 );
and ( n341 , n324 , n340 );
and ( n342 , n322 , n340 );
or ( n343 , n325 , n341 , n342 );
and ( n344 , n318 , n343 );
and ( n345 , n316 , n343 );
or ( n346 , n319 , n344 , n345 );
and ( n347 , n311 , n346 );
and ( n348 , n309 , n346 );
or ( n349 , n312 , n347 , n348 );
and ( n350 , n304 , n349 );
and ( n351 , n302 , n349 );
or ( n352 , n305 , n350 , n351 );
and ( n353 , n297 , n352 );
and ( n354 , n295 , n352 );
or ( n355 , n298 , n353 , n354 );
and ( n356 , n290 , n355 );
and ( n357 , n288 , n355 );
or ( n358 , n291 , n356 , n357 );
and ( n359 , n283 , n358 );
and ( n360 , n281 , n358 );
or ( n361 , n284 , n359 , n360 );
and ( n362 , n276 , n361 );
and ( n363 , n274 , n361 );
or ( n364 , n277 , n362 , n363 );
and ( n365 , n269 , n364 );
and ( n366 , n267 , n364 );
or ( n367 , n270 , n365 , n366 );
and ( n368 , n262 , n367 );
and ( n369 , n260 , n367 );
or ( n370 , n263 , n368 , n369 );
and ( n371 , n255 , n370 );
and ( n372 , n253 , n370 );
or ( n373 , n256 , n371 , n372 );
and ( n374 , n248 , n373 );
and ( n375 , n246 , n373 );
or ( n376 , n249 , n374 , n375 );
and ( n377 , n242 , n376 );
and ( n378 , n240 , n376 );
or ( n379 , n243 , n377 , n378 );
xor ( n380 , n237 , n379 );
buf ( n381 , n380 );
buf ( n382 , n381 );
xor ( n383 , n240 , n242 );
xor ( n384 , n383 , n376 );
buf ( n385 , n384 );
buf ( n386 , n385 );
xor ( n387 , n246 , n248 );
xor ( n388 , n387 , n373 );
buf ( n389 , n388 );
buf ( n390 , n389 );
xor ( n391 , n253 , n255 );
xor ( n392 , n391 , n370 );
buf ( n393 , n392 );
buf ( n394 , n393 );
xor ( n395 , n260 , n262 );
xor ( n396 , n395 , n367 );
buf ( n397 , n396 );
buf ( n398 , n397 );
xor ( n399 , n267 , n269 );
xor ( n400 , n399 , n364 );
buf ( n401 , n400 );
buf ( n402 , n401 );
xor ( n403 , n274 , n276 );
xor ( n404 , n403 , n361 );
buf ( n405 , n404 );
buf ( n406 , n405 );
xor ( n407 , n281 , n283 );
xor ( n408 , n407 , n358 );
buf ( n409 , n408 );
buf ( n410 , n409 );
xor ( n411 , n288 , n290 );
xor ( n412 , n411 , n355 );
buf ( n413 , n412 );
buf ( n414 , n413 );
xor ( n415 , n295 , n297 );
xor ( n416 , n415 , n352 );
buf ( n417 , n416 );
buf ( n418 , n417 );
xor ( n419 , n302 , n304 );
xor ( n420 , n419 , n349 );
buf ( n421 , n420 );
buf ( n422 , n421 );
xor ( n423 , n309 , n311 );
xor ( n424 , n423 , n346 );
buf ( n425 , n424 );
buf ( n426 , n425 );
xor ( n427 , n316 , n318 );
xor ( n428 , n427 , n343 );
buf ( n429 , n428 );
buf ( n430 , n429 );
xor ( n431 , n322 , n324 );
xor ( n432 , n431 , n340 );
buf ( n433 , n432 );
buf ( n434 , n433 );
xor ( n435 , n328 , n330 );
xor ( n436 , n435 , n337 );
buf ( n437 , n436 );
buf ( n438 , n437 );
xor ( n439 , n334 , n335 );
buf ( n440 , n439 );
buf ( n441 , n440 );
endmodule

