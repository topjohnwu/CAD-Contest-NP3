//
// Conformal-LEC Version 16.10-d160 ( 04-Jul-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
output n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;

wire n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , 
     n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , 
     n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , 
     n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , 
     n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , 
     n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , 
     n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , 
     n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
     n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
     n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , 
     n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , 
     n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , 
     n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , 
     n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , 
     n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , 
     n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , 
     n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , 
     n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , 
     n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , 
     n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , 
     n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , 
     n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
     n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
     n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
     n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
     n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , 
     n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , 
     n357 ;
buf ( n39 , n204 );
buf ( n36 , n221 );
buf ( n41 , n238 );
buf ( n43 , n255 );
buf ( n37 , n272 );
buf ( n34 , n289 );
buf ( n35 , n306 );
buf ( n38 , n316 );
buf ( n40 , n335 );
buf ( n42 , n349 );
buf ( n125 , n4 );
buf ( n126 , n27 );
buf ( n127 , n3 );
buf ( n128 , n12 );
buf ( n129 , n17 );
buf ( n130 , n18 );
buf ( n131 , n2 );
buf ( n132 , n31 );
buf ( n133 , n5 );
buf ( n134 , n33 );
buf ( n135 , n10 );
buf ( n136 , n11 );
buf ( n137 , n20 );
buf ( n138 , n22 );
buf ( n139 , n29 );
buf ( n140 , n24 );
buf ( n141 , n16 );
buf ( n142 , n8 );
buf ( n143 , n26 );
buf ( n144 , n14 );
buf ( n145 , n19 );
buf ( n146 , n13 );
buf ( n147 , n7 );
buf ( n148 , n23 );
buf ( n149 , n25 );
buf ( n150 , n0 );
buf ( n151 , n15 );
buf ( n152 , n30 );
buf ( n153 , n1 );
buf ( n154 , n28 );
buf ( n155 , n6 );
buf ( n156 , n9 );
buf ( n157 , n21 );
buf ( n158 , n32 );
not ( n159 , n156 );
not ( n160 , n146 );
not ( n161 , n147 );
not ( n162 , n148 );
not ( n163 , n149 );
not ( n164 , n151 );
not ( n165 , n152 );
nor ( n166 , n160 , n161 , n162 , n163 , n150 , n164 , n165 , n153 , n154 , n155 );
not ( n167 , n166 );
and ( n168 , n167 , n125 );
not ( n169 , n135 );
and ( n170 , n169 , n125 );
buf ( n171 , n125 );
buf ( n172 , n126 );
buf ( n173 , n127 );
buf ( n174 , n128 );
buf ( n175 , n129 );
buf ( n176 , n130 );
buf ( n177 , n131 );
buf ( n178 , n132 );
buf ( n179 , n133 );
buf ( n180 , n134 );
and ( n181 , n179 , n180 );
and ( n182 , n178 , n181 );
and ( n183 , n177 , n182 );
and ( n184 , n176 , n183 );
and ( n185 , n175 , n184 );
and ( n186 , n174 , n185 );
and ( n187 , n173 , n186 );
and ( n188 , n172 , n187 );
xor ( n189 , n171 , n188 );
buf ( n190 , n189 );
and ( n191 , n190 , n135 );
or ( n192 , n170 , n191 );
not ( n193 , n138 );
not ( n194 , n139 );
not ( n195 , n145 );
or ( n196 , n136 , n137 , n193 , n194 , n140 , n141 , n142 , n143 , n144 , n195 );
and ( n197 , n192 , n196 );
or ( n198 , 1'b0 , n197 );
and ( n199 , n198 , n166 );
or ( n200 , n168 , n199 );
and ( n201 , n159 , n200 );
or ( n202 , n201 , 1'b0 );
buf ( n203 , n202 );
buf ( n204 , n203 );
not ( n205 , n156 );
not ( n206 , n166 );
and ( n207 , n206 , n126 );
not ( n208 , n135 );
and ( n209 , n208 , n126 );
xor ( n210 , n172 , n187 );
buf ( n211 , n210 );
and ( n212 , n211 , n135 );
or ( n213 , n209 , n212 );
and ( n214 , n213 , n196 );
or ( n215 , 1'b0 , n214 );
and ( n216 , n215 , n166 );
or ( n217 , n207 , n216 );
and ( n218 , n205 , n217 );
or ( n219 , n218 , 1'b0 );
buf ( n220 , n219 );
buf ( n221 , n220 );
not ( n222 , n156 );
not ( n223 , n166 );
and ( n224 , n223 , n127 );
not ( n225 , n135 );
and ( n226 , n225 , n127 );
xor ( n227 , n173 , n186 );
buf ( n228 , n227 );
and ( n229 , n228 , n135 );
or ( n230 , n226 , n229 );
and ( n231 , n230 , n196 );
or ( n232 , 1'b0 , n231 );
and ( n233 , n232 , n166 );
or ( n234 , n224 , n233 );
and ( n235 , n222 , n234 );
or ( n236 , n235 , 1'b0 );
buf ( n237 , n236 );
buf ( n238 , n237 );
not ( n239 , n156 );
not ( n240 , n166 );
and ( n241 , n240 , n128 );
not ( n242 , n135 );
and ( n243 , n242 , n128 );
xor ( n244 , n174 , n185 );
buf ( n245 , n244 );
and ( n246 , n245 , n135 );
or ( n247 , n243 , n246 );
and ( n248 , n247 , n196 );
or ( n249 , 1'b0 , n248 );
and ( n250 , n249 , n166 );
or ( n251 , n241 , n250 );
and ( n252 , n239 , n251 );
or ( n253 , n252 , 1'b0 );
buf ( n254 , n253 );
buf ( n255 , n254 );
not ( n256 , n156 );
not ( n257 , n166 );
and ( n258 , n257 , n129 );
not ( n259 , n135 );
and ( n260 , n259 , n129 );
xor ( n261 , n175 , n184 );
buf ( n262 , n261 );
and ( n263 , n262 , n135 );
or ( n264 , n260 , n263 );
and ( n265 , n264 , n196 );
or ( n266 , 1'b0 , n265 );
and ( n267 , n266 , n166 );
or ( n268 , n258 , n267 );
and ( n269 , n256 , n268 );
or ( n270 , n269 , 1'b0 );
buf ( n271 , n270 );
buf ( n272 , n271 );
not ( n273 , n156 );
not ( n274 , n166 );
and ( n275 , n274 , n130 );
not ( n276 , n135 );
and ( n277 , n276 , n130 );
xor ( n278 , n176 , n183 );
buf ( n279 , n278 );
and ( n280 , n279 , n135 );
or ( n281 , n277 , n280 );
and ( n282 , n281 , n196 );
or ( n283 , 1'b0 , n282 );
and ( n284 , n283 , n166 );
or ( n285 , n275 , n284 );
and ( n286 , n273 , n285 );
or ( n287 , n286 , 1'b0 );
buf ( n288 , n287 );
buf ( n289 , n288 );
not ( n290 , n156 );
not ( n291 , n166 );
and ( n292 , n291 , n131 );
not ( n293 , n135 );
and ( n294 , n293 , n131 );
xor ( n295 , n177 , n182 );
buf ( n296 , n295 );
and ( n297 , n296 , n135 );
or ( n298 , n294 , n297 );
and ( n299 , n298 , n196 );
or ( n300 , 1'b0 , n299 );
and ( n301 , n300 , n166 );
or ( n302 , n292 , n301 );
and ( n303 , n290 , n302 );
or ( n304 , n303 , 1'b0 );
buf ( n305 , n304 );
buf ( n306 , n305 );
or ( n307 , n156 , n166 );
not ( n308 , n307 );
nor ( n309 , n160 , n161 , n162 , n163 , n150 , n151 , n152 , n153 , n154 , n155 );
not ( n310 , n309 );
and ( n311 , n157 , n310 );
and ( n312 , n308 , n311 );
and ( n313 , 1'b1 , n307 );
or ( n314 , n312 , n313 );
buf ( n315 , n314 );
buf ( n316 , n315 );
not ( n317 , n156 );
not ( n318 , n166 );
and ( n319 , n318 , n158 );
nor ( n320 , n136 , n137 , n193 , n194 , n140 , n141 , n142 , n143 , n144 , n145 );
not ( n321 , n320 );
not ( n322 , n137 );
nor ( n323 , n136 , n322 , n138 , n194 , n140 , n141 , n142 , n143 , n144 , n145 );
not ( n324 , n323 );
and ( n325 , n158 , n324 );
and ( n326 , n321 , n325 );
and ( n327 , 1'b1 , n320 );
or ( n328 , n326 , n327 );
and ( n329 , n328 , n166 );
or ( n330 , n319 , n329 );
and ( n331 , n317 , n330 );
and ( n332 , 1'b1 , n156 );
or ( n333 , n331 , n332 );
buf ( n334 , n333 );
buf ( n335 , n334 );
not ( n336 , n156 );
not ( n337 , n166 );
and ( n338 , n337 , n136 );
buf ( n339 , n136 );
not ( n340 , n339 );
buf ( n341 , n340 );
and ( n342 , n341 , n196 );
or ( n343 , 1'b0 , n342 );
and ( n344 , n343 , n166 );
or ( n345 , n338 , n344 );
and ( n346 , n336 , n345 );
or ( n347 , n346 , 1'b0 );
buf ( n348 , n347 );
buf ( n349 , n348 );
not ( n350 , n196 );
not ( n351 , n196 );
not ( n352 , n196 );
not ( n353 , n196 );
not ( n354 , n196 );
not ( n355 , n196 );
not ( n356 , n196 );
not ( n357 , n196 );
endmodule

