//
// Conformal-LEC Version 15.20-d235 ( 27-Mar-2016) ( 64 bit executable)
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 ;
output n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 ;

wire n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
     n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
     n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
     n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
     n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
     n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
     n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
     n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
     n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , 
     n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , 
     n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , 
     n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , 
     n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , 
     n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , 
     n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , 
     n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , 
     n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , 
     n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , 
     n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , 
     n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , 
     n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , 
     n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , 
     n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , 
     n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , 
     n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , 
     n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , 
     n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , 
     n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , 
     n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , 
     n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , 
     n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , 
     n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , 
     n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , 
     n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , 
     n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , 
     n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , 
     n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , 
     n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , 
     n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , 
     n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , 
     n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , 
     n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , 
     n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , 
     n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , 
     n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , 
     n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , 
     n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , 
     n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , 
     n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , 
     n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , 
     n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , 
     n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , 
     n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , 
     n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , 
     n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , 
     n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , 
     n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , 
     n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , 
     n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , 
     n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , 
     n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , 
     n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , 
     n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , 
     n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , 
     n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , 
     n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , 
     n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , 
     n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , 
     n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , 
     n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , 
     n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , 
     n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , 
     n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , 
     n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , 
     n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , 
     n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , 
     n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , 
     n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , 
     n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , 
     n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , 
     n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , 
     n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , 
     n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , 
     n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , 
     n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , 
     n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , 
     n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , 
     n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , 
     n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , 
     n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , 
     n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , 
     n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , 
     n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , 
     n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , 
     n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , 
     n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , 
     n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , 
     n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , 
     n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , 
     n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , 
     n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , 
     n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , 
     n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , 
     n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , 
     n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , 
     n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , 
     n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , 
     n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , 
     n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , 
     n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , 
     n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , 
     n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , 
     n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , 
     n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , 
     n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , 
     n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , 
     n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , 
     n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , 
     n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , 
     n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , 
     n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , 
     n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , 
     n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , 
     n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , 
     n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , 
     n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , 
     n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , 
     n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , 
     n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , 
     n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , 
     n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , 
     n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , 
     n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , 
     n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , 
     n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , 
     n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , 
     n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , 
     n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , 
     n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , 
     n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , 
     n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , 
     n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , 
     n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , 
     n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , 
     n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , 
     n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , 
     n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , 
     n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , 
     n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , 
     n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , 
     n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , 
     n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , 
     n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , 
     n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , 
     n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , 
     n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , 
     n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , 
     n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , 
     n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , 
     n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , 
     n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , 
     n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , 
     n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , 
     n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , 
     n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , 
     n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , 
     n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , 
     n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , 
     n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , 
     n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , 
     n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , 
     n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , 
     n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , 
     n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , 
     n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , 
     n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , 
     n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , 
     n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , 
     n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , 
     n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , 
     n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , 
     n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , 
     n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , 
     n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , 
     n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , 
     n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , 
     n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , 
     n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , 
     n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , 
     n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , 
     n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , 
     n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , 
     n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , 
     n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , 
     n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , 
     n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , 
     n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , 
     n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , 
     n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , 
     n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , 
     n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , 
     n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , 
     n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , 
     n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , 
     n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , 
     n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , 
     n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , 
     n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , 
     n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , 
     n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , 
     n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , 
     n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , 
     n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , 
     n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , 
     n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , 
     n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , 
     n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , 
     n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , 
     n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , 
     n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , 
     n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
     n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , 
     n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , 
     n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , 
     n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , 
     n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , 
     n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , 
     n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , 
     n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , 
     n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , 
     n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , 
     n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , 
     n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , 
     n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , 
     n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , 
     n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , 
     n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , 
     n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , 
     n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , 
     n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , 
     n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , 
     n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , 
     n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , 
     n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , 
     n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , 
     n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , 
     n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
     n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , 
     n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , 
     n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , 
     n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , 
     n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , 
     n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , 
     n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , 
     n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , 
     n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , 
     n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , 
     n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , 
     n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , 
     n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , 
     n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , 
     n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , 
     n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , 
     n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , 
     n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , 
     n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , 
     n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , 
     n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , 
     n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , 
     n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , 
     n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , 
     n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , 
     n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , 
     n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , 
     n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , 
     n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , 
     n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , 
     n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , 
     n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , 
     n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , 
     n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , 
     n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , 
     n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , 
     n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , 
     n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , 
     n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , 
     n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , 
     n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , 
     n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , 
     n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , 
     n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , 
     n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , 
     n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , 
     n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
     n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
     n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , 
     n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , 
     n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , 
     n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , 
     n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , 
     n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , 
     n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , 
     n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , 
     n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , 
     n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , 
     n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , 
     n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , 
     n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , 
     n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , 
     n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , 
     n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , 
     n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , 
     n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , 
     n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , 
     n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , 
     n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , 
     n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , 
     n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , 
     n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , 
     n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , 
     n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , 
     n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , 
     n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , 
     n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , 
     n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , 
     n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , 
     n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , 
     n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , 
     n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , 
     n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
     n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
     n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , 
     n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , 
     n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , 
     n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , 
     n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , 
     n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , 
     n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , 
     n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , 
     n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , 
     n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , 
     n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , 
     n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , 
     n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , 
     n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , 
     n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , 
     n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , 
     n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , 
     n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , 
     n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , 
     n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , 
     n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , 
     n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , 
     n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , 
     n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , 
     n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , 
     n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , 
     n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , 
     n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , 
     n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , 
     n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , 
     n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , 
     n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , 
     n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , 
     n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , 
     n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , 
     n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , 
     n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , 
     n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , 
     n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , 
     n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , 
     n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , 
     n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , 
     n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , 
     n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , 
     n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , 
     n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , 
     n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , 
     n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , 
     n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , 
     n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , 
     n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , 
     n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , 
     n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , 
     n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , 
     n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , 
     n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , 
     n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , 
     n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , 
     n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , 
     n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , 
     n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , 
     n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , 
     n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , 
     n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , 
     n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , 
     n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , 
     n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , 
     n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , 
     n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , 
     n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , 
     n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , 
     n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , 
     n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , 
     n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , 
     n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , 
     n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , 
     n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , 
     n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , 
     n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , 
     n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , 
     n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , 
     n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , 
     n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
     n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
     n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , 
     n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , 
     n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , 
     n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , 
     n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , 
     n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
     n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
     n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
     n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
     n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
     n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
     n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
     n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
     n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
     n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
     n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
     n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
     n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
     n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
     n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
     n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
     n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
     n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
     n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
     n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
     n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
     n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
     n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
     n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
     n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , 
     n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , 
     n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
     n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , 
     n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
     n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , 
     n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
     n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
     n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
     n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , 
     n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
     n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
     n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
     n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
     n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
     n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
     n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
     n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
     n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
     n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
     n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
     n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
     n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , 
     n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , 
     n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , 
     n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , 
     n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , 
     n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , 
     n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , 
     n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
     n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , 
     n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , 
     n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , 
     n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , 
     n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , 
     n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , 
     n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , 
     n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , 
     n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , 
     n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , 
     n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , 
     n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , 
     n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , 
     n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , 
     n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
     n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
     n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
     n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
     n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
     n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
     n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
     n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
     n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
     n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
     n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
     n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
     n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
     n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
     n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , 
     n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , 
     n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
     n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , 
     n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , 
     n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , 
     n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , 
     n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , 
     n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , 
     n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , 
     n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , 
     n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
     n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , 
     n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , 
     n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , 
     n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
     n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , 
     n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , 
     n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
     n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , 
     n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , 
     n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , 
     n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , 
     n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , 
     n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , 
     n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , 
     n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , 
     n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , 
     n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , 
     n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , 
     n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , 
     n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , 
     n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , 
     n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , 
     n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , 
     n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , 
     n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , 
     n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
     n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , 
     n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , 
     n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , 
     n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , 
     n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , 
     n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , 
     n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , 
     n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , 
     n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , 
     n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , 
     n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , 
     n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , 
     n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , 
     n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , 
     n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , 
     n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , 
     n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , 
     n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , 
     n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , 
     n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , 
     n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , 
     n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , 
     n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , 
     n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , 
     n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , 
     n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , 
     n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , 
     n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , 
     n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , 
     n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , 
     n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , 
     n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , 
     n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , 
     n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , 
     n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , 
     n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , 
     n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , 
     n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , 
     n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , 
     n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , 
     n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , 
     n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , 
     n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , 
     n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , 
     n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , 
     n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , 
     n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , 
     n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , 
     n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , 
     n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , 
     n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , 
     n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , 
     n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , 
     n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , 
     n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , 
     n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , 
     n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , 
     n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , 
     n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , 
     n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , 
     n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , 
     n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , 
     n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , 
     n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , 
     n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , 
     n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , 
     n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , 
     n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , 
     n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , 
     n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , 
     n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , 
     n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , 
     n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , 
     n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , 
     n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , 
     n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , 
     n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , 
     n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , 
     n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , 
     n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , 
     n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , 
     n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , 
     n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , 
     n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , 
     n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , 
     n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , 
     n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , 
     n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , 
     n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , 
     n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , 
     n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , 
     n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , 
     n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , 
     n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , 
     n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , 
     n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , 
     n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , 
     n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , 
     n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , 
     n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , 
     n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , 
     n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , 
     n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , 
     n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , 
     n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , 
     n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , 
     n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , 
     n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , 
     n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , 
     n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , 
     n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , 
     n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , 
     n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , 
     n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , 
     n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , 
     n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , 
     n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , 
     n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , 
     n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , 
     n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , 
     n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , 
     n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , 
     n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , 
     n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , 
     n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , 
     n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , 
     n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , 
     n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , 
     n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , 
     n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , 
     n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , 
     n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , 
     n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , 
     n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , 
     n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , 
     n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , 
     n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , 
     n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , 
     n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , 
     n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , 
     n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , 
     n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , 
     n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , 
     n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , 
     n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , 
     n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , 
     n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , 
     n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , 
     n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , 
     n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , 
     n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , 
     n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , 
     n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , 
     n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , 
     n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , 
     n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , 
     n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , 
     n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , 
     n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , 
     n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , 
     n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , 
     n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , 
     n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , 
     n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , 
     n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , 
     n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , 
     n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , 
     n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , 
     n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , 
     n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , 
     n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , 
     n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , 
     n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , 
     n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , 
     n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , 
     n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , 
     n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , 
     n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , 
     n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , 
     n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , 
     n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , 
     n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , 
     n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , 
     n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , 
     n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , 
     n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , 
     n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , 
     n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , 
     n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , 
     n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , 
     n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , 
     n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , 
     n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , 
     n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , 
     n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , 
     n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , 
     n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , 
     n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , 
     n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , 
     n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , 
     n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , 
     n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , 
     n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , 
     n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , 
     n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , 
     n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , 
     n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , 
     n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , 
     n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , 
     n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , 
     n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , 
     n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , 
     n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , 
     n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , 
     n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , 
     n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , 
     n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , 
     n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , 
     n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , 
     n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , 
     n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , 
     n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , 
     n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , 
     n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , 
     n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , 
     n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , 
     n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , 
     n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , 
     n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , 
     n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , 
     n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , 
     n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , 
     n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , 
     n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , 
     n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , 
     n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , 
     n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , 
     n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , 
     n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , 
     n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , 
     n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , 
     n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , 
     n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , 
     n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , 
     n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , 
     n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , 
     n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , 
     n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , 
     n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , 
     n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , 
     n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , 
     n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , 
     n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , 
     n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , 
     n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , 
     n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , 
     n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , 
     n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , 
     n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , 
     n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , 
     n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , 
     n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , 
     n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , 
     n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , 
     n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , 
     n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , 
     n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , 
     n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , 
     n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , 
     n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , 
     n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , 
     n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , 
     n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , 
     n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , 
     n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , 
     n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , 
     n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , 
     n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , 
     n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , 
     n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , 
     n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , 
     n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , 
     n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , 
     n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , 
     n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , 
     n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , 
     n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , 
     n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , 
     n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , 
     n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , 
     n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , 
     n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , 
     n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , 
     n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , 
     n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , 
     n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , 
     n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , 
     n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , 
     n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , 
     n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , 
     n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , 
     n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , 
     n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , 
     n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , 
     n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , 
     n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , 
     n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , 
     n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , 
     n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , 
     n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , 
     n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , 
     n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , 
     n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , 
     n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , 
     n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , 
     n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , 
     n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , 
     n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , 
     n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , 
     n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , 
     n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , 
     n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , 
     n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , 
     n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , 
     n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 ;
buf ( n88 , n8792 );
buf ( n91 , n8795 );
buf ( n94 , n8798 );
buf ( n95 , n8801 );
buf ( n80 , n8804 );
buf ( n85 , n8807 );
buf ( n86 , n8810 );
buf ( n89 , n8813 );
buf ( n81 , n8816 );
buf ( n83 , n8819 );
buf ( n93 , n8822 );
buf ( n87 , n8825 );
buf ( n90 , n8828 );
buf ( n82 , n8831 );
buf ( n84 , n8834 );
buf ( n92 , n8837 );
buf ( n195 , n21 );
buf ( n196 , n59 );
buf ( n197 , n25 );
buf ( n198 , n12 );
buf ( n199 , n47 );
buf ( n200 , n13 );
buf ( n201 , n36 );
buf ( n202 , n11 );
buf ( n203 , n2 );
buf ( n204 , n37 );
buf ( n205 , n1 );
buf ( n206 , n31 );
buf ( n207 , n8 );
buf ( n208 , n51 );
buf ( n209 , n15 );
buf ( n210 , n20 );
buf ( n211 , n42 );
buf ( n212 , n4 );
buf ( n213 , n50 );
buf ( n214 , n71 );
buf ( n215 , n5 );
buf ( n216 , n32 );
buf ( n217 , n38 );
buf ( n218 , n62 );
buf ( n219 , n57 );
buf ( n220 , n9 );
buf ( n221 , n23 );
buf ( n222 , n67 );
buf ( n223 , n3 );
buf ( n224 , n27 );
buf ( n225 , n41 );
buf ( n226 , n65 );
buf ( n227 , n54 );
buf ( n228 , n18 );
buf ( n229 , n7 );
buf ( n230 , n69 );
buf ( n231 , n6 );
buf ( n232 , n30 );
buf ( n233 , n61 );
buf ( n234 , n63 );
buf ( n235 , n60 );
buf ( n236 , n73 );
buf ( n237 , n49 );
buf ( n238 , n17 );
buf ( n239 , n66 );
buf ( n240 , n48 );
buf ( n241 , n72 );
buf ( n242 , n74 );
buf ( n243 , n46 );
buf ( n244 , n35 );
buf ( n245 , n43 );
buf ( n246 , n40 );
buf ( n247 , n53 );
buf ( n248 , n55 );
buf ( n249 , n79 );
buf ( n250 , n29 );
buf ( n251 , n70 );
buf ( n252 , n56 );
buf ( n253 , n33 );
buf ( n254 , n10 );
buf ( n255 , n19 );
buf ( n256 , n76 );
buf ( n257 , n68 );
buf ( n258 , n39 );
buf ( n259 , n75 );
buf ( n260 , n26 );
buf ( n261 , n0 );
buf ( n262 , n28 );
buf ( n263 , n78 );
buf ( n264 , n52 );
buf ( n265 , n34 );
buf ( n266 , n14 );
buf ( n267 , n44 );
buf ( n268 , n16 );
buf ( n269 , n22 );
buf ( n270 , n24 );
buf ( n271 , n58 );
buf ( n272 , n77 );
buf ( n273 , n225 );
buf ( n274 , n256 );
and ( n275 , n273 , n274 );
buf ( n276 , n275 );
buf ( n277 , n276 );
not ( n278 , n238 );
buf ( n279 , n278 );
and ( n280 , n277 , n279 );
buf ( n281 , n280 );
buf ( n282 , n281 );
not ( n283 , n282 );
buf ( n284 , n195 );
not ( n285 , n284 );
and ( n286 , n285 , n282 );
nor ( n287 , n283 , n286 );
buf ( n288 , n240 );
and ( n289 , n277 , n288 );
buf ( n290 , n289 );
buf ( n291 , n255 );
and ( n292 , n273 , n291 );
buf ( n293 , n292 );
buf ( n294 , n224 );
and ( n295 , n294 , n274 );
xor ( n296 , n293 , n295 );
buf ( n297 , n296 );
buf ( n298 , n297 );
and ( n299 , n298 , n279 );
xor ( n300 , n290 , n299 );
buf ( n301 , n300 );
buf ( n302 , n301 );
not ( n303 , n302 );
buf ( n304 , n196 );
not ( n305 , n304 );
nor ( n306 , n303 , n305 );
xor ( n307 , n287 , n306 );
buf ( n308 , n307 );
and ( n309 , n289 , n299 );
buf ( n310 , n309 );
buf ( n311 , n310 );
buf ( n312 , n239 );
and ( n313 , n277 , n312 );
and ( n314 , n298 , n288 );
xor ( n315 , n313 , n314 );
and ( n316 , n292 , n295 );
buf ( n317 , n316 );
buf ( n318 , n223 );
and ( n319 , n318 , n274 );
xor ( n320 , n317 , n319 );
buf ( n321 , n254 );
and ( n322 , n273 , n321 );
buf ( n323 , n322 );
and ( n324 , n294 , n291 );
xor ( n325 , n323 , n324 );
xor ( n326 , n320 , n325 );
buf ( n327 , n326 );
buf ( n328 , n327 );
and ( n329 , n328 , n279 );
xor ( n330 , n315 , n329 );
xor ( n331 , n311 , n330 );
buf ( n332 , n331 );
buf ( n333 , n332 );
not ( n334 , n333 );
buf ( n335 , n197 );
not ( n336 , n335 );
nor ( n337 , n334 , n336 );
xor ( n338 , n308 , n337 );
nor ( n339 , n283 , n305 );
buf ( n340 , n339 );
nor ( n341 , n303 , n336 );
and ( n342 , n340 , n341 );
buf ( n343 , n342 );
xor ( n344 , n338 , n343 );
and ( n345 , n313 , n314 );
and ( n346 , n314 , n329 );
and ( n347 , n313 , n329 );
or ( n348 , n345 , n346 , n347 );
and ( n349 , n298 , n312 );
and ( n350 , n328 , n288 );
xor ( n351 , n349 , n350 );
and ( n352 , n322 , n324 );
buf ( n353 , n352 );
buf ( n354 , n253 );
and ( n355 , n273 , n354 );
buf ( n356 , n355 );
and ( n357 , n294 , n321 );
xor ( n358 , n356 , n357 );
xor ( n359 , n353 , n358 );
and ( n360 , n318 , n291 );
buf ( n361 , n222 );
and ( n362 , n361 , n274 );
xor ( n363 , n360 , n362 );
xor ( n364 , n359 , n363 );
and ( n365 , n317 , n319 );
and ( n366 , n319 , n325 );
and ( n367 , n317 , n325 );
or ( n368 , n365 , n366 , n367 );
xor ( n369 , n364 , n368 );
buf ( n370 , n369 );
buf ( n371 , n370 );
and ( n372 , n371 , n279 );
xor ( n373 , n351 , n372 );
xor ( n374 , n348 , n373 );
buf ( n375 , n238 );
and ( n376 , n277 , n375 );
buf ( n377 , n376 );
xor ( n378 , n374 , n377 );
and ( n379 , n310 , n330 );
buf ( n380 , n379 );
xor ( n381 , n378 , n380 );
buf ( n382 , n381 );
buf ( n383 , n382 );
not ( n384 , n383 );
buf ( n385 , n198 );
not ( n386 , n385 );
nor ( n387 , n384 , n386 );
xor ( n388 , n344 , n387 );
xor ( n389 , n340 , n341 );
buf ( n390 , n389 );
nor ( n391 , n334 , n386 );
and ( n392 , n390 , n391 );
xor ( n393 , n390 , n391 );
nor ( n394 , n283 , n336 );
buf ( n395 , n394 );
nor ( n396 , n303 , n386 );
and ( n397 , n395 , n396 );
buf ( n398 , n397 );
and ( n399 , n393 , n398 );
or ( n400 , n392 , n399 );
xor ( n401 , n388 , n400 );
and ( n402 , n348 , n373 );
and ( n403 , n373 , n377 );
and ( n404 , n348 , n377 );
or ( n405 , n402 , n403 , n404 );
buf ( n406 , n405 );
and ( n407 , n349 , n350 );
and ( n408 , n350 , n372 );
and ( n409 , n349 , n372 );
or ( n410 , n407 , n408 , n409 );
buf ( n411 , n237 );
and ( n412 , n277 , n411 );
buf ( n413 , n412 );
and ( n414 , n298 , n375 );
xor ( n415 , n413 , n414 );
xor ( n416 , n410 , n415 );
and ( n417 , n328 , n312 );
and ( n418 , n371 , n288 );
xor ( n419 , n417 , n418 );
and ( n420 , n360 , n362 );
and ( n421 , n353 , n358 );
and ( n422 , n358 , n363 );
and ( n423 , n353 , n363 );
or ( n424 , n421 , n422 , n423 );
xor ( n425 , n420 , n424 );
and ( n426 , n355 , n357 );
buf ( n427 , n426 );
and ( n428 , n318 , n321 );
and ( n429 , n361 , n291 );
xor ( n430 , n428 , n429 );
buf ( n431 , n221 );
and ( n432 , n431 , n274 );
xor ( n433 , n430 , n432 );
xor ( n434 , n427 , n433 );
buf ( n435 , n252 );
and ( n436 , n273 , n435 );
buf ( n437 , n436 );
and ( n438 , n294 , n354 );
xor ( n439 , n437 , n438 );
xor ( n440 , n434 , n439 );
xor ( n441 , n425 , n440 );
and ( n442 , n364 , n368 );
buf ( n443 , n442 );
xor ( n444 , n441 , n443 );
buf ( n445 , n444 );
buf ( n446 , n445 );
and ( n447 , n446 , n279 );
xor ( n448 , n419 , n447 );
xor ( n449 , n416 , n448 );
xor ( n450 , n406 , n449 );
and ( n451 , n378 , n380 );
buf ( n452 , n451 );
xor ( n453 , n450 , n452 );
buf ( n454 , n453 );
buf ( n455 , n454 );
not ( n456 , n455 );
buf ( n457 , n199 );
not ( n458 , n457 );
nor ( n459 , n456 , n458 );
xor ( n460 , n401 , n459 );
xor ( n461 , n393 , n398 );
nor ( n462 , n384 , n458 );
and ( n463 , n461 , n462 );
xor ( n464 , n461 , n462 );
xor ( n465 , n395 , n396 );
buf ( n466 , n465 );
nor ( n467 , n334 , n458 );
and ( n468 , n466 , n467 );
xor ( n469 , n466 , n467 );
nor ( n470 , n283 , n386 );
buf ( n471 , n470 );
nor ( n472 , n303 , n458 );
and ( n473 , n471 , n472 );
buf ( n474 , n473 );
and ( n475 , n469 , n474 );
or ( n476 , n468 , n475 );
and ( n477 , n464 , n476 );
or ( n478 , n463 , n477 );
xor ( n479 , n460 , n478 );
and ( n480 , n410 , n415 );
and ( n481 , n415 , n448 );
and ( n482 , n410 , n448 );
or ( n483 , n480 , n481 , n482 );
and ( n484 , n417 , n418 );
and ( n485 , n418 , n447 );
and ( n486 , n417 , n447 );
or ( n487 , n484 , n485 , n486 );
buf ( n488 , n236 );
and ( n489 , n277 , n488 );
and ( n490 , n298 , n411 );
xor ( n491 , n489 , n490 );
and ( n492 , n328 , n375 );
xor ( n493 , n491 , n492 );
xor ( n494 , n487 , n493 );
and ( n495 , n371 , n312 );
and ( n496 , n446 , n288 );
xor ( n497 , n495 , n496 );
and ( n498 , n427 , n433 );
and ( n499 , n433 , n439 );
and ( n500 , n427 , n439 );
or ( n501 , n498 , n499 , n500 );
and ( n502 , n436 , n438 );
buf ( n503 , n502 );
and ( n504 , n318 , n354 );
and ( n505 , n361 , n321 );
xor ( n506 , n504 , n505 );
and ( n507 , n431 , n291 );
xor ( n508 , n506 , n507 );
xor ( n509 , n503 , n508 );
buf ( n510 , n251 );
and ( n511 , n273 , n510 );
buf ( n512 , n511 );
and ( n513 , n294 , n435 );
xor ( n514 , n512 , n513 );
xor ( n515 , n509 , n514 );
xor ( n516 , n501 , n515 );
and ( n517 , n428 , n429 );
and ( n518 , n429 , n432 );
and ( n519 , n428 , n432 );
or ( n520 , n517 , n518 , n519 );
buf ( n521 , n220 );
and ( n522 , n521 , n274 );
xor ( n523 , n520 , n522 );
xor ( n524 , n516 , n523 );
and ( n525 , n420 , n424 );
and ( n526 , n424 , n440 );
and ( n527 , n420 , n440 );
or ( n528 , n525 , n526 , n527 );
xor ( n529 , n524 , n528 );
and ( n530 , n441 , n443 );
xor ( n531 , n529 , n530 );
buf ( n532 , n531 );
buf ( n533 , n532 );
and ( n534 , n533 , n279 );
xor ( n535 , n497 , n534 );
xor ( n536 , n494 , n535 );
xor ( n537 , n483 , n536 );
and ( n538 , n412 , n414 );
buf ( n539 , n538 );
buf ( n540 , n539 );
xor ( n541 , n537 , n540 );
and ( n542 , n405 , n449 );
buf ( n543 , n542 );
xor ( n544 , n541 , n543 );
and ( n545 , n450 , n452 );
xor ( n546 , n544 , n545 );
buf ( n547 , n546 );
buf ( n548 , n547 );
not ( n549 , n548 );
buf ( n550 , n200 );
not ( n551 , n550 );
nor ( n552 , n549 , n551 );
xor ( n553 , n479 , n552 );
xor ( n554 , n464 , n476 );
nor ( n555 , n456 , n551 );
and ( n556 , n554 , n555 );
xor ( n557 , n554 , n555 );
xor ( n558 , n469 , n474 );
nor ( n559 , n384 , n551 );
and ( n560 , n558 , n559 );
xor ( n561 , n558 , n559 );
xor ( n562 , n471 , n472 );
buf ( n563 , n562 );
nor ( n564 , n334 , n551 );
and ( n565 , n563 , n564 );
xor ( n566 , n563 , n564 );
nor ( n567 , n283 , n458 );
buf ( n568 , n567 );
nor ( n569 , n303 , n551 );
and ( n570 , n568 , n569 );
buf ( n571 , n570 );
and ( n572 , n566 , n571 );
or ( n573 , n565 , n572 );
and ( n574 , n561 , n573 );
or ( n575 , n560 , n574 );
and ( n576 , n557 , n575 );
or ( n577 , n556 , n576 );
xor ( n578 , n553 , n577 );
and ( n579 , n483 , n536 );
and ( n580 , n536 , n540 );
and ( n581 , n483 , n540 );
or ( n582 , n579 , n580 , n581 );
buf ( n583 , n582 );
and ( n584 , n487 , n493 );
and ( n585 , n493 , n535 );
and ( n586 , n487 , n535 );
or ( n587 , n584 , n585 , n586 );
and ( n588 , n495 , n496 );
and ( n589 , n496 , n534 );
and ( n590 , n495 , n534 );
or ( n591 , n588 , n589 , n590 );
and ( n592 , n446 , n312 );
and ( n593 , n533 , n288 );
xor ( n594 , n592 , n593 );
and ( n595 , n520 , n522 );
and ( n596 , n501 , n515 );
and ( n597 , n515 , n523 );
and ( n598 , n501 , n523 );
or ( n599 , n596 , n597 , n598 );
xor ( n600 , n595 , n599 );
and ( n601 , n503 , n508 );
and ( n602 , n508 , n514 );
and ( n603 , n503 , n514 );
or ( n604 , n601 , n602 , n603 );
and ( n605 , n511 , n513 );
buf ( n606 , n605 );
buf ( n607 , n250 );
and ( n608 , n273 , n607 );
buf ( n609 , n608 );
and ( n610 , n294 , n510 );
xor ( n611 , n609 , n610 );
xor ( n612 , n606 , n611 );
and ( n613 , n318 , n435 );
and ( n614 , n361 , n354 );
xor ( n615 , n613 , n614 );
and ( n616 , n431 , n321 );
xor ( n617 , n615 , n616 );
xor ( n618 , n612 , n617 );
xor ( n619 , n604 , n618 );
and ( n620 , n504 , n505 );
and ( n621 , n505 , n507 );
and ( n622 , n504 , n507 );
or ( n623 , n620 , n621 , n622 );
and ( n624 , n521 , n291 );
buf ( n625 , n219 );
and ( n626 , n625 , n274 );
xor ( n627 , n624 , n626 );
xor ( n628 , n623 , n627 );
xor ( n629 , n619 , n628 );
xor ( n630 , n600 , n629 );
and ( n631 , n524 , n528 );
and ( n632 , n529 , n530 );
or ( n633 , n631 , n632 );
xor ( n634 , n630 , n633 );
buf ( n635 , n634 );
buf ( n636 , n635 );
and ( n637 , n636 , n279 );
xor ( n638 , n594 , n637 );
xor ( n639 , n591 , n638 );
and ( n640 , n298 , n488 );
and ( n641 , n328 , n411 );
xor ( n642 , n640 , n641 );
and ( n643 , n371 , n375 );
xor ( n644 , n642 , n643 );
xor ( n645 , n639 , n644 );
xor ( n646 , n587 , n645 );
and ( n647 , n489 , n490 );
and ( n648 , n490 , n492 );
and ( n649 , n489 , n492 );
or ( n650 , n647 , n648 , n649 );
buf ( n651 , n235 );
and ( n652 , n277 , n651 );
buf ( n653 , n652 );
xor ( n654 , n650 , n653 );
xor ( n655 , n646 , n654 );
xor ( n656 , n583 , n655 );
and ( n657 , n541 , n543 );
and ( n658 , n544 , n545 );
or ( n659 , n657 , n658 );
xor ( n660 , n656 , n659 );
buf ( n661 , n660 );
buf ( n662 , n661 );
not ( n663 , n662 );
buf ( n664 , n201 );
not ( n665 , n664 );
nor ( n666 , n663 , n665 );
xor ( n667 , n578 , n666 );
xor ( n668 , n557 , n575 );
nor ( n669 , n549 , n665 );
and ( n670 , n668 , n669 );
xor ( n671 , n668 , n669 );
xor ( n672 , n561 , n573 );
nor ( n673 , n456 , n665 );
and ( n674 , n672 , n673 );
xor ( n675 , n672 , n673 );
xor ( n676 , n566 , n571 );
nor ( n677 , n384 , n665 );
and ( n678 , n676 , n677 );
xor ( n679 , n676 , n677 );
xor ( n680 , n568 , n569 );
buf ( n681 , n680 );
nor ( n682 , n334 , n665 );
and ( n683 , n681 , n682 );
xor ( n684 , n681 , n682 );
nor ( n685 , n283 , n551 );
buf ( n686 , n685 );
nor ( n687 , n303 , n665 );
and ( n688 , n686 , n687 );
buf ( n689 , n688 );
and ( n690 , n684 , n689 );
or ( n691 , n683 , n690 );
and ( n692 , n679 , n691 );
or ( n693 , n678 , n692 );
and ( n694 , n675 , n693 );
or ( n695 , n674 , n694 );
and ( n696 , n671 , n695 );
or ( n697 , n670 , n696 );
xor ( n698 , n667 , n697 );
and ( n699 , n650 , n653 );
and ( n700 , n587 , n645 );
and ( n701 , n645 , n654 );
and ( n702 , n587 , n654 );
or ( n703 , n700 , n701 , n702 );
xor ( n704 , n699 , n703 );
and ( n705 , n591 , n638 );
and ( n706 , n638 , n644 );
and ( n707 , n591 , n644 );
or ( n708 , n705 , n706 , n707 );
and ( n709 , n640 , n641 );
and ( n710 , n641 , n643 );
and ( n711 , n640 , n643 );
or ( n712 , n709 , n710 , n711 );
buf ( n713 , n712 );
buf ( n714 , n234 );
and ( n715 , n277 , n714 );
buf ( n716 , n715 );
and ( n717 , n298 , n651 );
xor ( n718 , n716 , n717 );
xor ( n719 , n713 , n718 );
xor ( n720 , n708 , n719 );
and ( n721 , n592 , n593 );
and ( n722 , n593 , n637 );
and ( n723 , n592 , n637 );
or ( n724 , n721 , n722 , n723 );
and ( n725 , n328 , n488 );
and ( n726 , n371 , n411 );
xor ( n727 , n725 , n726 );
and ( n728 , n446 , n375 );
xor ( n729 , n727 , n728 );
xor ( n730 , n724 , n729 );
and ( n731 , n533 , n312 );
and ( n732 , n636 , n288 );
xor ( n733 , n731 , n732 );
and ( n734 , n623 , n627 );
and ( n735 , n604 , n618 );
and ( n736 , n618 , n628 );
and ( n737 , n604 , n628 );
or ( n738 , n735 , n736 , n737 );
xor ( n739 , n734 , n738 );
and ( n740 , n606 , n611 );
and ( n741 , n611 , n617 );
and ( n742 , n606 , n617 );
or ( n743 , n740 , n741 , n742 );
and ( n744 , n613 , n614 );
and ( n745 , n614 , n616 );
and ( n746 , n613 , n616 );
or ( n747 , n744 , n745 , n746 );
and ( n748 , n624 , n626 );
xor ( n749 , n747 , n748 );
and ( n750 , n521 , n321 );
and ( n751 , n625 , n291 );
xor ( n752 , n750 , n751 );
buf ( n753 , n218 );
and ( n754 , n753 , n274 );
xor ( n755 , n752 , n754 );
xor ( n756 , n749 , n755 );
xor ( n757 , n743 , n756 );
and ( n758 , n608 , n610 );
buf ( n759 , n758 );
and ( n760 , n318 , n510 );
and ( n761 , n361 , n435 );
xor ( n762 , n760 , n761 );
and ( n763 , n431 , n354 );
xor ( n764 , n762 , n763 );
xor ( n765 , n759 , n764 );
buf ( n766 , n249 );
and ( n767 , n273 , n766 );
buf ( n768 , n767 );
and ( n769 , n294 , n607 );
xor ( n770 , n768 , n769 );
xor ( n771 , n765 , n770 );
xor ( n772 , n757 , n771 );
xor ( n773 , n739 , n772 );
and ( n774 , n595 , n599 );
and ( n775 , n599 , n629 );
and ( n776 , n595 , n629 );
or ( n777 , n774 , n775 , n776 );
xor ( n778 , n773 , n777 );
and ( n779 , n630 , n633 );
xor ( n780 , n778 , n779 );
buf ( n781 , n780 );
buf ( n782 , n781 );
and ( n783 , n782 , n279 );
xor ( n784 , n733 , n783 );
xor ( n785 , n730 , n784 );
xor ( n786 , n720 , n785 );
xor ( n787 , n704 , n786 );
and ( n788 , n582 , n655 );
buf ( n789 , n788 );
xor ( n790 , n787 , n789 );
and ( n791 , n656 , n659 );
xor ( n792 , n790 , n791 );
buf ( n793 , n792 );
buf ( n794 , n793 );
not ( n795 , n794 );
buf ( n796 , n202 );
not ( n797 , n796 );
nor ( n798 , n795 , n797 );
xor ( n799 , n698 , n798 );
xor ( n800 , n671 , n695 );
nor ( n801 , n663 , n797 );
and ( n802 , n800 , n801 );
xor ( n803 , n800 , n801 );
xor ( n804 , n675 , n693 );
nor ( n805 , n549 , n797 );
and ( n806 , n804 , n805 );
xor ( n807 , n804 , n805 );
xor ( n808 , n679 , n691 );
nor ( n809 , n456 , n797 );
and ( n810 , n808 , n809 );
xor ( n811 , n808 , n809 );
xor ( n812 , n684 , n689 );
nor ( n813 , n384 , n797 );
and ( n814 , n812 , n813 );
xor ( n815 , n812 , n813 );
xor ( n816 , n686 , n687 );
buf ( n817 , n816 );
nor ( n818 , n334 , n797 );
and ( n819 , n817 , n818 );
xor ( n820 , n817 , n818 );
nor ( n821 , n283 , n665 );
buf ( n822 , n821 );
nor ( n823 , n303 , n797 );
and ( n824 , n822 , n823 );
buf ( n825 , n824 );
and ( n826 , n820 , n825 );
or ( n827 , n819 , n826 );
and ( n828 , n815 , n827 );
or ( n829 , n814 , n828 );
and ( n830 , n811 , n829 );
or ( n831 , n810 , n830 );
and ( n832 , n807 , n831 );
or ( n833 , n806 , n832 );
and ( n834 , n803 , n833 );
or ( n835 , n802 , n834 );
xor ( n836 , n799 , n835 );
and ( n837 , n708 , n719 );
and ( n838 , n719 , n785 );
and ( n839 , n708 , n785 );
or ( n840 , n837 , n838 , n839 );
and ( n841 , n724 , n729 );
and ( n842 , n729 , n784 );
and ( n843 , n724 , n784 );
or ( n844 , n841 , n842 , n843 );
and ( n845 , n715 , n717 );
buf ( n846 , n845 );
and ( n847 , n725 , n726 );
and ( n848 , n726 , n728 );
and ( n849 , n725 , n728 );
or ( n850 , n847 , n848 , n849 );
xor ( n851 , n846 , n850 );
buf ( n852 , n233 );
and ( n853 , n277 , n852 );
and ( n854 , n298 , n714 );
xor ( n855 , n853 , n854 );
and ( n856 , n328 , n651 );
xor ( n857 , n855 , n856 );
xor ( n858 , n851 , n857 );
xor ( n859 , n844 , n858 );
and ( n860 , n731 , n732 );
and ( n861 , n732 , n783 );
and ( n862 , n731 , n783 );
or ( n863 , n860 , n861 , n862 );
and ( n864 , n371 , n488 );
and ( n865 , n446 , n411 );
xor ( n866 , n864 , n865 );
and ( n867 , n533 , n375 );
xor ( n868 , n866 , n867 );
xor ( n869 , n863 , n868 );
and ( n870 , n636 , n312 );
and ( n871 , n782 , n288 );
xor ( n872 , n870 , n871 );
and ( n873 , n743 , n756 );
and ( n874 , n756 , n771 );
and ( n875 , n743 , n771 );
or ( n876 , n873 , n874 , n875 );
and ( n877 , n759 , n764 );
and ( n878 , n764 , n770 );
and ( n879 , n759 , n770 );
or ( n880 , n877 , n878 , n879 );
and ( n881 , n750 , n751 );
and ( n882 , n751 , n754 );
and ( n883 , n750 , n754 );
or ( n884 , n881 , n882 , n883 );
and ( n885 , n760 , n761 );
and ( n886 , n761 , n763 );
and ( n887 , n760 , n763 );
or ( n888 , n885 , n886 , n887 );
xor ( n889 , n884 , n888 );
and ( n890 , n521 , n354 );
and ( n891 , n625 , n321 );
xor ( n892 , n890 , n891 );
and ( n893 , n753 , n291 );
xor ( n894 , n892 , n893 );
xor ( n895 , n889 , n894 );
xor ( n896 , n880 , n895 );
and ( n897 , n767 , n769 );
buf ( n898 , n897 );
and ( n899 , n318 , n607 );
and ( n900 , n361 , n510 );
xor ( n901 , n899 , n900 );
and ( n902 , n431 , n435 );
xor ( n903 , n901 , n902 );
xor ( n904 , n898 , n903 );
buf ( n905 , n248 );
and ( n906 , n273 , n905 );
buf ( n907 , n906 );
and ( n908 , n294 , n766 );
xor ( n909 , n907 , n908 );
xor ( n910 , n904 , n909 );
xor ( n911 , n896 , n910 );
xor ( n912 , n876 , n911 );
and ( n913 , n747 , n748 );
and ( n914 , n748 , n755 );
and ( n915 , n747 , n755 );
or ( n916 , n913 , n914 , n915 );
buf ( n917 , n217 );
and ( n918 , n917 , n274 );
xor ( n919 , n916 , n918 );
xor ( n920 , n912 , n919 );
and ( n921 , n734 , n738 );
and ( n922 , n738 , n772 );
and ( n923 , n734 , n772 );
or ( n924 , n921 , n922 , n923 );
xor ( n925 , n920 , n924 );
and ( n926 , n773 , n777 );
and ( n927 , n778 , n779 );
or ( n928 , n926 , n927 );
xor ( n929 , n925 , n928 );
buf ( n930 , n929 );
buf ( n931 , n930 );
and ( n932 , n931 , n279 );
xor ( n933 , n872 , n932 );
xor ( n934 , n869 , n933 );
xor ( n935 , n859 , n934 );
xor ( n936 , n840 , n935 );
and ( n937 , n712 , n718 );
buf ( n938 , n937 );
buf ( n939 , n938 );
xor ( n940 , n936 , n939 );
and ( n941 , n699 , n703 );
and ( n942 , n703 , n786 );
and ( n943 , n699 , n786 );
or ( n944 , n941 , n942 , n943 );
xor ( n945 , n940 , n944 );
and ( n946 , n787 , n789 );
and ( n947 , n790 , n791 );
or ( n948 , n946 , n947 );
xor ( n949 , n945 , n948 );
buf ( n950 , n949 );
buf ( n951 , n950 );
not ( n952 , n951 );
buf ( n953 , n203 );
not ( n954 , n953 );
nor ( n955 , n952 , n954 );
xor ( n956 , n836 , n955 );
xor ( n957 , n803 , n833 );
nor ( n958 , n795 , n954 );
and ( n959 , n957 , n958 );
xor ( n960 , n957 , n958 );
xor ( n961 , n807 , n831 );
nor ( n962 , n663 , n954 );
and ( n963 , n961 , n962 );
xor ( n964 , n961 , n962 );
xor ( n965 , n811 , n829 );
nor ( n966 , n549 , n954 );
and ( n967 , n965 , n966 );
xor ( n968 , n965 , n966 );
xor ( n969 , n815 , n827 );
nor ( n970 , n456 , n954 );
and ( n971 , n969 , n970 );
xor ( n972 , n969 , n970 );
xor ( n973 , n820 , n825 );
nor ( n974 , n384 , n954 );
and ( n975 , n973 , n974 );
xor ( n976 , n973 , n974 );
xor ( n977 , n822 , n823 );
buf ( n978 , n977 );
nor ( n979 , n334 , n954 );
and ( n980 , n978 , n979 );
xor ( n981 , n978 , n979 );
nor ( n982 , n283 , n797 );
buf ( n983 , n982 );
nor ( n984 , n303 , n954 );
and ( n985 , n983 , n984 );
buf ( n986 , n985 );
and ( n987 , n981 , n986 );
or ( n988 , n980 , n987 );
and ( n989 , n976 , n988 );
or ( n990 , n975 , n989 );
and ( n991 , n972 , n990 );
or ( n992 , n971 , n991 );
and ( n993 , n968 , n992 );
or ( n994 , n967 , n993 );
and ( n995 , n964 , n994 );
or ( n996 , n963 , n995 );
and ( n997 , n960 , n996 );
or ( n998 , n959 , n997 );
xor ( n999 , n956 , n998 );
and ( n1000 , n840 , n935 );
and ( n1001 , n935 , n939 );
and ( n1002 , n840 , n939 );
or ( n1003 , n1000 , n1001 , n1002 );
buf ( n1004 , n1003 );
and ( n1005 , n844 , n858 );
and ( n1006 , n858 , n934 );
and ( n1007 , n844 , n934 );
or ( n1008 , n1005 , n1006 , n1007 );
and ( n1009 , n863 , n868 );
and ( n1010 , n868 , n933 );
and ( n1011 , n863 , n933 );
or ( n1012 , n1009 , n1010 , n1011 );
and ( n1013 , n870 , n871 );
and ( n1014 , n871 , n932 );
and ( n1015 , n870 , n932 );
or ( n1016 , n1013 , n1014 , n1015 );
and ( n1017 , n446 , n488 );
and ( n1018 , n533 , n411 );
xor ( n1019 , n1017 , n1018 );
and ( n1020 , n636 , n375 );
xor ( n1021 , n1019 , n1020 );
xor ( n1022 , n1016 , n1021 );
and ( n1023 , n782 , n312 );
and ( n1024 , n931 , n288 );
xor ( n1025 , n1023 , n1024 );
and ( n1026 , n916 , n918 );
and ( n1027 , n876 , n911 );
and ( n1028 , n911 , n919 );
and ( n1029 , n876 , n919 );
or ( n1030 , n1027 , n1028 , n1029 );
xor ( n1031 , n1026 , n1030 );
and ( n1032 , n880 , n895 );
and ( n1033 , n895 , n910 );
and ( n1034 , n880 , n910 );
or ( n1035 , n1032 , n1033 , n1034 );
and ( n1036 , n898 , n903 );
and ( n1037 , n903 , n909 );
and ( n1038 , n898 , n909 );
or ( n1039 , n1036 , n1037 , n1038 );
and ( n1040 , n906 , n908 );
buf ( n1041 , n1040 );
and ( n1042 , n318 , n766 );
and ( n1043 , n361 , n607 );
xor ( n1044 , n1042 , n1043 );
and ( n1045 , n431 , n510 );
xor ( n1046 , n1044 , n1045 );
xor ( n1047 , n1041 , n1046 );
buf ( n1048 , n247 );
and ( n1049 , n273 , n1048 );
buf ( n1050 , n1049 );
and ( n1051 , n294 , n905 );
xor ( n1052 , n1050 , n1051 );
xor ( n1053 , n1047 , n1052 );
xor ( n1054 , n1039 , n1053 );
and ( n1055 , n890 , n891 );
and ( n1056 , n891 , n893 );
and ( n1057 , n890 , n893 );
or ( n1058 , n1055 , n1056 , n1057 );
and ( n1059 , n899 , n900 );
and ( n1060 , n900 , n902 );
and ( n1061 , n899 , n902 );
or ( n1062 , n1059 , n1060 , n1061 );
xor ( n1063 , n1058 , n1062 );
and ( n1064 , n521 , n435 );
and ( n1065 , n625 , n354 );
xor ( n1066 , n1064 , n1065 );
and ( n1067 , n753 , n321 );
xor ( n1068 , n1066 , n1067 );
xor ( n1069 , n1063 , n1068 );
xor ( n1070 , n1054 , n1069 );
xor ( n1071 , n1035 , n1070 );
and ( n1072 , n884 , n888 );
and ( n1073 , n888 , n894 );
and ( n1074 , n884 , n894 );
or ( n1075 , n1072 , n1073 , n1074 );
and ( n1076 , n917 , n291 );
buf ( n1077 , n216 );
and ( n1078 , n1077 , n274 );
xor ( n1079 , n1076 , n1078 );
xor ( n1080 , n1075 , n1079 );
xor ( n1081 , n1071 , n1080 );
xor ( n1082 , n1031 , n1081 );
and ( n1083 , n920 , n924 );
and ( n1084 , n925 , n928 );
or ( n1085 , n1083 , n1084 );
xor ( n1086 , n1082 , n1085 );
buf ( n1087 , n1086 );
buf ( n1088 , n1087 );
and ( n1089 , n1088 , n279 );
xor ( n1090 , n1025 , n1089 );
xor ( n1091 , n1022 , n1090 );
xor ( n1092 , n1012 , n1091 );
and ( n1093 , n853 , n854 );
and ( n1094 , n854 , n856 );
and ( n1095 , n853 , n856 );
or ( n1096 , n1093 , n1094 , n1095 );
and ( n1097 , n864 , n865 );
and ( n1098 , n865 , n867 );
and ( n1099 , n864 , n867 );
or ( n1100 , n1097 , n1098 , n1099 );
xor ( n1101 , n1096 , n1100 );
and ( n1102 , n298 , n852 );
and ( n1103 , n328 , n714 );
xor ( n1104 , n1102 , n1103 );
and ( n1105 , n371 , n651 );
xor ( n1106 , n1104 , n1105 );
xor ( n1107 , n1101 , n1106 );
xor ( n1108 , n1092 , n1107 );
xor ( n1109 , n1008 , n1108 );
and ( n1110 , n846 , n850 );
and ( n1111 , n850 , n857 );
and ( n1112 , n846 , n857 );
or ( n1113 , n1110 , n1111 , n1112 );
buf ( n1114 , n232 );
and ( n1115 , n277 , n1114 );
buf ( n1116 , n1115 );
xor ( n1117 , n1113 , n1116 );
xor ( n1118 , n1109 , n1117 );
xor ( n1119 , n1004 , n1118 );
and ( n1120 , n940 , n944 );
and ( n1121 , n945 , n948 );
or ( n1122 , n1120 , n1121 );
xor ( n1123 , n1119 , n1122 );
buf ( n1124 , n1123 );
buf ( n1125 , n1124 );
not ( n1126 , n1125 );
buf ( n1127 , n204 );
not ( n1128 , n1127 );
nor ( n1129 , n1126 , n1128 );
xor ( n1130 , n999 , n1129 );
xor ( n1131 , n960 , n996 );
nor ( n1132 , n952 , n1128 );
and ( n1133 , n1131 , n1132 );
xor ( n1134 , n1131 , n1132 );
xor ( n1135 , n964 , n994 );
nor ( n1136 , n795 , n1128 );
and ( n1137 , n1135 , n1136 );
xor ( n1138 , n1135 , n1136 );
xor ( n1139 , n968 , n992 );
nor ( n1140 , n663 , n1128 );
and ( n1141 , n1139 , n1140 );
xor ( n1142 , n1139 , n1140 );
xor ( n1143 , n972 , n990 );
nor ( n1144 , n549 , n1128 );
and ( n1145 , n1143 , n1144 );
xor ( n1146 , n1143 , n1144 );
xor ( n1147 , n976 , n988 );
nor ( n1148 , n456 , n1128 );
and ( n1149 , n1147 , n1148 );
xor ( n1150 , n1147 , n1148 );
xor ( n1151 , n981 , n986 );
nor ( n1152 , n384 , n1128 );
and ( n1153 , n1151 , n1152 );
xor ( n1154 , n1151 , n1152 );
xor ( n1155 , n983 , n984 );
buf ( n1156 , n1155 );
nor ( n1157 , n334 , n1128 );
and ( n1158 , n1156 , n1157 );
xor ( n1159 , n1156 , n1157 );
nor ( n1160 , n283 , n954 );
buf ( n1161 , n1160 );
nor ( n1162 , n303 , n1128 );
and ( n1163 , n1161 , n1162 );
buf ( n1164 , n1163 );
and ( n1165 , n1159 , n1164 );
or ( n1166 , n1158 , n1165 );
and ( n1167 , n1154 , n1166 );
or ( n1168 , n1153 , n1167 );
and ( n1169 , n1150 , n1168 );
or ( n1170 , n1149 , n1169 );
and ( n1171 , n1146 , n1170 );
or ( n1172 , n1145 , n1171 );
and ( n1173 , n1142 , n1172 );
or ( n1174 , n1141 , n1173 );
and ( n1175 , n1138 , n1174 );
or ( n1176 , n1137 , n1175 );
and ( n1177 , n1134 , n1176 );
or ( n1178 , n1133 , n1177 );
xor ( n1179 , n1130 , n1178 );
and ( n1180 , n1113 , n1116 );
and ( n1181 , n1008 , n1108 );
and ( n1182 , n1108 , n1117 );
and ( n1183 , n1008 , n1117 );
or ( n1184 , n1181 , n1182 , n1183 );
xor ( n1185 , n1180 , n1184 );
and ( n1186 , n1012 , n1091 );
and ( n1187 , n1091 , n1107 );
and ( n1188 , n1012 , n1107 );
or ( n1189 , n1186 , n1187 , n1188 );
and ( n1190 , n1016 , n1021 );
and ( n1191 , n1021 , n1090 );
and ( n1192 , n1016 , n1090 );
or ( n1193 , n1190 , n1191 , n1192 );
and ( n1194 , n1017 , n1018 );
and ( n1195 , n1018 , n1020 );
and ( n1196 , n1017 , n1020 );
or ( n1197 , n1194 , n1195 , n1196 );
and ( n1198 , n1102 , n1103 );
and ( n1199 , n1103 , n1105 );
and ( n1200 , n1102 , n1105 );
or ( n1201 , n1198 , n1199 , n1200 );
xor ( n1202 , n1197 , n1201 );
and ( n1203 , n328 , n852 );
and ( n1204 , n371 , n714 );
xor ( n1205 , n1203 , n1204 );
and ( n1206 , n446 , n651 );
xor ( n1207 , n1205 , n1206 );
xor ( n1208 , n1202 , n1207 );
xor ( n1209 , n1193 , n1208 );
and ( n1210 , n1023 , n1024 );
and ( n1211 , n1024 , n1089 );
and ( n1212 , n1023 , n1089 );
or ( n1213 , n1210 , n1211 , n1212 );
and ( n1214 , n533 , n488 );
and ( n1215 , n636 , n411 );
xor ( n1216 , n1214 , n1215 );
and ( n1217 , n782 , n375 );
xor ( n1218 , n1216 , n1217 );
xor ( n1219 , n1213 , n1218 );
and ( n1220 , n931 , n312 );
and ( n1221 , n1088 , n288 );
xor ( n1222 , n1220 , n1221 );
and ( n1223 , n1075 , n1079 );
and ( n1224 , n1035 , n1070 );
and ( n1225 , n1070 , n1080 );
and ( n1226 , n1035 , n1080 );
or ( n1227 , n1224 , n1225 , n1226 );
xor ( n1228 , n1223 , n1227 );
and ( n1229 , n1039 , n1053 );
and ( n1230 , n1053 , n1069 );
and ( n1231 , n1039 , n1069 );
or ( n1232 , n1229 , n1230 , n1231 );
and ( n1233 , n1041 , n1046 );
and ( n1234 , n1046 , n1052 );
and ( n1235 , n1041 , n1052 );
or ( n1236 , n1233 , n1234 , n1235 );
and ( n1237 , n1042 , n1043 );
and ( n1238 , n1043 , n1045 );
and ( n1239 , n1042 , n1045 );
or ( n1240 , n1237 , n1238 , n1239 );
and ( n1241 , n1064 , n1065 );
and ( n1242 , n1065 , n1067 );
and ( n1243 , n1064 , n1067 );
or ( n1244 , n1241 , n1242 , n1243 );
xor ( n1245 , n1240 , n1244 );
and ( n1246 , n521 , n510 );
and ( n1247 , n625 , n435 );
xor ( n1248 , n1246 , n1247 );
and ( n1249 , n753 , n354 );
xor ( n1250 , n1248 , n1249 );
xor ( n1251 , n1245 , n1250 );
xor ( n1252 , n1236 , n1251 );
and ( n1253 , n1049 , n1051 );
buf ( n1254 , n1253 );
and ( n1255 , n318 , n905 );
and ( n1256 , n361 , n766 );
xor ( n1257 , n1255 , n1256 );
and ( n1258 , n431 , n607 );
xor ( n1259 , n1257 , n1258 );
xor ( n1260 , n1254 , n1259 );
buf ( n1261 , n246 );
and ( n1262 , n273 , n1261 );
buf ( n1263 , n1262 );
and ( n1264 , n294 , n1048 );
xor ( n1265 , n1263 , n1264 );
xor ( n1266 , n1260 , n1265 );
xor ( n1267 , n1252 , n1266 );
xor ( n1268 , n1232 , n1267 );
and ( n1269 , n1058 , n1062 );
and ( n1270 , n1062 , n1068 );
and ( n1271 , n1058 , n1068 );
or ( n1272 , n1269 , n1270 , n1271 );
and ( n1273 , n1076 , n1078 );
and ( n1274 , n917 , n321 );
and ( n1275 , n1077 , n291 );
xor ( n1276 , n1274 , n1275 );
buf ( n1277 , n215 );
and ( n1278 , n1277 , n274 );
xor ( n1279 , n1276 , n1278 );
xor ( n1280 , n1273 , n1279 );
xor ( n1281 , n1272 , n1280 );
xor ( n1282 , n1268 , n1281 );
xor ( n1283 , n1228 , n1282 );
and ( n1284 , n1026 , n1030 );
and ( n1285 , n1030 , n1081 );
and ( n1286 , n1026 , n1081 );
or ( n1287 , n1284 , n1285 , n1286 );
xor ( n1288 , n1283 , n1287 );
and ( n1289 , n1082 , n1085 );
xor ( n1290 , n1288 , n1289 );
buf ( n1291 , n1290 );
buf ( n1292 , n1291 );
and ( n1293 , n1292 , n279 );
xor ( n1294 , n1222 , n1293 );
xor ( n1295 , n1219 , n1294 );
xor ( n1296 , n1209 , n1295 );
xor ( n1297 , n1189 , n1296 );
and ( n1298 , n1096 , n1100 );
and ( n1299 , n1100 , n1106 );
and ( n1300 , n1096 , n1106 );
or ( n1301 , n1298 , n1299 , n1300 );
buf ( n1302 , n231 );
and ( n1303 , n277 , n1302 );
buf ( n1304 , n1303 );
and ( n1305 , n298 , n1114 );
xor ( n1306 , n1304 , n1305 );
buf ( n1307 , n1306 );
xor ( n1308 , n1301 , n1307 );
xor ( n1309 , n1297 , n1308 );
xor ( n1310 , n1185 , n1309 );
and ( n1311 , n1003 , n1118 );
buf ( n1312 , n1311 );
xor ( n1313 , n1310 , n1312 );
and ( n1314 , n1119 , n1122 );
xor ( n1315 , n1313 , n1314 );
buf ( n1316 , n1315 );
buf ( n1317 , n1316 );
not ( n1318 , n1317 );
buf ( n1319 , n205 );
not ( n1320 , n1319 );
nor ( n1321 , n1318 , n1320 );
xor ( n1322 , n1179 , n1321 );
xor ( n1323 , n1134 , n1176 );
nor ( n1324 , n1126 , n1320 );
and ( n1325 , n1323 , n1324 );
xor ( n1326 , n1323 , n1324 );
xor ( n1327 , n1138 , n1174 );
nor ( n1328 , n952 , n1320 );
and ( n1329 , n1327 , n1328 );
xor ( n1330 , n1327 , n1328 );
xor ( n1331 , n1142 , n1172 );
nor ( n1332 , n795 , n1320 );
and ( n1333 , n1331 , n1332 );
xor ( n1334 , n1331 , n1332 );
xor ( n1335 , n1146 , n1170 );
nor ( n1336 , n663 , n1320 );
and ( n1337 , n1335 , n1336 );
xor ( n1338 , n1335 , n1336 );
xor ( n1339 , n1150 , n1168 );
nor ( n1340 , n549 , n1320 );
and ( n1341 , n1339 , n1340 );
xor ( n1342 , n1339 , n1340 );
xor ( n1343 , n1154 , n1166 );
nor ( n1344 , n456 , n1320 );
and ( n1345 , n1343 , n1344 );
xor ( n1346 , n1343 , n1344 );
xor ( n1347 , n1159 , n1164 );
nor ( n1348 , n384 , n1320 );
and ( n1349 , n1347 , n1348 );
xor ( n1350 , n1347 , n1348 );
xor ( n1351 , n1161 , n1162 );
buf ( n1352 , n1351 );
nor ( n1353 , n334 , n1320 );
and ( n1354 , n1352 , n1353 );
xor ( n1355 , n1352 , n1353 );
nor ( n1356 , n283 , n1128 );
buf ( n1357 , n1356 );
nor ( n1358 , n303 , n1320 );
and ( n1359 , n1357 , n1358 );
buf ( n1360 , n1359 );
and ( n1361 , n1355 , n1360 );
or ( n1362 , n1354 , n1361 );
and ( n1363 , n1350 , n1362 );
or ( n1364 , n1349 , n1363 );
and ( n1365 , n1346 , n1364 );
or ( n1366 , n1345 , n1365 );
and ( n1367 , n1342 , n1366 );
or ( n1368 , n1341 , n1367 );
and ( n1369 , n1338 , n1368 );
or ( n1370 , n1337 , n1369 );
and ( n1371 , n1334 , n1370 );
or ( n1372 , n1333 , n1371 );
and ( n1373 , n1330 , n1372 );
or ( n1374 , n1329 , n1373 );
and ( n1375 , n1326 , n1374 );
or ( n1376 , n1325 , n1375 );
xor ( n1377 , n1322 , n1376 );
and ( n1378 , n1301 , n1307 );
and ( n1379 , n1189 , n1296 );
and ( n1380 , n1296 , n1308 );
and ( n1381 , n1189 , n1308 );
or ( n1382 , n1379 , n1380 , n1381 );
xor ( n1383 , n1378 , n1382 );
and ( n1384 , n1193 , n1208 );
and ( n1385 , n1208 , n1295 );
and ( n1386 , n1193 , n1295 );
or ( n1387 , n1384 , n1385 , n1386 );
and ( n1388 , n1197 , n1201 );
and ( n1389 , n1201 , n1207 );
and ( n1390 , n1197 , n1207 );
or ( n1391 , n1388 , n1389 , n1390 );
buf ( n1392 , n1391 );
and ( n1393 , n1303 , n1305 );
buf ( n1394 , n1393 );
buf ( n1395 , n1394 );
buf ( n1396 , n230 );
and ( n1397 , n277 , n1396 );
and ( n1398 , n298 , n1302 );
xor ( n1399 , n1397 , n1398 );
and ( n1400 , n328 , n1114 );
xor ( n1401 , n1399 , n1400 );
xor ( n1402 , n1395 , n1401 );
xor ( n1403 , n1392 , n1402 );
xor ( n1404 , n1387 , n1403 );
and ( n1405 , n1213 , n1218 );
and ( n1406 , n1218 , n1294 );
and ( n1407 , n1213 , n1294 );
or ( n1408 , n1405 , n1406 , n1407 );
and ( n1409 , n1203 , n1204 );
and ( n1410 , n1204 , n1206 );
and ( n1411 , n1203 , n1206 );
or ( n1412 , n1409 , n1410 , n1411 );
and ( n1413 , n1214 , n1215 );
and ( n1414 , n1215 , n1217 );
and ( n1415 , n1214 , n1217 );
or ( n1416 , n1413 , n1414 , n1415 );
xor ( n1417 , n1412 , n1416 );
and ( n1418 , n371 , n852 );
and ( n1419 , n446 , n714 );
xor ( n1420 , n1418 , n1419 );
and ( n1421 , n533 , n651 );
xor ( n1422 , n1420 , n1421 );
xor ( n1423 , n1417 , n1422 );
xor ( n1424 , n1408 , n1423 );
and ( n1425 , n1220 , n1221 );
and ( n1426 , n1221 , n1293 );
and ( n1427 , n1220 , n1293 );
or ( n1428 , n1425 , n1426 , n1427 );
and ( n1429 , n636 , n488 );
and ( n1430 , n782 , n411 );
xor ( n1431 , n1429 , n1430 );
and ( n1432 , n931 , n375 );
xor ( n1433 , n1431 , n1432 );
xor ( n1434 , n1428 , n1433 );
and ( n1435 , n1088 , n312 );
and ( n1436 , n1292 , n288 );
xor ( n1437 , n1435 , n1436 );
and ( n1438 , n1272 , n1280 );
and ( n1439 , n1232 , n1267 );
and ( n1440 , n1267 , n1281 );
and ( n1441 , n1232 , n1281 );
or ( n1442 , n1439 , n1440 , n1441 );
xor ( n1443 , n1438 , n1442 );
and ( n1444 , n1236 , n1251 );
and ( n1445 , n1251 , n1266 );
and ( n1446 , n1236 , n1266 );
or ( n1447 , n1444 , n1445 , n1446 );
and ( n1448 , n1240 , n1244 );
and ( n1449 , n1244 , n1250 );
and ( n1450 , n1240 , n1250 );
or ( n1451 , n1448 , n1449 , n1450 );
and ( n1452 , n1273 , n1279 );
xor ( n1453 , n1451 , n1452 );
and ( n1454 , n1274 , n1275 );
and ( n1455 , n1275 , n1278 );
and ( n1456 , n1274 , n1278 );
or ( n1457 , n1454 , n1455 , n1456 );
buf ( n1458 , n214 );
and ( n1459 , n1458 , n274 );
xor ( n1460 , n1457 , n1459 );
and ( n1461 , n917 , n354 );
and ( n1462 , n1077 , n321 );
xor ( n1463 , n1461 , n1462 );
and ( n1464 , n1277 , n291 );
xor ( n1465 , n1463 , n1464 );
xor ( n1466 , n1460 , n1465 );
xor ( n1467 , n1453 , n1466 );
xor ( n1468 , n1447 , n1467 );
and ( n1469 , n1254 , n1259 );
and ( n1470 , n1259 , n1265 );
and ( n1471 , n1254 , n1265 );
or ( n1472 , n1469 , n1470 , n1471 );
and ( n1473 , n1246 , n1247 );
and ( n1474 , n1247 , n1249 );
and ( n1475 , n1246 , n1249 );
or ( n1476 , n1473 , n1474 , n1475 );
and ( n1477 , n1255 , n1256 );
and ( n1478 , n1256 , n1258 );
and ( n1479 , n1255 , n1258 );
or ( n1480 , n1477 , n1478 , n1479 );
xor ( n1481 , n1476 , n1480 );
and ( n1482 , n521 , n607 );
and ( n1483 , n625 , n510 );
xor ( n1484 , n1482 , n1483 );
and ( n1485 , n753 , n435 );
xor ( n1486 , n1484 , n1485 );
xor ( n1487 , n1481 , n1486 );
xor ( n1488 , n1472 , n1487 );
and ( n1489 , n1262 , n1264 );
buf ( n1490 , n1489 );
and ( n1491 , n318 , n1048 );
and ( n1492 , n361 , n905 );
xor ( n1493 , n1491 , n1492 );
and ( n1494 , n431 , n766 );
xor ( n1495 , n1493 , n1494 );
xor ( n1496 , n1490 , n1495 );
buf ( n1497 , n245 );
and ( n1498 , n273 , n1497 );
buf ( n1499 , n1498 );
and ( n1500 , n294 , n1261 );
xor ( n1501 , n1499 , n1500 );
xor ( n1502 , n1496 , n1501 );
xor ( n1503 , n1488 , n1502 );
xor ( n1504 , n1468 , n1503 );
xor ( n1505 , n1443 , n1504 );
and ( n1506 , n1223 , n1227 );
and ( n1507 , n1227 , n1282 );
and ( n1508 , n1223 , n1282 );
or ( n1509 , n1506 , n1507 , n1508 );
xor ( n1510 , n1505 , n1509 );
and ( n1511 , n1283 , n1287 );
and ( n1512 , n1288 , n1289 );
or ( n1513 , n1511 , n1512 );
xor ( n1514 , n1510 , n1513 );
buf ( n1515 , n1514 );
buf ( n1516 , n1515 );
and ( n1517 , n1516 , n279 );
xor ( n1518 , n1437 , n1517 );
xor ( n1519 , n1434 , n1518 );
xor ( n1520 , n1424 , n1519 );
xor ( n1521 , n1404 , n1520 );
xor ( n1522 , n1383 , n1521 );
and ( n1523 , n1180 , n1184 );
and ( n1524 , n1184 , n1309 );
and ( n1525 , n1180 , n1309 );
or ( n1526 , n1523 , n1524 , n1525 );
xor ( n1527 , n1522 , n1526 );
and ( n1528 , n1310 , n1312 );
and ( n1529 , n1313 , n1314 );
or ( n1530 , n1528 , n1529 );
xor ( n1531 , n1527 , n1530 );
buf ( n1532 , n1531 );
buf ( n1533 , n1532 );
not ( n1534 , n1533 );
buf ( n1535 , n206 );
not ( n1536 , n1535 );
nor ( n1537 , n1534 , n1536 );
xor ( n1538 , n1377 , n1537 );
xor ( n1539 , n1326 , n1374 );
nor ( n1540 , n1318 , n1536 );
and ( n1541 , n1539 , n1540 );
xor ( n1542 , n1539 , n1540 );
xor ( n1543 , n1330 , n1372 );
nor ( n1544 , n1126 , n1536 );
and ( n1545 , n1543 , n1544 );
xor ( n1546 , n1543 , n1544 );
xor ( n1547 , n1334 , n1370 );
nor ( n1548 , n952 , n1536 );
and ( n1549 , n1547 , n1548 );
xor ( n1550 , n1547 , n1548 );
xor ( n1551 , n1338 , n1368 );
nor ( n1552 , n795 , n1536 );
and ( n1553 , n1551 , n1552 );
xor ( n1554 , n1551 , n1552 );
xor ( n1555 , n1342 , n1366 );
nor ( n1556 , n663 , n1536 );
and ( n1557 , n1555 , n1556 );
xor ( n1558 , n1555 , n1556 );
xor ( n1559 , n1346 , n1364 );
nor ( n1560 , n549 , n1536 );
and ( n1561 , n1559 , n1560 );
xor ( n1562 , n1559 , n1560 );
xor ( n1563 , n1350 , n1362 );
nor ( n1564 , n456 , n1536 );
and ( n1565 , n1563 , n1564 );
xor ( n1566 , n1563 , n1564 );
xor ( n1567 , n1355 , n1360 );
nor ( n1568 , n384 , n1536 );
and ( n1569 , n1567 , n1568 );
xor ( n1570 , n1567 , n1568 );
xor ( n1571 , n1357 , n1358 );
buf ( n1572 , n1571 );
nor ( n1573 , n334 , n1536 );
and ( n1574 , n1572 , n1573 );
xor ( n1575 , n1572 , n1573 );
nor ( n1576 , n283 , n1320 );
buf ( n1577 , n1576 );
nor ( n1578 , n303 , n1536 );
and ( n1579 , n1577 , n1578 );
buf ( n1580 , n1579 );
and ( n1581 , n1575 , n1580 );
or ( n1582 , n1574 , n1581 );
and ( n1583 , n1570 , n1582 );
or ( n1584 , n1569 , n1583 );
and ( n1585 , n1566 , n1584 );
or ( n1586 , n1565 , n1585 );
and ( n1587 , n1562 , n1586 );
or ( n1588 , n1561 , n1587 );
and ( n1589 , n1558 , n1588 );
or ( n1590 , n1557 , n1589 );
and ( n1591 , n1554 , n1590 );
or ( n1592 , n1553 , n1591 );
and ( n1593 , n1550 , n1592 );
or ( n1594 , n1549 , n1593 );
and ( n1595 , n1546 , n1594 );
or ( n1596 , n1545 , n1595 );
and ( n1597 , n1542 , n1596 );
or ( n1598 , n1541 , n1597 );
xor ( n1599 , n1538 , n1598 );
and ( n1600 , n1391 , n1402 );
buf ( n1601 , n1600 );
and ( n1602 , n1387 , n1403 );
and ( n1603 , n1403 , n1520 );
and ( n1604 , n1387 , n1520 );
or ( n1605 , n1602 , n1603 , n1604 );
xor ( n1606 , n1601 , n1605 );
and ( n1607 , n1408 , n1423 );
and ( n1608 , n1423 , n1519 );
and ( n1609 , n1408 , n1519 );
or ( n1610 , n1607 , n1608 , n1609 );
and ( n1611 , n1428 , n1433 );
and ( n1612 , n1433 , n1518 );
and ( n1613 , n1428 , n1518 );
or ( n1614 , n1611 , n1612 , n1613 );
and ( n1615 , n1418 , n1419 );
and ( n1616 , n1419 , n1421 );
and ( n1617 , n1418 , n1421 );
or ( n1618 , n1615 , n1616 , n1617 );
and ( n1619 , n1429 , n1430 );
and ( n1620 , n1430 , n1432 );
and ( n1621 , n1429 , n1432 );
or ( n1622 , n1619 , n1620 , n1621 );
xor ( n1623 , n1618 , n1622 );
and ( n1624 , n446 , n852 );
and ( n1625 , n533 , n714 );
xor ( n1626 , n1624 , n1625 );
and ( n1627 , n636 , n651 );
xor ( n1628 , n1626 , n1627 );
xor ( n1629 , n1623 , n1628 );
xor ( n1630 , n1614 , n1629 );
and ( n1631 , n1435 , n1436 );
and ( n1632 , n1436 , n1517 );
and ( n1633 , n1435 , n1517 );
or ( n1634 , n1631 , n1632 , n1633 );
and ( n1635 , n782 , n488 );
and ( n1636 , n931 , n411 );
xor ( n1637 , n1635 , n1636 );
and ( n1638 , n1088 , n375 );
xor ( n1639 , n1637 , n1638 );
xor ( n1640 , n1634 , n1639 );
and ( n1641 , n1292 , n312 );
and ( n1642 , n1516 , n288 );
xor ( n1643 , n1641 , n1642 );
and ( n1644 , n1451 , n1452 );
and ( n1645 , n1452 , n1466 );
and ( n1646 , n1451 , n1466 );
or ( n1647 , n1644 , n1645 , n1646 );
and ( n1648 , n1447 , n1467 );
and ( n1649 , n1467 , n1503 );
and ( n1650 , n1447 , n1503 );
or ( n1651 , n1648 , n1649 , n1650 );
xor ( n1652 , n1647 , n1651 );
and ( n1653 , n1472 , n1487 );
and ( n1654 , n1487 , n1502 );
and ( n1655 , n1472 , n1502 );
or ( n1656 , n1653 , n1654 , n1655 );
and ( n1657 , n1490 , n1495 );
and ( n1658 , n1495 , n1501 );
and ( n1659 , n1490 , n1501 );
or ( n1660 , n1657 , n1658 , n1659 );
and ( n1661 , n1482 , n1483 );
and ( n1662 , n1483 , n1485 );
and ( n1663 , n1482 , n1485 );
or ( n1664 , n1661 , n1662 , n1663 );
and ( n1665 , n1491 , n1492 );
and ( n1666 , n1492 , n1494 );
and ( n1667 , n1491 , n1494 );
or ( n1668 , n1665 , n1666 , n1667 );
xor ( n1669 , n1664 , n1668 );
and ( n1670 , n521 , n766 );
and ( n1671 , n625 , n607 );
xor ( n1672 , n1670 , n1671 );
and ( n1673 , n753 , n510 );
xor ( n1674 , n1672 , n1673 );
xor ( n1675 , n1669 , n1674 );
xor ( n1676 , n1660 , n1675 );
and ( n1677 , n1498 , n1500 );
buf ( n1678 , n1677 );
and ( n1679 , n318 , n1261 );
and ( n1680 , n361 , n1048 );
xor ( n1681 , n1679 , n1680 );
and ( n1682 , n431 , n905 );
xor ( n1683 , n1681 , n1682 );
xor ( n1684 , n1678 , n1683 );
buf ( n1685 , n244 );
and ( n1686 , n273 , n1685 );
buf ( n1687 , n1686 );
and ( n1688 , n294 , n1497 );
xor ( n1689 , n1687 , n1688 );
xor ( n1690 , n1684 , n1689 );
xor ( n1691 , n1676 , n1690 );
xor ( n1692 , n1656 , n1691 );
and ( n1693 , n1457 , n1459 );
and ( n1694 , n1459 , n1465 );
and ( n1695 , n1457 , n1465 );
or ( n1696 , n1693 , n1694 , n1695 );
and ( n1697 , n1476 , n1480 );
and ( n1698 , n1480 , n1486 );
and ( n1699 , n1476 , n1486 );
or ( n1700 , n1697 , n1698 , n1699 );
xor ( n1701 , n1696 , n1700 );
and ( n1702 , n1461 , n1462 );
and ( n1703 , n1462 , n1464 );
and ( n1704 , n1461 , n1464 );
or ( n1705 , n1702 , n1703 , n1704 );
and ( n1706 , n917 , n435 );
and ( n1707 , n1077 , n354 );
xor ( n1708 , n1706 , n1707 );
and ( n1709 , n1277 , n321 );
xor ( n1710 , n1708 , n1709 );
xor ( n1711 , n1705 , n1710 );
and ( n1712 , n1458 , n291 );
buf ( n1713 , n213 );
and ( n1714 , n1713 , n274 );
xor ( n1715 , n1712 , n1714 );
xor ( n1716 , n1711 , n1715 );
xor ( n1717 , n1701 , n1716 );
xor ( n1718 , n1692 , n1717 );
xor ( n1719 , n1652 , n1718 );
and ( n1720 , n1438 , n1442 );
and ( n1721 , n1442 , n1504 );
and ( n1722 , n1438 , n1504 );
or ( n1723 , n1720 , n1721 , n1722 );
xor ( n1724 , n1719 , n1723 );
and ( n1725 , n1505 , n1509 );
and ( n1726 , n1510 , n1513 );
or ( n1727 , n1725 , n1726 );
xor ( n1728 , n1724 , n1727 );
buf ( n1729 , n1728 );
buf ( n1730 , n1729 );
and ( n1731 , n1730 , n279 );
xor ( n1732 , n1643 , n1731 );
xor ( n1733 , n1640 , n1732 );
xor ( n1734 , n1630 , n1733 );
xor ( n1735 , n1610 , n1734 );
and ( n1736 , n1394 , n1401 );
buf ( n1737 , n1736 );
and ( n1738 , n1412 , n1416 );
and ( n1739 , n1416 , n1422 );
and ( n1740 , n1412 , n1422 );
or ( n1741 , n1738 , n1739 , n1740 );
xor ( n1742 , n1737 , n1741 );
and ( n1743 , n1397 , n1398 );
and ( n1744 , n1398 , n1400 );
and ( n1745 , n1397 , n1400 );
or ( n1746 , n1743 , n1744 , n1745 );
and ( n1747 , n298 , n1396 );
and ( n1748 , n328 , n1302 );
xor ( n1749 , n1747 , n1748 );
and ( n1750 , n371 , n1114 );
xor ( n1751 , n1749 , n1750 );
xor ( n1752 , n1746 , n1751 );
buf ( n1753 , n229 );
and ( n1754 , n277 , n1753 );
buf ( n1755 , n1754 );
xor ( n1756 , n1752 , n1755 );
xor ( n1757 , n1742 , n1756 );
xor ( n1758 , n1735 , n1757 );
xor ( n1759 , n1606 , n1758 );
and ( n1760 , n1378 , n1382 );
and ( n1761 , n1382 , n1521 );
and ( n1762 , n1378 , n1521 );
or ( n1763 , n1760 , n1761 , n1762 );
xor ( n1764 , n1759 , n1763 );
and ( n1765 , n1522 , n1526 );
and ( n1766 , n1527 , n1530 );
or ( n1767 , n1765 , n1766 );
xor ( n1768 , n1764 , n1767 );
buf ( n1769 , n1768 );
buf ( n1770 , n1769 );
not ( n1771 , n1770 );
buf ( n1772 , n207 );
not ( n1773 , n1772 );
nor ( n1774 , n1771 , n1773 );
xor ( n1775 , n1599 , n1774 );
xor ( n1776 , n1542 , n1596 );
nor ( n1777 , n1534 , n1773 );
and ( n1778 , n1776 , n1777 );
xor ( n1779 , n1776 , n1777 );
xor ( n1780 , n1546 , n1594 );
nor ( n1781 , n1318 , n1773 );
and ( n1782 , n1780 , n1781 );
xor ( n1783 , n1780 , n1781 );
xor ( n1784 , n1550 , n1592 );
nor ( n1785 , n1126 , n1773 );
and ( n1786 , n1784 , n1785 );
xor ( n1787 , n1784 , n1785 );
xor ( n1788 , n1554 , n1590 );
nor ( n1789 , n952 , n1773 );
and ( n1790 , n1788 , n1789 );
xor ( n1791 , n1788 , n1789 );
xor ( n1792 , n1558 , n1588 );
nor ( n1793 , n795 , n1773 );
and ( n1794 , n1792 , n1793 );
xor ( n1795 , n1792 , n1793 );
xor ( n1796 , n1562 , n1586 );
nor ( n1797 , n663 , n1773 );
and ( n1798 , n1796 , n1797 );
xor ( n1799 , n1796 , n1797 );
xor ( n1800 , n1566 , n1584 );
nor ( n1801 , n549 , n1773 );
and ( n1802 , n1800 , n1801 );
xor ( n1803 , n1800 , n1801 );
xor ( n1804 , n1570 , n1582 );
nor ( n1805 , n456 , n1773 );
and ( n1806 , n1804 , n1805 );
xor ( n1807 , n1804 , n1805 );
xor ( n1808 , n1575 , n1580 );
nor ( n1809 , n384 , n1773 );
and ( n1810 , n1808 , n1809 );
xor ( n1811 , n1808 , n1809 );
xor ( n1812 , n1577 , n1578 );
buf ( n1813 , n1812 );
nor ( n1814 , n334 , n1773 );
and ( n1815 , n1813 , n1814 );
xor ( n1816 , n1813 , n1814 );
nor ( n1817 , n283 , n1536 );
buf ( n1818 , n1817 );
nor ( n1819 , n303 , n1773 );
and ( n1820 , n1818 , n1819 );
buf ( n1821 , n1820 );
and ( n1822 , n1816 , n1821 );
or ( n1823 , n1815 , n1822 );
and ( n1824 , n1811 , n1823 );
or ( n1825 , n1810 , n1824 );
and ( n1826 , n1807 , n1825 );
or ( n1827 , n1806 , n1826 );
and ( n1828 , n1803 , n1827 );
or ( n1829 , n1802 , n1828 );
and ( n1830 , n1799 , n1829 );
or ( n1831 , n1798 , n1830 );
and ( n1832 , n1795 , n1831 );
or ( n1833 , n1794 , n1832 );
and ( n1834 , n1791 , n1833 );
or ( n1835 , n1790 , n1834 );
and ( n1836 , n1787 , n1835 );
or ( n1837 , n1786 , n1836 );
and ( n1838 , n1783 , n1837 );
or ( n1839 , n1782 , n1838 );
and ( n1840 , n1779 , n1839 );
or ( n1841 , n1778 , n1840 );
xor ( n1842 , n1775 , n1841 );
and ( n1843 , n1610 , n1734 );
and ( n1844 , n1734 , n1757 );
and ( n1845 , n1610 , n1757 );
or ( n1846 , n1843 , n1844 , n1845 );
and ( n1847 , n1614 , n1629 );
and ( n1848 , n1629 , n1733 );
and ( n1849 , n1614 , n1733 );
or ( n1850 , n1847 , n1848 , n1849 );
and ( n1851 , n1618 , n1622 );
and ( n1852 , n1622 , n1628 );
and ( n1853 , n1618 , n1628 );
or ( n1854 , n1851 , n1852 , n1853 );
and ( n1855 , n1746 , n1751 );
and ( n1856 , n1751 , n1755 );
and ( n1857 , n1746 , n1755 );
or ( n1858 , n1855 , n1856 , n1857 );
xor ( n1859 , n1854 , n1858 );
and ( n1860 , n1747 , n1748 );
and ( n1861 , n1748 , n1750 );
and ( n1862 , n1747 , n1750 );
or ( n1863 , n1860 , n1861 , n1862 );
buf ( n1864 , n228 );
and ( n1865 , n277 , n1864 );
buf ( n1866 , n1865 );
and ( n1867 , n298 , n1753 );
xor ( n1868 , n1866 , n1867 );
xor ( n1869 , n1863 , n1868 );
and ( n1870 , n328 , n1396 );
and ( n1871 , n371 , n1302 );
xor ( n1872 , n1870 , n1871 );
and ( n1873 , n446 , n1114 );
xor ( n1874 , n1872 , n1873 );
xor ( n1875 , n1869 , n1874 );
xor ( n1876 , n1859 , n1875 );
xor ( n1877 , n1850 , n1876 );
and ( n1878 , n1634 , n1639 );
and ( n1879 , n1639 , n1732 );
and ( n1880 , n1634 , n1732 );
or ( n1881 , n1878 , n1879 , n1880 );
and ( n1882 , n1624 , n1625 );
and ( n1883 , n1625 , n1627 );
and ( n1884 , n1624 , n1627 );
or ( n1885 , n1882 , n1883 , n1884 );
and ( n1886 , n1635 , n1636 );
and ( n1887 , n1636 , n1638 );
and ( n1888 , n1635 , n1638 );
or ( n1889 , n1886 , n1887 , n1888 );
xor ( n1890 , n1885 , n1889 );
and ( n1891 , n533 , n852 );
and ( n1892 , n636 , n714 );
xor ( n1893 , n1891 , n1892 );
and ( n1894 , n782 , n651 );
xor ( n1895 , n1893 , n1894 );
xor ( n1896 , n1890 , n1895 );
xor ( n1897 , n1881 , n1896 );
and ( n1898 , n1641 , n1642 );
and ( n1899 , n1642 , n1731 );
and ( n1900 , n1641 , n1731 );
or ( n1901 , n1898 , n1899 , n1900 );
and ( n1902 , n931 , n488 );
and ( n1903 , n1088 , n411 );
xor ( n1904 , n1902 , n1903 );
and ( n1905 , n1292 , n375 );
xor ( n1906 , n1904 , n1905 );
xor ( n1907 , n1901 , n1906 );
and ( n1908 , n1516 , n312 );
and ( n1909 , n1730 , n288 );
xor ( n1910 , n1908 , n1909 );
and ( n1911 , n1656 , n1691 );
and ( n1912 , n1691 , n1717 );
and ( n1913 , n1656 , n1717 );
or ( n1914 , n1911 , n1912 , n1913 );
and ( n1915 , n1660 , n1675 );
and ( n1916 , n1675 , n1690 );
and ( n1917 , n1660 , n1690 );
or ( n1918 , n1915 , n1916 , n1917 );
and ( n1919 , n1664 , n1668 );
and ( n1920 , n1668 , n1674 );
and ( n1921 , n1664 , n1674 );
or ( n1922 , n1919 , n1920 , n1921 );
and ( n1923 , n1705 , n1710 );
and ( n1924 , n1710 , n1715 );
and ( n1925 , n1705 , n1715 );
or ( n1926 , n1923 , n1924 , n1925 );
xor ( n1927 , n1922 , n1926 );
and ( n1928 , n1706 , n1707 );
and ( n1929 , n1707 , n1709 );
and ( n1930 , n1706 , n1709 );
or ( n1931 , n1928 , n1929 , n1930 );
and ( n1932 , n1458 , n321 );
and ( n1933 , n1713 , n291 );
xor ( n1934 , n1932 , n1933 );
buf ( n1935 , n212 );
and ( n1936 , n1935 , n274 );
xor ( n1937 , n1934 , n1936 );
xor ( n1938 , n1931 , n1937 );
and ( n1939 , n917 , n510 );
and ( n1940 , n1077 , n435 );
xor ( n1941 , n1939 , n1940 );
and ( n1942 , n1277 , n354 );
xor ( n1943 , n1941 , n1942 );
xor ( n1944 , n1938 , n1943 );
xor ( n1945 , n1927 , n1944 );
xor ( n1946 , n1918 , n1945 );
and ( n1947 , n1678 , n1683 );
and ( n1948 , n1683 , n1689 );
and ( n1949 , n1678 , n1689 );
or ( n1950 , n1947 , n1948 , n1949 );
and ( n1951 , n1670 , n1671 );
and ( n1952 , n1671 , n1673 );
and ( n1953 , n1670 , n1673 );
or ( n1954 , n1951 , n1952 , n1953 );
and ( n1955 , n1679 , n1680 );
and ( n1956 , n1680 , n1682 );
and ( n1957 , n1679 , n1682 );
or ( n1958 , n1955 , n1956 , n1957 );
xor ( n1959 , n1954 , n1958 );
and ( n1960 , n521 , n905 );
and ( n1961 , n625 , n766 );
xor ( n1962 , n1960 , n1961 );
and ( n1963 , n753 , n607 );
xor ( n1964 , n1962 , n1963 );
xor ( n1965 , n1959 , n1964 );
xor ( n1966 , n1950 , n1965 );
and ( n1967 , n1686 , n1688 );
buf ( n1968 , n1967 );
and ( n1969 , n318 , n1497 );
and ( n1970 , n361 , n1261 );
xor ( n1971 , n1969 , n1970 );
and ( n1972 , n431 , n1048 );
xor ( n1973 , n1971 , n1972 );
xor ( n1974 , n1968 , n1973 );
buf ( n1975 , n243 );
and ( n1976 , n273 , n1975 );
buf ( n1977 , n1976 );
and ( n1978 , n294 , n1685 );
xor ( n1979 , n1977 , n1978 );
xor ( n1980 , n1974 , n1979 );
xor ( n1981 , n1966 , n1980 );
xor ( n1982 , n1946 , n1981 );
xor ( n1983 , n1914 , n1982 );
and ( n1984 , n1712 , n1714 );
and ( n1985 , n1696 , n1700 );
and ( n1986 , n1700 , n1716 );
and ( n1987 , n1696 , n1716 );
or ( n1988 , n1985 , n1986 , n1987 );
xor ( n1989 , n1984 , n1988 );
xor ( n1990 , n1983 , n1989 );
and ( n1991 , n1647 , n1651 );
and ( n1992 , n1651 , n1718 );
and ( n1993 , n1647 , n1718 );
or ( n1994 , n1991 , n1992 , n1993 );
xor ( n1995 , n1990 , n1994 );
and ( n1996 , n1719 , n1723 );
and ( n1997 , n1724 , n1727 );
or ( n1998 , n1996 , n1997 );
xor ( n1999 , n1995 , n1998 );
buf ( n2000 , n1999 );
buf ( n2001 , n2000 );
and ( n2002 , n2001 , n279 );
xor ( n2003 , n1910 , n2002 );
xor ( n2004 , n1907 , n2003 );
xor ( n2005 , n1897 , n2004 );
xor ( n2006 , n1877 , n2005 );
xor ( n2007 , n1846 , n2006 );
and ( n2008 , n1737 , n1741 );
and ( n2009 , n1741 , n1756 );
and ( n2010 , n1737 , n1756 );
or ( n2011 , n2008 , n2009 , n2010 );
buf ( n2012 , n2011 );
xor ( n2013 , n2007 , n2012 );
and ( n2014 , n1601 , n1605 );
and ( n2015 , n1605 , n1758 );
and ( n2016 , n1601 , n1758 );
or ( n2017 , n2014 , n2015 , n2016 );
xor ( n2018 , n2013 , n2017 );
and ( n2019 , n1759 , n1763 );
and ( n2020 , n1764 , n1767 );
or ( n2021 , n2019 , n2020 );
xor ( n2022 , n2018 , n2021 );
buf ( n2023 , n2022 );
buf ( n2024 , n2023 );
not ( n2025 , n2024 );
buf ( n2026 , n208 );
not ( n2027 , n2026 );
nor ( n2028 , n2025 , n2027 );
xor ( n2029 , n1842 , n2028 );
xor ( n2030 , n1779 , n1839 );
nor ( n2031 , n1771 , n2027 );
and ( n2032 , n2030 , n2031 );
xor ( n2033 , n2030 , n2031 );
xor ( n2034 , n1783 , n1837 );
nor ( n2035 , n1534 , n2027 );
and ( n2036 , n2034 , n2035 );
xor ( n2037 , n2034 , n2035 );
xor ( n2038 , n1787 , n1835 );
nor ( n2039 , n1318 , n2027 );
and ( n2040 , n2038 , n2039 );
xor ( n2041 , n2038 , n2039 );
xor ( n2042 , n1791 , n1833 );
nor ( n2043 , n1126 , n2027 );
and ( n2044 , n2042 , n2043 );
xor ( n2045 , n2042 , n2043 );
xor ( n2046 , n1795 , n1831 );
nor ( n2047 , n952 , n2027 );
and ( n2048 , n2046 , n2047 );
xor ( n2049 , n2046 , n2047 );
xor ( n2050 , n1799 , n1829 );
nor ( n2051 , n795 , n2027 );
and ( n2052 , n2050 , n2051 );
xor ( n2053 , n2050 , n2051 );
xor ( n2054 , n1803 , n1827 );
nor ( n2055 , n663 , n2027 );
and ( n2056 , n2054 , n2055 );
xor ( n2057 , n2054 , n2055 );
xor ( n2058 , n1807 , n1825 );
nor ( n2059 , n549 , n2027 );
and ( n2060 , n2058 , n2059 );
xor ( n2061 , n2058 , n2059 );
xor ( n2062 , n1811 , n1823 );
nor ( n2063 , n456 , n2027 );
and ( n2064 , n2062 , n2063 );
xor ( n2065 , n2062 , n2063 );
xor ( n2066 , n1816 , n1821 );
nor ( n2067 , n384 , n2027 );
and ( n2068 , n2066 , n2067 );
xor ( n2069 , n2066 , n2067 );
xor ( n2070 , n1818 , n1819 );
buf ( n2071 , n2070 );
nor ( n2072 , n334 , n2027 );
and ( n2073 , n2071 , n2072 );
xor ( n2074 , n2071 , n2072 );
nor ( n2075 , n283 , n1773 );
buf ( n2076 , n2075 );
nor ( n2077 , n303 , n2027 );
and ( n2078 , n2076 , n2077 );
buf ( n2079 , n2078 );
and ( n2080 , n2074 , n2079 );
or ( n2081 , n2073 , n2080 );
and ( n2082 , n2069 , n2081 );
or ( n2083 , n2068 , n2082 );
and ( n2084 , n2065 , n2083 );
or ( n2085 , n2064 , n2084 );
and ( n2086 , n2061 , n2085 );
or ( n2087 , n2060 , n2086 );
and ( n2088 , n2057 , n2087 );
or ( n2089 , n2056 , n2088 );
and ( n2090 , n2053 , n2089 );
or ( n2091 , n2052 , n2090 );
and ( n2092 , n2049 , n2091 );
or ( n2093 , n2048 , n2092 );
and ( n2094 , n2045 , n2093 );
or ( n2095 , n2044 , n2094 );
and ( n2096 , n2041 , n2095 );
or ( n2097 , n2040 , n2096 );
and ( n2098 , n2037 , n2097 );
or ( n2099 , n2036 , n2098 );
and ( n2100 , n2033 , n2099 );
or ( n2101 , n2032 , n2100 );
xor ( n2102 , n2029 , n2101 );
and ( n2103 , n1846 , n2006 );
and ( n2104 , n2006 , n2012 );
and ( n2105 , n1846 , n2012 );
or ( n2106 , n2103 , n2104 , n2105 );
buf ( n2107 , n2106 );
and ( n2108 , n1850 , n1876 );
and ( n2109 , n1876 , n2005 );
and ( n2110 , n1850 , n2005 );
or ( n2111 , n2108 , n2109 , n2110 );
and ( n2112 , n1865 , n1867 );
buf ( n2113 , n2112 );
and ( n2114 , n1854 , n1858 );
and ( n2115 , n1858 , n1875 );
and ( n2116 , n1854 , n1875 );
or ( n2117 , n2114 , n2115 , n2116 );
xor ( n2118 , n2113 , n2117 );
buf ( n2119 , n2118 );
xor ( n2120 , n2111 , n2119 );
and ( n2121 , n1881 , n1896 );
and ( n2122 , n1896 , n2004 );
and ( n2123 , n1881 , n2004 );
or ( n2124 , n2121 , n2122 , n2123 );
and ( n2125 , n1863 , n1868 );
and ( n2126 , n1868 , n1874 );
and ( n2127 , n1863 , n1874 );
or ( n2128 , n2125 , n2126 , n2127 );
and ( n2129 , n1885 , n1889 );
and ( n2130 , n1889 , n1895 );
and ( n2131 , n1885 , n1895 );
or ( n2132 , n2129 , n2130 , n2131 );
xor ( n2133 , n2128 , n2132 );
and ( n2134 , n1870 , n1871 );
and ( n2135 , n1871 , n1873 );
and ( n2136 , n1870 , n1873 );
or ( n2137 , n2134 , n2135 , n2136 );
buf ( n2138 , n227 );
and ( n2139 , n277 , n2138 );
and ( n2140 , n298 , n1864 );
xor ( n2141 , n2139 , n2140 );
and ( n2142 , n328 , n1753 );
xor ( n2143 , n2141 , n2142 );
xor ( n2144 , n2137 , n2143 );
and ( n2145 , n371 , n1396 );
and ( n2146 , n446 , n1302 );
xor ( n2147 , n2145 , n2146 );
and ( n2148 , n533 , n1114 );
xor ( n2149 , n2147 , n2148 );
xor ( n2150 , n2144 , n2149 );
xor ( n2151 , n2133 , n2150 );
xor ( n2152 , n2124 , n2151 );
and ( n2153 , n1901 , n1906 );
and ( n2154 , n1906 , n2003 );
and ( n2155 , n1901 , n2003 );
or ( n2156 , n2153 , n2154 , n2155 );
and ( n2157 , n1891 , n1892 );
and ( n2158 , n1892 , n1894 );
and ( n2159 , n1891 , n1894 );
or ( n2160 , n2157 , n2158 , n2159 );
and ( n2161 , n1902 , n1903 );
and ( n2162 , n1903 , n1905 );
and ( n2163 , n1902 , n1905 );
or ( n2164 , n2161 , n2162 , n2163 );
xor ( n2165 , n2160 , n2164 );
and ( n2166 , n636 , n852 );
and ( n2167 , n782 , n714 );
xor ( n2168 , n2166 , n2167 );
and ( n2169 , n931 , n651 );
xor ( n2170 , n2168 , n2169 );
xor ( n2171 , n2165 , n2170 );
xor ( n2172 , n2156 , n2171 );
and ( n2173 , n1908 , n1909 );
and ( n2174 , n1909 , n2002 );
and ( n2175 , n1908 , n2002 );
or ( n2176 , n2173 , n2174 , n2175 );
and ( n2177 , n1088 , n488 );
and ( n2178 , n1292 , n411 );
xor ( n2179 , n2177 , n2178 );
and ( n2180 , n1516 , n375 );
xor ( n2181 , n2179 , n2180 );
xor ( n2182 , n2176 , n2181 );
and ( n2183 , n1730 , n312 );
and ( n2184 , n2001 , n288 );
xor ( n2185 , n2183 , n2184 );
and ( n2186 , n1984 , n1988 );
and ( n2187 , n1914 , n1982 );
and ( n2188 , n1982 , n1989 );
and ( n2189 , n1914 , n1989 );
or ( n2190 , n2187 , n2188 , n2189 );
xor ( n2191 , n2186 , n2190 );
and ( n2192 , n1918 , n1945 );
and ( n2193 , n1945 , n1981 );
and ( n2194 , n1918 , n1981 );
or ( n2195 , n2192 , n2193 , n2194 );
and ( n2196 , n1932 , n1933 );
and ( n2197 , n1933 , n1936 );
and ( n2198 , n1932 , n1936 );
or ( n2199 , n2196 , n2197 , n2198 );
and ( n2200 , n1922 , n1926 );
and ( n2201 , n1926 , n1944 );
and ( n2202 , n1922 , n1944 );
or ( n2203 , n2200 , n2201 , n2202 );
xor ( n2204 , n2199 , n2203 );
buf ( n2205 , n211 );
not ( n2206 , n2205 );
and ( n2207 , n2206 , n274 );
not ( n2208 , n274 );
nor ( n2209 , n2207 , n2208 );
xor ( n2210 , n2204 , n2209 );
xor ( n2211 , n2195 , n2210 );
and ( n2212 , n1950 , n1965 );
and ( n2213 , n1965 , n1980 );
and ( n2214 , n1950 , n1980 );
or ( n2215 , n2212 , n2213 , n2214 );
and ( n2216 , n1931 , n1937 );
and ( n2217 , n1937 , n1943 );
and ( n2218 , n1931 , n1943 );
or ( n2219 , n2216 , n2217 , n2218 );
and ( n2220 , n1954 , n1958 );
and ( n2221 , n1958 , n1964 );
and ( n2222 , n1954 , n1964 );
or ( n2223 , n2220 , n2221 , n2222 );
xor ( n2224 , n2219 , n2223 );
and ( n2225 , n1939 , n1940 );
and ( n2226 , n1940 , n1942 );
and ( n2227 , n1939 , n1942 );
or ( n2228 , n2225 , n2226 , n2227 );
and ( n2229 , n1458 , n354 );
and ( n2230 , n1713 , n321 );
xor ( n2231 , n2229 , n2230 );
and ( n2232 , n1935 , n291 );
xor ( n2233 , n2231 , n2232 );
xor ( n2234 , n2228 , n2233 );
and ( n2235 , n917 , n607 );
and ( n2236 , n1077 , n510 );
xor ( n2237 , n2235 , n2236 );
and ( n2238 , n1277 , n435 );
xor ( n2239 , n2237 , n2238 );
xor ( n2240 , n2234 , n2239 );
xor ( n2241 , n2224 , n2240 );
xor ( n2242 , n2215 , n2241 );
and ( n2243 , n1968 , n1973 );
and ( n2244 , n1973 , n1979 );
and ( n2245 , n1968 , n1979 );
or ( n2246 , n2243 , n2244 , n2245 );
and ( n2247 , n1960 , n1961 );
and ( n2248 , n1961 , n1963 );
and ( n2249 , n1960 , n1963 );
or ( n2250 , n2247 , n2248 , n2249 );
and ( n2251 , n1969 , n1970 );
and ( n2252 , n1970 , n1972 );
and ( n2253 , n1969 , n1972 );
or ( n2254 , n2251 , n2252 , n2253 );
xor ( n2255 , n2250 , n2254 );
and ( n2256 , n521 , n1048 );
and ( n2257 , n625 , n905 );
xor ( n2258 , n2256 , n2257 );
and ( n2259 , n753 , n766 );
xor ( n2260 , n2258 , n2259 );
xor ( n2261 , n2255 , n2260 );
xor ( n2262 , n2246 , n2261 );
and ( n2263 , n1976 , n1978 );
buf ( n2264 , n2263 );
and ( n2265 , n318 , n1685 );
and ( n2266 , n361 , n1497 );
xor ( n2267 , n2265 , n2266 );
and ( n2268 , n431 , n1261 );
xor ( n2269 , n2267 , n2268 );
xor ( n2270 , n2264 , n2269 );
buf ( n2271 , n242 );
and ( n2272 , n273 , n2271 );
buf ( n2273 , n2272 );
and ( n2274 , n294 , n1975 );
xor ( n2275 , n2273 , n2274 );
xor ( n2276 , n2270 , n2275 );
xor ( n2277 , n2262 , n2276 );
xor ( n2278 , n2242 , n2277 );
xor ( n2279 , n2211 , n2278 );
xor ( n2280 , n2191 , n2279 );
and ( n2281 , n1990 , n1994 );
and ( n2282 , n1995 , n1998 );
or ( n2283 , n2281 , n2282 );
xor ( n2284 , n2280 , n2283 );
buf ( n2285 , n2284 );
buf ( n2286 , n2285 );
and ( n2287 , n2286 , n279 );
xor ( n2288 , n2185 , n2287 );
xor ( n2289 , n2182 , n2288 );
xor ( n2290 , n2172 , n2289 );
xor ( n2291 , n2152 , n2290 );
xor ( n2292 , n2120 , n2291 );
xor ( n2293 , n2107 , n2292 );
and ( n2294 , n2013 , n2017 );
and ( n2295 , n2018 , n2021 );
or ( n2296 , n2294 , n2295 );
xor ( n2297 , n2293 , n2296 );
buf ( n2298 , n2297 );
buf ( n2299 , n2298 );
not ( n2300 , n2299 );
buf ( n2301 , n209 );
not ( n2302 , n2301 );
nor ( n2303 , n2300 , n2302 );
xor ( n2304 , n2102 , n2303 );
xor ( n2305 , n2033 , n2099 );
nor ( n2306 , n2025 , n2302 );
and ( n2307 , n2305 , n2306 );
xor ( n2308 , n2305 , n2306 );
xor ( n2309 , n2037 , n2097 );
nor ( n2310 , n1771 , n2302 );
and ( n2311 , n2309 , n2310 );
xor ( n2312 , n2309 , n2310 );
xor ( n2313 , n2041 , n2095 );
nor ( n2314 , n1534 , n2302 );
and ( n2315 , n2313 , n2314 );
xor ( n2316 , n2313 , n2314 );
xor ( n2317 , n2045 , n2093 );
nor ( n2318 , n1318 , n2302 );
and ( n2319 , n2317 , n2318 );
xor ( n2320 , n2317 , n2318 );
xor ( n2321 , n2049 , n2091 );
nor ( n2322 , n1126 , n2302 );
and ( n2323 , n2321 , n2322 );
xor ( n2324 , n2321 , n2322 );
xor ( n2325 , n2053 , n2089 );
nor ( n2326 , n952 , n2302 );
and ( n2327 , n2325 , n2326 );
xor ( n2328 , n2325 , n2326 );
xor ( n2329 , n2057 , n2087 );
nor ( n2330 , n795 , n2302 );
and ( n2331 , n2329 , n2330 );
xor ( n2332 , n2329 , n2330 );
xor ( n2333 , n2061 , n2085 );
nor ( n2334 , n663 , n2302 );
and ( n2335 , n2333 , n2334 );
xor ( n2336 , n2333 , n2334 );
xor ( n2337 , n2065 , n2083 );
nor ( n2338 , n549 , n2302 );
and ( n2339 , n2337 , n2338 );
xor ( n2340 , n2337 , n2338 );
xor ( n2341 , n2069 , n2081 );
nor ( n2342 , n456 , n2302 );
and ( n2343 , n2341 , n2342 );
xor ( n2344 , n2341 , n2342 );
xor ( n2345 , n2074 , n2079 );
nor ( n2346 , n384 , n2302 );
and ( n2347 , n2345 , n2346 );
xor ( n2348 , n2345 , n2346 );
xor ( n2349 , n2076 , n2077 );
buf ( n2350 , n2349 );
nor ( n2351 , n334 , n2302 );
and ( n2352 , n2350 , n2351 );
xor ( n2353 , n2350 , n2351 );
nor ( n2354 , n283 , n2027 );
buf ( n2355 , n2354 );
nor ( n2356 , n303 , n2302 );
and ( n2357 , n2355 , n2356 );
buf ( n2358 , n2357 );
and ( n2359 , n2353 , n2358 );
or ( n2360 , n2352 , n2359 );
and ( n2361 , n2348 , n2360 );
or ( n2362 , n2347 , n2361 );
and ( n2363 , n2344 , n2362 );
or ( n2364 , n2343 , n2363 );
and ( n2365 , n2340 , n2364 );
or ( n2366 , n2339 , n2365 );
and ( n2367 , n2336 , n2366 );
or ( n2368 , n2335 , n2367 );
and ( n2369 , n2332 , n2368 );
or ( n2370 , n2331 , n2369 );
and ( n2371 , n2328 , n2370 );
or ( n2372 , n2327 , n2371 );
and ( n2373 , n2324 , n2372 );
or ( n2374 , n2323 , n2373 );
and ( n2375 , n2320 , n2374 );
or ( n2376 , n2319 , n2375 );
and ( n2377 , n2316 , n2376 );
or ( n2378 , n2315 , n2377 );
and ( n2379 , n2312 , n2378 );
or ( n2380 , n2311 , n2379 );
and ( n2381 , n2308 , n2380 );
or ( n2382 , n2307 , n2381 );
xor ( n2383 , n2304 , n2382 );
and ( n2384 , n2113 , n2117 );
buf ( n2385 , n2384 );
and ( n2386 , n2111 , n2119 );
and ( n2387 , n2119 , n2291 );
and ( n2388 , n2111 , n2291 );
or ( n2389 , n2386 , n2387 , n2388 );
xor ( n2390 , n2385 , n2389 );
and ( n2391 , n2124 , n2151 );
and ( n2392 , n2151 , n2290 );
and ( n2393 , n2124 , n2290 );
or ( n2394 , n2391 , n2392 , n2393 );
and ( n2395 , n2139 , n2140 );
and ( n2396 , n2140 , n2142 );
and ( n2397 , n2139 , n2142 );
or ( n2398 , n2395 , n2396 , n2397 );
and ( n2399 , n2128 , n2132 );
and ( n2400 , n2132 , n2150 );
and ( n2401 , n2128 , n2150 );
or ( n2402 , n2399 , n2400 , n2401 );
xor ( n2403 , n2398 , n2402 );
not ( n2404 , n277 );
buf ( n2405 , n226 );
not ( n2406 , n2405 );
and ( n2407 , n2406 , n277 );
nor ( n2408 , n2404 , n2407 );
xor ( n2409 , n2403 , n2408 );
xor ( n2410 , n2394 , n2409 );
and ( n2411 , n2156 , n2171 );
and ( n2412 , n2171 , n2289 );
and ( n2413 , n2156 , n2289 );
or ( n2414 , n2411 , n2412 , n2413 );
and ( n2415 , n2137 , n2143 );
and ( n2416 , n2143 , n2149 );
and ( n2417 , n2137 , n2149 );
or ( n2418 , n2415 , n2416 , n2417 );
and ( n2419 , n2160 , n2164 );
and ( n2420 , n2164 , n2170 );
and ( n2421 , n2160 , n2170 );
or ( n2422 , n2419 , n2420 , n2421 );
xor ( n2423 , n2418 , n2422 );
and ( n2424 , n2145 , n2146 );
and ( n2425 , n2146 , n2148 );
and ( n2426 , n2145 , n2148 );
or ( n2427 , n2424 , n2425 , n2426 );
and ( n2428 , n298 , n2138 );
and ( n2429 , n328 , n1864 );
xor ( n2430 , n2428 , n2429 );
and ( n2431 , n371 , n1753 );
xor ( n2432 , n2430 , n2431 );
xor ( n2433 , n2427 , n2432 );
and ( n2434 , n446 , n1396 );
and ( n2435 , n533 , n1302 );
xor ( n2436 , n2434 , n2435 );
and ( n2437 , n636 , n1114 );
xor ( n2438 , n2436 , n2437 );
xor ( n2439 , n2433 , n2438 );
xor ( n2440 , n2423 , n2439 );
xor ( n2441 , n2414 , n2440 );
and ( n2442 , n2176 , n2181 );
and ( n2443 , n2181 , n2288 );
and ( n2444 , n2176 , n2288 );
or ( n2445 , n2442 , n2443 , n2444 );
and ( n2446 , n2166 , n2167 );
and ( n2447 , n2167 , n2169 );
and ( n2448 , n2166 , n2169 );
or ( n2449 , n2446 , n2447 , n2448 );
and ( n2450 , n2177 , n2178 );
and ( n2451 , n2178 , n2180 );
and ( n2452 , n2177 , n2180 );
or ( n2453 , n2450 , n2451 , n2452 );
xor ( n2454 , n2449 , n2453 );
and ( n2455 , n782 , n852 );
and ( n2456 , n931 , n714 );
xor ( n2457 , n2455 , n2456 );
and ( n2458 , n1088 , n651 );
xor ( n2459 , n2457 , n2458 );
xor ( n2460 , n2454 , n2459 );
xor ( n2461 , n2445 , n2460 );
and ( n2462 , n2183 , n2184 );
and ( n2463 , n2184 , n2287 );
and ( n2464 , n2183 , n2287 );
or ( n2465 , n2462 , n2463 , n2464 );
and ( n2466 , n1292 , n488 );
and ( n2467 , n1516 , n411 );
xor ( n2468 , n2466 , n2467 );
and ( n2469 , n1730 , n375 );
xor ( n2470 , n2468 , n2469 );
xor ( n2471 , n2465 , n2470 );
and ( n2472 , n2001 , n312 );
and ( n2473 , n2286 , n288 );
xor ( n2474 , n2472 , n2473 );
and ( n2475 , n2199 , n2203 );
and ( n2476 , n2203 , n2209 );
and ( n2477 , n2199 , n2209 );
or ( n2478 , n2475 , n2476 , n2477 );
and ( n2479 , n2195 , n2210 );
and ( n2480 , n2210 , n2278 );
and ( n2481 , n2195 , n2278 );
or ( n2482 , n2479 , n2480 , n2481 );
xor ( n2483 , n2478 , n2482 );
and ( n2484 , n2215 , n2241 );
and ( n2485 , n2241 , n2277 );
and ( n2486 , n2215 , n2277 );
or ( n2487 , n2484 , n2485 , n2486 );
and ( n2488 , n2229 , n2230 );
and ( n2489 , n2230 , n2232 );
and ( n2490 , n2229 , n2232 );
or ( n2491 , n2488 , n2489 , n2490 );
and ( n2492 , n2219 , n2223 );
and ( n2493 , n2223 , n2240 );
and ( n2494 , n2219 , n2240 );
or ( n2495 , n2492 , n2493 , n2494 );
xor ( n2496 , n2491 , n2495 );
and ( n2497 , n2206 , n291 );
not ( n2498 , n291 );
nor ( n2499 , n2497 , n2498 );
xor ( n2500 , n2496 , n2499 );
xor ( n2501 , n2487 , n2500 );
and ( n2502 , n2246 , n2261 );
and ( n2503 , n2261 , n2276 );
and ( n2504 , n2246 , n2276 );
or ( n2505 , n2502 , n2503 , n2504 );
and ( n2506 , n2228 , n2233 );
and ( n2507 , n2233 , n2239 );
and ( n2508 , n2228 , n2239 );
or ( n2509 , n2506 , n2507 , n2508 );
and ( n2510 , n2250 , n2254 );
and ( n2511 , n2254 , n2260 );
and ( n2512 , n2250 , n2260 );
or ( n2513 , n2510 , n2511 , n2512 );
xor ( n2514 , n2509 , n2513 );
and ( n2515 , n2235 , n2236 );
and ( n2516 , n2236 , n2238 );
and ( n2517 , n2235 , n2238 );
or ( n2518 , n2515 , n2516 , n2517 );
and ( n2519 , n1458 , n435 );
and ( n2520 , n1713 , n354 );
xor ( n2521 , n2519 , n2520 );
and ( n2522 , n1935 , n321 );
xor ( n2523 , n2521 , n2522 );
xor ( n2524 , n2518 , n2523 );
and ( n2525 , n917 , n766 );
and ( n2526 , n1077 , n607 );
xor ( n2527 , n2525 , n2526 );
and ( n2528 , n1277 , n510 );
xor ( n2529 , n2527 , n2528 );
xor ( n2530 , n2524 , n2529 );
xor ( n2531 , n2514 , n2530 );
xor ( n2532 , n2505 , n2531 );
and ( n2533 , n2264 , n2269 );
and ( n2534 , n2269 , n2275 );
and ( n2535 , n2264 , n2275 );
or ( n2536 , n2533 , n2534 , n2535 );
and ( n2537 , n2256 , n2257 );
and ( n2538 , n2257 , n2259 );
and ( n2539 , n2256 , n2259 );
or ( n2540 , n2537 , n2538 , n2539 );
and ( n2541 , n2265 , n2266 );
and ( n2542 , n2266 , n2268 );
and ( n2543 , n2265 , n2268 );
or ( n2544 , n2541 , n2542 , n2543 );
xor ( n2545 , n2540 , n2544 );
and ( n2546 , n521 , n1261 );
and ( n2547 , n625 , n1048 );
xor ( n2548 , n2546 , n2547 );
and ( n2549 , n753 , n905 );
xor ( n2550 , n2548 , n2549 );
xor ( n2551 , n2545 , n2550 );
xor ( n2552 , n2536 , n2551 );
and ( n2553 , n2272 , n2274 );
buf ( n2554 , n2553 );
and ( n2555 , n318 , n1975 );
and ( n2556 , n361 , n1685 );
xor ( n2557 , n2555 , n2556 );
and ( n2558 , n431 , n1497 );
xor ( n2559 , n2557 , n2558 );
xor ( n2560 , n2554 , n2559 );
not ( n2561 , n273 );
buf ( n2562 , n241 );
not ( n2563 , n2562 );
and ( n2564 , n2563 , n273 );
nor ( n2565 , n2561 , n2564 );
and ( n2566 , n294 , n2271 );
xor ( n2567 , n2565 , n2566 );
xor ( n2568 , n2560 , n2567 );
xor ( n2569 , n2552 , n2568 );
xor ( n2570 , n2532 , n2569 );
xor ( n2571 , n2501 , n2570 );
xor ( n2572 , n2483 , n2571 );
and ( n2573 , n2186 , n2190 );
and ( n2574 , n2190 , n2279 );
and ( n2575 , n2186 , n2279 );
or ( n2576 , n2573 , n2574 , n2575 );
xor ( n2577 , n2572 , n2576 );
and ( n2578 , n2280 , n2283 );
xor ( n2579 , n2577 , n2578 );
buf ( n2580 , n2579 );
buf ( n2581 , n2580 );
and ( n2582 , n2581 , n279 );
xor ( n2583 , n2474 , n2582 );
xor ( n2584 , n2471 , n2583 );
xor ( n2585 , n2461 , n2584 );
xor ( n2586 , n2441 , n2585 );
xor ( n2587 , n2410 , n2586 );
xor ( n2588 , n2390 , n2587 );
and ( n2589 , n2106 , n2292 );
buf ( n2590 , n2589 );
xor ( n2591 , n2588 , n2590 );
and ( n2592 , n2293 , n2296 );
xor ( n2593 , n2591 , n2592 );
buf ( n2594 , n2593 );
buf ( n2595 , n2594 );
not ( n2596 , n2595 );
buf ( n2597 , n210 );
not ( n2598 , n2597 );
nor ( n2599 , n2596 , n2598 );
xor ( n2600 , n2383 , n2599 );
xor ( n2601 , n2308 , n2380 );
nor ( n2602 , n2300 , n2598 );
and ( n2603 , n2601 , n2602 );
xor ( n2604 , n2601 , n2602 );
xor ( n2605 , n2312 , n2378 );
nor ( n2606 , n2025 , n2598 );
and ( n2607 , n2605 , n2606 );
xor ( n2608 , n2605 , n2606 );
xor ( n2609 , n2316 , n2376 );
nor ( n2610 , n1771 , n2598 );
and ( n2611 , n2609 , n2610 );
xor ( n2612 , n2609 , n2610 );
xor ( n2613 , n2320 , n2374 );
nor ( n2614 , n1534 , n2598 );
and ( n2615 , n2613 , n2614 );
xor ( n2616 , n2613 , n2614 );
xor ( n2617 , n2324 , n2372 );
nor ( n2618 , n1318 , n2598 );
and ( n2619 , n2617 , n2618 );
xor ( n2620 , n2617 , n2618 );
xor ( n2621 , n2328 , n2370 );
nor ( n2622 , n1126 , n2598 );
and ( n2623 , n2621 , n2622 );
xor ( n2624 , n2621 , n2622 );
xor ( n2625 , n2332 , n2368 );
nor ( n2626 , n952 , n2598 );
and ( n2627 , n2625 , n2626 );
xor ( n2628 , n2625 , n2626 );
xor ( n2629 , n2336 , n2366 );
nor ( n2630 , n795 , n2598 );
and ( n2631 , n2629 , n2630 );
xor ( n2632 , n2629 , n2630 );
xor ( n2633 , n2340 , n2364 );
nor ( n2634 , n663 , n2598 );
and ( n2635 , n2633 , n2634 );
xor ( n2636 , n2633 , n2634 );
xor ( n2637 , n2344 , n2362 );
nor ( n2638 , n549 , n2598 );
and ( n2639 , n2637 , n2638 );
xor ( n2640 , n2637 , n2638 );
xor ( n2641 , n2348 , n2360 );
nor ( n2642 , n456 , n2598 );
and ( n2643 , n2641 , n2642 );
xor ( n2644 , n2641 , n2642 );
xor ( n2645 , n2353 , n2358 );
nor ( n2646 , n384 , n2598 );
and ( n2647 , n2645 , n2646 );
xor ( n2648 , n2645 , n2646 );
xor ( n2649 , n2355 , n2356 );
buf ( n2650 , n2649 );
nor ( n2651 , n334 , n2598 );
and ( n2652 , n2650 , n2651 );
xor ( n2653 , n2650 , n2651 );
nor ( n2654 , n283 , n2302 );
buf ( n2655 , n2654 );
nor ( n2656 , n303 , n2598 );
and ( n2657 , n2655 , n2656 );
buf ( n2658 , n2657 );
and ( n2659 , n2653 , n2658 );
or ( n2660 , n2652 , n2659 );
and ( n2661 , n2648 , n2660 );
or ( n2662 , n2647 , n2661 );
and ( n2663 , n2644 , n2662 );
or ( n2664 , n2643 , n2663 );
and ( n2665 , n2640 , n2664 );
or ( n2666 , n2639 , n2665 );
and ( n2667 , n2636 , n2666 );
or ( n2668 , n2635 , n2667 );
and ( n2669 , n2632 , n2668 );
or ( n2670 , n2631 , n2669 );
and ( n2671 , n2628 , n2670 );
or ( n2672 , n2627 , n2671 );
and ( n2673 , n2624 , n2672 );
or ( n2674 , n2623 , n2673 );
and ( n2675 , n2620 , n2674 );
or ( n2676 , n2619 , n2675 );
and ( n2677 , n2616 , n2676 );
or ( n2678 , n2615 , n2677 );
and ( n2679 , n2612 , n2678 );
or ( n2680 , n2611 , n2679 );
and ( n2681 , n2608 , n2680 );
or ( n2682 , n2607 , n2681 );
and ( n2683 , n2604 , n2682 );
or ( n2684 , n2603 , n2683 );
xor ( n2685 , n2600 , n2684 );
buf ( n2686 , n2685 );
buf ( n2687 , n2686 );
not ( n2688 , n2687 );
buf ( n2689 , n257 );
not ( n2690 , n2689 );
and ( n2691 , n2690 , n2687 );
nor ( n2692 , n2688 , n2691 );
and ( n2693 , n285 , n302 );
nor ( n2694 , n303 , n2693 );
nor ( n2695 , n334 , n305 );
xor ( n2696 , n2694 , n2695 );
and ( n2697 , n287 , n306 );
buf ( n2698 , n2697 );
xor ( n2699 , n2696 , n2698 );
nor ( n2700 , n384 , n336 );
xor ( n2701 , n2699 , n2700 );
and ( n2702 , n308 , n337 );
and ( n2703 , n338 , n343 );
or ( n2704 , n2702 , n2703 );
xor ( n2705 , n2701 , n2704 );
nor ( n2706 , n456 , n386 );
xor ( n2707 , n2705 , n2706 );
and ( n2708 , n344 , n387 );
and ( n2709 , n388 , n400 );
or ( n2710 , n2708 , n2709 );
xor ( n2711 , n2707 , n2710 );
nor ( n2712 , n549 , n458 );
xor ( n2713 , n2711 , n2712 );
and ( n2714 , n401 , n459 );
and ( n2715 , n460 , n478 );
or ( n2716 , n2714 , n2715 );
xor ( n2717 , n2713 , n2716 );
nor ( n2718 , n663 , n551 );
xor ( n2719 , n2717 , n2718 );
and ( n2720 , n479 , n552 );
and ( n2721 , n553 , n577 );
or ( n2722 , n2720 , n2721 );
xor ( n2723 , n2719 , n2722 );
nor ( n2724 , n795 , n665 );
xor ( n2725 , n2723 , n2724 );
and ( n2726 , n578 , n666 );
and ( n2727 , n667 , n697 );
or ( n2728 , n2726 , n2727 );
xor ( n2729 , n2725 , n2728 );
nor ( n2730 , n952 , n797 );
xor ( n2731 , n2729 , n2730 );
and ( n2732 , n698 , n798 );
and ( n2733 , n799 , n835 );
or ( n2734 , n2732 , n2733 );
xor ( n2735 , n2731 , n2734 );
nor ( n2736 , n1126 , n954 );
xor ( n2737 , n2735 , n2736 );
and ( n2738 , n836 , n955 );
and ( n2739 , n956 , n998 );
or ( n2740 , n2738 , n2739 );
xor ( n2741 , n2737 , n2740 );
nor ( n2742 , n1318 , n1128 );
xor ( n2743 , n2741 , n2742 );
and ( n2744 , n999 , n1129 );
and ( n2745 , n1130 , n1178 );
or ( n2746 , n2744 , n2745 );
xor ( n2747 , n2743 , n2746 );
nor ( n2748 , n1534 , n1320 );
xor ( n2749 , n2747 , n2748 );
and ( n2750 , n1179 , n1321 );
and ( n2751 , n1322 , n1376 );
or ( n2752 , n2750 , n2751 );
xor ( n2753 , n2749 , n2752 );
nor ( n2754 , n1771 , n1536 );
xor ( n2755 , n2753 , n2754 );
and ( n2756 , n1377 , n1537 );
and ( n2757 , n1538 , n1598 );
or ( n2758 , n2756 , n2757 );
xor ( n2759 , n2755 , n2758 );
nor ( n2760 , n2025 , n1773 );
xor ( n2761 , n2759 , n2760 );
and ( n2762 , n1599 , n1774 );
and ( n2763 , n1775 , n1841 );
or ( n2764 , n2762 , n2763 );
xor ( n2765 , n2761 , n2764 );
nor ( n2766 , n2300 , n2027 );
xor ( n2767 , n2765 , n2766 );
and ( n2768 , n1842 , n2028 );
and ( n2769 , n2029 , n2101 );
or ( n2770 , n2768 , n2769 );
xor ( n2771 , n2767 , n2770 );
nor ( n2772 , n2596 , n2302 );
xor ( n2773 , n2771 , n2772 );
and ( n2774 , n2102 , n2303 );
and ( n2775 , n2304 , n2382 );
or ( n2776 , n2774 , n2775 );
xor ( n2777 , n2773 , n2776 );
and ( n2778 , n2398 , n2402 );
and ( n2779 , n2402 , n2408 );
and ( n2780 , n2398 , n2408 );
or ( n2781 , n2778 , n2779 , n2780 );
and ( n2782 , n2394 , n2409 );
and ( n2783 , n2409 , n2586 );
and ( n2784 , n2394 , n2586 );
or ( n2785 , n2782 , n2783 , n2784 );
xor ( n2786 , n2781 , n2785 );
and ( n2787 , n2414 , n2440 );
and ( n2788 , n2440 , n2585 );
and ( n2789 , n2414 , n2585 );
or ( n2790 , n2787 , n2788 , n2789 );
and ( n2791 , n2428 , n2429 );
and ( n2792 , n2429 , n2431 );
and ( n2793 , n2428 , n2431 );
or ( n2794 , n2791 , n2792 , n2793 );
and ( n2795 , n2418 , n2422 );
and ( n2796 , n2422 , n2439 );
and ( n2797 , n2418 , n2439 );
or ( n2798 , n2795 , n2796 , n2797 );
xor ( n2799 , n2794 , n2798 );
not ( n2800 , n298 );
and ( n2801 , n2406 , n298 );
nor ( n2802 , n2800 , n2801 );
xor ( n2803 , n2799 , n2802 );
xor ( n2804 , n2790 , n2803 );
and ( n2805 , n2445 , n2460 );
and ( n2806 , n2460 , n2584 );
and ( n2807 , n2445 , n2584 );
or ( n2808 , n2805 , n2806 , n2807 );
and ( n2809 , n2427 , n2432 );
and ( n2810 , n2432 , n2438 );
and ( n2811 , n2427 , n2438 );
or ( n2812 , n2809 , n2810 , n2811 );
and ( n2813 , n2449 , n2453 );
and ( n2814 , n2453 , n2459 );
and ( n2815 , n2449 , n2459 );
or ( n2816 , n2813 , n2814 , n2815 );
xor ( n2817 , n2812 , n2816 );
and ( n2818 , n2434 , n2435 );
and ( n2819 , n2435 , n2437 );
and ( n2820 , n2434 , n2437 );
or ( n2821 , n2818 , n2819 , n2820 );
and ( n2822 , n328 , n2138 );
and ( n2823 , n371 , n1864 );
xor ( n2824 , n2822 , n2823 );
and ( n2825 , n446 , n1753 );
xor ( n2826 , n2824 , n2825 );
xor ( n2827 , n2821 , n2826 );
and ( n2828 , n533 , n1396 );
and ( n2829 , n636 , n1302 );
xor ( n2830 , n2828 , n2829 );
and ( n2831 , n782 , n1114 );
xor ( n2832 , n2830 , n2831 );
xor ( n2833 , n2827 , n2832 );
xor ( n2834 , n2817 , n2833 );
xor ( n2835 , n2808 , n2834 );
and ( n2836 , n2465 , n2470 );
and ( n2837 , n2470 , n2583 );
and ( n2838 , n2465 , n2583 );
or ( n2839 , n2836 , n2837 , n2838 );
and ( n2840 , n2455 , n2456 );
and ( n2841 , n2456 , n2458 );
and ( n2842 , n2455 , n2458 );
or ( n2843 , n2840 , n2841 , n2842 );
and ( n2844 , n2466 , n2467 );
and ( n2845 , n2467 , n2469 );
and ( n2846 , n2466 , n2469 );
or ( n2847 , n2844 , n2845 , n2846 );
xor ( n2848 , n2843 , n2847 );
and ( n2849 , n931 , n852 );
and ( n2850 , n1088 , n714 );
xor ( n2851 , n2849 , n2850 );
and ( n2852 , n1292 , n651 );
xor ( n2853 , n2851 , n2852 );
xor ( n2854 , n2848 , n2853 );
xor ( n2855 , n2839 , n2854 );
and ( n2856 , n2472 , n2473 );
and ( n2857 , n2473 , n2582 );
and ( n2858 , n2472 , n2582 );
or ( n2859 , n2856 , n2857 , n2858 );
and ( n2860 , n1516 , n488 );
and ( n2861 , n1730 , n411 );
xor ( n2862 , n2860 , n2861 );
and ( n2863 , n2001 , n375 );
xor ( n2864 , n2862 , n2863 );
xor ( n2865 , n2859 , n2864 );
and ( n2866 , n2286 , n312 );
and ( n2867 , n2581 , n288 );
xor ( n2868 , n2866 , n2867 );
and ( n2869 , n2491 , n2495 );
and ( n2870 , n2495 , n2499 );
and ( n2871 , n2491 , n2499 );
or ( n2872 , n2869 , n2870 , n2871 );
and ( n2873 , n2487 , n2500 );
and ( n2874 , n2500 , n2570 );
and ( n2875 , n2487 , n2570 );
or ( n2876 , n2873 , n2874 , n2875 );
xor ( n2877 , n2872 , n2876 );
and ( n2878 , n2505 , n2531 );
and ( n2879 , n2531 , n2569 );
and ( n2880 , n2505 , n2569 );
or ( n2881 , n2878 , n2879 , n2880 );
and ( n2882 , n2519 , n2520 );
and ( n2883 , n2520 , n2522 );
and ( n2884 , n2519 , n2522 );
or ( n2885 , n2882 , n2883 , n2884 );
and ( n2886 , n2509 , n2513 );
and ( n2887 , n2513 , n2530 );
and ( n2888 , n2509 , n2530 );
or ( n2889 , n2886 , n2887 , n2888 );
xor ( n2890 , n2885 , n2889 );
and ( n2891 , n2206 , n321 );
not ( n2892 , n321 );
nor ( n2893 , n2891 , n2892 );
xor ( n2894 , n2890 , n2893 );
xor ( n2895 , n2881 , n2894 );
and ( n2896 , n2536 , n2551 );
and ( n2897 , n2551 , n2568 );
and ( n2898 , n2536 , n2568 );
or ( n2899 , n2896 , n2897 , n2898 );
and ( n2900 , n2518 , n2523 );
and ( n2901 , n2523 , n2529 );
and ( n2902 , n2518 , n2529 );
or ( n2903 , n2900 , n2901 , n2902 );
and ( n2904 , n2540 , n2544 );
and ( n2905 , n2544 , n2550 );
and ( n2906 , n2540 , n2550 );
or ( n2907 , n2904 , n2905 , n2906 );
xor ( n2908 , n2903 , n2907 );
and ( n2909 , n2525 , n2526 );
and ( n2910 , n2526 , n2528 );
and ( n2911 , n2525 , n2528 );
or ( n2912 , n2909 , n2910 , n2911 );
and ( n2913 , n1458 , n510 );
and ( n2914 , n1713 , n435 );
xor ( n2915 , n2913 , n2914 );
and ( n2916 , n1935 , n354 );
xor ( n2917 , n2915 , n2916 );
xor ( n2918 , n2912 , n2917 );
and ( n2919 , n917 , n905 );
and ( n2920 , n1077 , n766 );
xor ( n2921 , n2919 , n2920 );
and ( n2922 , n1277 , n607 );
xor ( n2923 , n2921 , n2922 );
xor ( n2924 , n2918 , n2923 );
xor ( n2925 , n2908 , n2924 );
xor ( n2926 , n2899 , n2925 );
and ( n2927 , n2554 , n2559 );
and ( n2928 , n2559 , n2567 );
and ( n2929 , n2554 , n2567 );
or ( n2930 , n2927 , n2928 , n2929 );
and ( n2931 , n2546 , n2547 );
and ( n2932 , n2547 , n2549 );
and ( n2933 , n2546 , n2549 );
or ( n2934 , n2931 , n2932 , n2933 );
and ( n2935 , n2555 , n2556 );
and ( n2936 , n2556 , n2558 );
and ( n2937 , n2555 , n2558 );
or ( n2938 , n2935 , n2936 , n2937 );
xor ( n2939 , n2934 , n2938 );
and ( n2940 , n521 , n1497 );
and ( n2941 , n625 , n1261 );
xor ( n2942 , n2940 , n2941 );
and ( n2943 , n753 , n1048 );
xor ( n2944 , n2942 , n2943 );
xor ( n2945 , n2939 , n2944 );
xor ( n2946 , n2930 , n2945 );
and ( n2947 , n2565 , n2566 );
not ( n2948 , n294 );
and ( n2949 , n2563 , n294 );
nor ( n2950 , n2948 , n2949 );
xor ( n2951 , n2947 , n2950 );
and ( n2952 , n318 , n2271 );
and ( n2953 , n361 , n1975 );
xor ( n2954 , n2952 , n2953 );
and ( n2955 , n431 , n1685 );
xor ( n2956 , n2954 , n2955 );
xor ( n2957 , n2951 , n2956 );
xor ( n2958 , n2946 , n2957 );
xor ( n2959 , n2926 , n2958 );
xor ( n2960 , n2895 , n2959 );
xor ( n2961 , n2877 , n2960 );
and ( n2962 , n2478 , n2482 );
and ( n2963 , n2482 , n2571 );
and ( n2964 , n2478 , n2571 );
or ( n2965 , n2962 , n2963 , n2964 );
xor ( n2966 , n2961 , n2965 );
and ( n2967 , n2572 , n2576 );
and ( n2968 , n2577 , n2578 );
or ( n2969 , n2967 , n2968 );
xor ( n2970 , n2966 , n2969 );
buf ( n2971 , n2970 );
buf ( n2972 , n2971 );
and ( n2973 , n2972 , n279 );
xor ( n2974 , n2868 , n2973 );
xor ( n2975 , n2865 , n2974 );
xor ( n2976 , n2855 , n2975 );
xor ( n2977 , n2835 , n2976 );
xor ( n2978 , n2804 , n2977 );
xor ( n2979 , n2786 , n2978 );
and ( n2980 , n2385 , n2389 );
and ( n2981 , n2389 , n2587 );
and ( n2982 , n2385 , n2587 );
or ( n2983 , n2980 , n2981 , n2982 );
xor ( n2984 , n2979 , n2983 );
and ( n2985 , n2588 , n2590 );
and ( n2986 , n2591 , n2592 );
or ( n2987 , n2985 , n2986 );
xor ( n2988 , n2984 , n2987 );
buf ( n2989 , n2988 );
buf ( n2990 , n2989 );
not ( n2991 , n2990 );
nor ( n2992 , n2991 , n2598 );
xor ( n2993 , n2777 , n2992 );
and ( n2994 , n2383 , n2599 );
and ( n2995 , n2600 , n2684 );
or ( n2996 , n2994 , n2995 );
xor ( n2997 , n2993 , n2996 );
buf ( n2998 , n2997 );
buf ( n2999 , n2998 );
not ( n3000 , n2999 );
buf ( n3001 , n258 );
not ( n3002 , n3001 );
nor ( n3003 , n3000 , n3002 );
xor ( n3004 , n2692 , n3003 );
xor ( n3005 , n2604 , n2682 );
buf ( n3006 , n3005 );
buf ( n3007 , n3006 );
not ( n3008 , n3007 );
and ( n3009 , n2690 , n3007 );
nor ( n3010 , n3008 , n3009 );
nor ( n3011 , n2688 , n3002 );
and ( n3012 , n3010 , n3011 );
xor ( n3013 , n3010 , n3011 );
xor ( n3014 , n2608 , n2680 );
buf ( n3015 , n3014 );
buf ( n3016 , n3015 );
not ( n3017 , n3016 );
and ( n3018 , n2690 , n3016 );
nor ( n3019 , n3017 , n3018 );
nor ( n3020 , n3008 , n3002 );
and ( n3021 , n3019 , n3020 );
xor ( n3022 , n3019 , n3020 );
xor ( n3023 , n2612 , n2678 );
buf ( n3024 , n3023 );
buf ( n3025 , n3024 );
not ( n3026 , n3025 );
and ( n3027 , n2690 , n3025 );
nor ( n3028 , n3026 , n3027 );
nor ( n3029 , n3017 , n3002 );
and ( n3030 , n3028 , n3029 );
xor ( n3031 , n3028 , n3029 );
xor ( n3032 , n2616 , n2676 );
buf ( n3033 , n3032 );
buf ( n3034 , n3033 );
not ( n3035 , n3034 );
and ( n3036 , n2690 , n3034 );
nor ( n3037 , n3035 , n3036 );
nor ( n3038 , n3026 , n3002 );
and ( n3039 , n3037 , n3038 );
xor ( n3040 , n3037 , n3038 );
xor ( n3041 , n2620 , n2674 );
buf ( n3042 , n3041 );
buf ( n3043 , n3042 );
not ( n3044 , n3043 );
and ( n3045 , n2690 , n3043 );
nor ( n3046 , n3044 , n3045 );
nor ( n3047 , n3035 , n3002 );
and ( n3048 , n3046 , n3047 );
xor ( n3049 , n3046 , n3047 );
xor ( n3050 , n2624 , n2672 );
buf ( n3051 , n3050 );
buf ( n3052 , n3051 );
not ( n3053 , n3052 );
and ( n3054 , n2690 , n3052 );
nor ( n3055 , n3053 , n3054 );
nor ( n3056 , n3044 , n3002 );
and ( n3057 , n3055 , n3056 );
xor ( n3058 , n3055 , n3056 );
xor ( n3059 , n2628 , n2670 );
buf ( n3060 , n3059 );
buf ( n3061 , n3060 );
not ( n3062 , n3061 );
and ( n3063 , n2690 , n3061 );
nor ( n3064 , n3062 , n3063 );
nor ( n3065 , n3053 , n3002 );
and ( n3066 , n3064 , n3065 );
xor ( n3067 , n3064 , n3065 );
xor ( n3068 , n2632 , n2668 );
buf ( n3069 , n3068 );
buf ( n3070 , n3069 );
not ( n3071 , n3070 );
and ( n3072 , n2690 , n3070 );
nor ( n3073 , n3071 , n3072 );
nor ( n3074 , n3062 , n3002 );
and ( n3075 , n3073 , n3074 );
xor ( n3076 , n3073 , n3074 );
xor ( n3077 , n2636 , n2666 );
buf ( n3078 , n3077 );
buf ( n3079 , n3078 );
not ( n3080 , n3079 );
and ( n3081 , n2690 , n3079 );
nor ( n3082 , n3080 , n3081 );
nor ( n3083 , n3071 , n3002 );
and ( n3084 , n3082 , n3083 );
xor ( n3085 , n3082 , n3083 );
xor ( n3086 , n2640 , n2664 );
buf ( n3087 , n3086 );
buf ( n3088 , n3087 );
not ( n3089 , n3088 );
and ( n3090 , n2690 , n3088 );
nor ( n3091 , n3089 , n3090 );
nor ( n3092 , n3080 , n3002 );
and ( n3093 , n3091 , n3092 );
xor ( n3094 , n3091 , n3092 );
xor ( n3095 , n2644 , n2662 );
buf ( n3096 , n3095 );
buf ( n3097 , n3096 );
not ( n3098 , n3097 );
and ( n3099 , n2690 , n3097 );
nor ( n3100 , n3098 , n3099 );
nor ( n3101 , n3089 , n3002 );
and ( n3102 , n3100 , n3101 );
xor ( n3103 , n3100 , n3101 );
xor ( n3104 , n2648 , n2660 );
buf ( n3105 , n3104 );
buf ( n3106 , n3105 );
not ( n3107 , n3106 );
and ( n3108 , n2690 , n3106 );
nor ( n3109 , n3107 , n3108 );
nor ( n3110 , n3098 , n3002 );
and ( n3111 , n3109 , n3110 );
xor ( n3112 , n3109 , n3110 );
xor ( n3113 , n2653 , n2658 );
buf ( n3114 , n3113 );
buf ( n3115 , n3114 );
not ( n3116 , n3115 );
and ( n3117 , n2690 , n3115 );
nor ( n3118 , n3116 , n3117 );
nor ( n3119 , n3107 , n3002 );
and ( n3120 , n3118 , n3119 );
xor ( n3121 , n3118 , n3119 );
xor ( n3122 , n2655 , n2656 );
buf ( n3123 , n3122 );
buf ( n3124 , n3123 );
not ( n3125 , n3124 );
and ( n3126 , n2690 , n3124 );
nor ( n3127 , n3125 , n3126 );
nor ( n3128 , n3116 , n3002 );
and ( n3129 , n3127 , n3128 );
xor ( n3130 , n3127 , n3128 );
nor ( n3131 , n283 , n2598 );
buf ( n3132 , n3131 );
buf ( n3133 , n3132 );
not ( n3134 , n3133 );
and ( n3135 , n2690 , n3133 );
nor ( n3136 , n3134 , n3135 );
nor ( n3137 , n3125 , n3002 );
and ( n3138 , n3136 , n3137 );
buf ( n3139 , n3138 );
and ( n3140 , n3130 , n3139 );
or ( n3141 , n3129 , n3140 );
and ( n3142 , n3121 , n3141 );
or ( n3143 , n3120 , n3142 );
and ( n3144 , n3112 , n3143 );
or ( n3145 , n3111 , n3144 );
and ( n3146 , n3103 , n3145 );
or ( n3147 , n3102 , n3146 );
and ( n3148 , n3094 , n3147 );
or ( n3149 , n3093 , n3148 );
and ( n3150 , n3085 , n3149 );
or ( n3151 , n3084 , n3150 );
and ( n3152 , n3076 , n3151 );
or ( n3153 , n3075 , n3152 );
and ( n3154 , n3067 , n3153 );
or ( n3155 , n3066 , n3154 );
and ( n3156 , n3058 , n3155 );
or ( n3157 , n3057 , n3156 );
and ( n3158 , n3049 , n3157 );
or ( n3159 , n3048 , n3158 );
and ( n3160 , n3040 , n3159 );
or ( n3161 , n3039 , n3160 );
and ( n3162 , n3031 , n3161 );
or ( n3163 , n3030 , n3162 );
and ( n3164 , n3022 , n3163 );
or ( n3165 , n3021 , n3164 );
and ( n3166 , n3013 , n3165 );
or ( n3167 , n3012 , n3166 );
xor ( n3168 , n3004 , n3167 );
and ( n3169 , n285 , n333 );
nor ( n3170 , n334 , n3169 );
nor ( n3171 , n384 , n305 );
xor ( n3172 , n3170 , n3171 );
and ( n3173 , n2694 , n2695 );
and ( n3174 , n2696 , n2698 );
or ( n3175 , n3173 , n3174 );
xor ( n3176 , n3172 , n3175 );
nor ( n3177 , n456 , n336 );
xor ( n3178 , n3176 , n3177 );
and ( n3179 , n2699 , n2700 );
and ( n3180 , n2701 , n2704 );
or ( n3181 , n3179 , n3180 );
xor ( n3182 , n3178 , n3181 );
nor ( n3183 , n549 , n386 );
xor ( n3184 , n3182 , n3183 );
and ( n3185 , n2705 , n2706 );
and ( n3186 , n2707 , n2710 );
or ( n3187 , n3185 , n3186 );
xor ( n3188 , n3184 , n3187 );
nor ( n3189 , n663 , n458 );
xor ( n3190 , n3188 , n3189 );
and ( n3191 , n2711 , n2712 );
and ( n3192 , n2713 , n2716 );
or ( n3193 , n3191 , n3192 );
xor ( n3194 , n3190 , n3193 );
nor ( n3195 , n795 , n551 );
xor ( n3196 , n3194 , n3195 );
and ( n3197 , n2717 , n2718 );
and ( n3198 , n2719 , n2722 );
or ( n3199 , n3197 , n3198 );
xor ( n3200 , n3196 , n3199 );
nor ( n3201 , n952 , n665 );
xor ( n3202 , n3200 , n3201 );
and ( n3203 , n2723 , n2724 );
and ( n3204 , n2725 , n2728 );
or ( n3205 , n3203 , n3204 );
xor ( n3206 , n3202 , n3205 );
nor ( n3207 , n1126 , n797 );
xor ( n3208 , n3206 , n3207 );
and ( n3209 , n2729 , n2730 );
and ( n3210 , n2731 , n2734 );
or ( n3211 , n3209 , n3210 );
xor ( n3212 , n3208 , n3211 );
nor ( n3213 , n1318 , n954 );
xor ( n3214 , n3212 , n3213 );
and ( n3215 , n2735 , n2736 );
and ( n3216 , n2737 , n2740 );
or ( n3217 , n3215 , n3216 );
xor ( n3218 , n3214 , n3217 );
nor ( n3219 , n1534 , n1128 );
xor ( n3220 , n3218 , n3219 );
and ( n3221 , n2741 , n2742 );
and ( n3222 , n2743 , n2746 );
or ( n3223 , n3221 , n3222 );
xor ( n3224 , n3220 , n3223 );
nor ( n3225 , n1771 , n1320 );
xor ( n3226 , n3224 , n3225 );
and ( n3227 , n2747 , n2748 );
and ( n3228 , n2749 , n2752 );
or ( n3229 , n3227 , n3228 );
xor ( n3230 , n3226 , n3229 );
nor ( n3231 , n2025 , n1536 );
xor ( n3232 , n3230 , n3231 );
and ( n3233 , n2753 , n2754 );
and ( n3234 , n2755 , n2758 );
or ( n3235 , n3233 , n3234 );
xor ( n3236 , n3232 , n3235 );
nor ( n3237 , n2300 , n1773 );
xor ( n3238 , n3236 , n3237 );
and ( n3239 , n2759 , n2760 );
and ( n3240 , n2761 , n2764 );
or ( n3241 , n3239 , n3240 );
xor ( n3242 , n3238 , n3241 );
nor ( n3243 , n2596 , n2027 );
xor ( n3244 , n3242 , n3243 );
and ( n3245 , n2765 , n2766 );
and ( n3246 , n2767 , n2770 );
or ( n3247 , n3245 , n3246 );
xor ( n3248 , n3244 , n3247 );
nor ( n3249 , n2991 , n2302 );
xor ( n3250 , n3248 , n3249 );
and ( n3251 , n2771 , n2772 );
and ( n3252 , n2773 , n2776 );
or ( n3253 , n3251 , n3252 );
xor ( n3254 , n3250 , n3253 );
and ( n3255 , n2794 , n2798 );
and ( n3256 , n2798 , n2802 );
and ( n3257 , n2794 , n2802 );
or ( n3258 , n3255 , n3256 , n3257 );
and ( n3259 , n2790 , n2803 );
and ( n3260 , n2803 , n2977 );
and ( n3261 , n2790 , n2977 );
or ( n3262 , n3259 , n3260 , n3261 );
xor ( n3263 , n3258 , n3262 );
and ( n3264 , n2808 , n2834 );
and ( n3265 , n2834 , n2976 );
and ( n3266 , n2808 , n2976 );
or ( n3267 , n3264 , n3265 , n3266 );
and ( n3268 , n2822 , n2823 );
and ( n3269 , n2823 , n2825 );
and ( n3270 , n2822 , n2825 );
or ( n3271 , n3268 , n3269 , n3270 );
and ( n3272 , n2812 , n2816 );
and ( n3273 , n2816 , n2833 );
and ( n3274 , n2812 , n2833 );
or ( n3275 , n3272 , n3273 , n3274 );
xor ( n3276 , n3271 , n3275 );
not ( n3277 , n328 );
and ( n3278 , n2406 , n328 );
nor ( n3279 , n3277 , n3278 );
xor ( n3280 , n3276 , n3279 );
xor ( n3281 , n3267 , n3280 );
and ( n3282 , n2839 , n2854 );
and ( n3283 , n2854 , n2975 );
and ( n3284 , n2839 , n2975 );
or ( n3285 , n3282 , n3283 , n3284 );
and ( n3286 , n2821 , n2826 );
and ( n3287 , n2826 , n2832 );
and ( n3288 , n2821 , n2832 );
or ( n3289 , n3286 , n3287 , n3288 );
and ( n3290 , n2843 , n2847 );
and ( n3291 , n2847 , n2853 );
and ( n3292 , n2843 , n2853 );
or ( n3293 , n3290 , n3291 , n3292 );
xor ( n3294 , n3289 , n3293 );
and ( n3295 , n2828 , n2829 );
and ( n3296 , n2829 , n2831 );
and ( n3297 , n2828 , n2831 );
or ( n3298 , n3295 , n3296 , n3297 );
and ( n3299 , n371 , n2138 );
and ( n3300 , n446 , n1864 );
xor ( n3301 , n3299 , n3300 );
and ( n3302 , n533 , n1753 );
xor ( n3303 , n3301 , n3302 );
xor ( n3304 , n3298 , n3303 );
and ( n3305 , n636 , n1396 );
and ( n3306 , n782 , n1302 );
xor ( n3307 , n3305 , n3306 );
and ( n3308 , n931 , n1114 );
xor ( n3309 , n3307 , n3308 );
xor ( n3310 , n3304 , n3309 );
xor ( n3311 , n3294 , n3310 );
xor ( n3312 , n3285 , n3311 );
and ( n3313 , n2859 , n2864 );
and ( n3314 , n2864 , n2974 );
and ( n3315 , n2859 , n2974 );
or ( n3316 , n3313 , n3314 , n3315 );
and ( n3317 , n2849 , n2850 );
and ( n3318 , n2850 , n2852 );
and ( n3319 , n2849 , n2852 );
or ( n3320 , n3317 , n3318 , n3319 );
and ( n3321 , n2860 , n2861 );
and ( n3322 , n2861 , n2863 );
and ( n3323 , n2860 , n2863 );
or ( n3324 , n3321 , n3322 , n3323 );
xor ( n3325 , n3320 , n3324 );
and ( n3326 , n1088 , n852 );
and ( n3327 , n1292 , n714 );
xor ( n3328 , n3326 , n3327 );
and ( n3329 , n1516 , n651 );
xor ( n3330 , n3328 , n3329 );
xor ( n3331 , n3325 , n3330 );
xor ( n3332 , n3316 , n3331 );
and ( n3333 , n2866 , n2867 );
and ( n3334 , n2867 , n2973 );
and ( n3335 , n2866 , n2973 );
or ( n3336 , n3333 , n3334 , n3335 );
and ( n3337 , n1730 , n488 );
and ( n3338 , n2001 , n411 );
xor ( n3339 , n3337 , n3338 );
and ( n3340 , n2286 , n375 );
xor ( n3341 , n3339 , n3340 );
xor ( n3342 , n3336 , n3341 );
and ( n3343 , n2581 , n312 );
and ( n3344 , n2972 , n288 );
xor ( n3345 , n3343 , n3344 );
and ( n3346 , n2885 , n2889 );
and ( n3347 , n2889 , n2893 );
and ( n3348 , n2885 , n2893 );
or ( n3349 , n3346 , n3347 , n3348 );
and ( n3350 , n2881 , n2894 );
and ( n3351 , n2894 , n2959 );
and ( n3352 , n2881 , n2959 );
or ( n3353 , n3350 , n3351 , n3352 );
xor ( n3354 , n3349 , n3353 );
and ( n3355 , n2899 , n2925 );
and ( n3356 , n2925 , n2958 );
and ( n3357 , n2899 , n2958 );
or ( n3358 , n3355 , n3356 , n3357 );
and ( n3359 , n2913 , n2914 );
and ( n3360 , n2914 , n2916 );
and ( n3361 , n2913 , n2916 );
or ( n3362 , n3359 , n3360 , n3361 );
and ( n3363 , n2903 , n2907 );
and ( n3364 , n2907 , n2924 );
and ( n3365 , n2903 , n2924 );
or ( n3366 , n3363 , n3364 , n3365 );
xor ( n3367 , n3362 , n3366 );
and ( n3368 , n2206 , n354 );
not ( n3369 , n354 );
nor ( n3370 , n3368 , n3369 );
xor ( n3371 , n3367 , n3370 );
xor ( n3372 , n3358 , n3371 );
and ( n3373 , n2930 , n2945 );
and ( n3374 , n2945 , n2957 );
and ( n3375 , n2930 , n2957 );
or ( n3376 , n3373 , n3374 , n3375 );
and ( n3377 , n2912 , n2917 );
and ( n3378 , n2917 , n2923 );
and ( n3379 , n2912 , n2923 );
or ( n3380 , n3377 , n3378 , n3379 );
and ( n3381 , n2934 , n2938 );
and ( n3382 , n2938 , n2944 );
and ( n3383 , n2934 , n2944 );
or ( n3384 , n3381 , n3382 , n3383 );
xor ( n3385 , n3380 , n3384 );
and ( n3386 , n2919 , n2920 );
and ( n3387 , n2920 , n2922 );
and ( n3388 , n2919 , n2922 );
or ( n3389 , n3386 , n3387 , n3388 );
and ( n3390 , n917 , n1048 );
and ( n3391 , n1077 , n905 );
xor ( n3392 , n3390 , n3391 );
and ( n3393 , n1277 , n766 );
xor ( n3394 , n3392 , n3393 );
xor ( n3395 , n3389 , n3394 );
and ( n3396 , n1458 , n607 );
and ( n3397 , n1713 , n510 );
xor ( n3398 , n3396 , n3397 );
and ( n3399 , n1935 , n435 );
xor ( n3400 , n3398 , n3399 );
xor ( n3401 , n3395 , n3400 );
xor ( n3402 , n3385 , n3401 );
xor ( n3403 , n3376 , n3402 );
and ( n3404 , n2947 , n2950 );
and ( n3405 , n2950 , n2956 );
and ( n3406 , n2947 , n2956 );
or ( n3407 , n3404 , n3405 , n3406 );
not ( n3408 , n318 );
and ( n3409 , n2563 , n318 );
nor ( n3410 , n3408 , n3409 );
and ( n3411 , n361 , n2271 );
xor ( n3412 , n3410 , n3411 );
and ( n3413 , n431 , n1975 );
xor ( n3414 , n3412 , n3413 );
xor ( n3415 , n3407 , n3414 );
and ( n3416 , n2940 , n2941 );
and ( n3417 , n2941 , n2943 );
and ( n3418 , n2940 , n2943 );
or ( n3419 , n3416 , n3417 , n3418 );
and ( n3420 , n2952 , n2953 );
and ( n3421 , n2953 , n2955 );
and ( n3422 , n2952 , n2955 );
or ( n3423 , n3420 , n3421 , n3422 );
xor ( n3424 , n3419 , n3423 );
and ( n3425 , n521 , n1685 );
and ( n3426 , n625 , n1497 );
xor ( n3427 , n3425 , n3426 );
and ( n3428 , n753 , n1261 );
xor ( n3429 , n3427 , n3428 );
xor ( n3430 , n3424 , n3429 );
xor ( n3431 , n3415 , n3430 );
xor ( n3432 , n3403 , n3431 );
xor ( n3433 , n3372 , n3432 );
xor ( n3434 , n3354 , n3433 );
and ( n3435 , n2872 , n2876 );
and ( n3436 , n2876 , n2960 );
and ( n3437 , n2872 , n2960 );
or ( n3438 , n3435 , n3436 , n3437 );
xor ( n3439 , n3434 , n3438 );
and ( n3440 , n2961 , n2965 );
and ( n3441 , n2966 , n2969 );
or ( n3442 , n3440 , n3441 );
xor ( n3443 , n3439 , n3442 );
buf ( n3444 , n3443 );
buf ( n3445 , n3444 );
and ( n3446 , n3445 , n279 );
xor ( n3447 , n3345 , n3446 );
xor ( n3448 , n3342 , n3447 );
xor ( n3449 , n3332 , n3448 );
xor ( n3450 , n3312 , n3449 );
xor ( n3451 , n3281 , n3450 );
xor ( n3452 , n3263 , n3451 );
and ( n3453 , n2781 , n2785 );
and ( n3454 , n2785 , n2978 );
and ( n3455 , n2781 , n2978 );
or ( n3456 , n3453 , n3454 , n3455 );
xor ( n3457 , n3452 , n3456 );
and ( n3458 , n2979 , n2983 );
and ( n3459 , n2984 , n2987 );
or ( n3460 , n3458 , n3459 );
xor ( n3461 , n3457 , n3460 );
buf ( n3462 , n3461 );
buf ( n3463 , n3462 );
not ( n3464 , n3463 );
nor ( n3465 , n3464 , n2598 );
xor ( n3466 , n3254 , n3465 );
and ( n3467 , n2777 , n2992 );
and ( n3468 , n2993 , n2996 );
or ( n3469 , n3467 , n3468 );
xor ( n3470 , n3466 , n3469 );
buf ( n3471 , n3470 );
buf ( n3472 , n3471 );
not ( n3473 , n3472 );
buf ( n3474 , n259 );
not ( n3475 , n3474 );
nor ( n3476 , n3473 , n3475 );
xor ( n3477 , n3168 , n3476 );
xor ( n3478 , n3013 , n3165 );
nor ( n3479 , n3000 , n3475 );
and ( n3480 , n3478 , n3479 );
xor ( n3481 , n3478 , n3479 );
xor ( n3482 , n3022 , n3163 );
nor ( n3483 , n2688 , n3475 );
and ( n3484 , n3482 , n3483 );
xor ( n3485 , n3482 , n3483 );
xor ( n3486 , n3031 , n3161 );
nor ( n3487 , n3008 , n3475 );
and ( n3488 , n3486 , n3487 );
xor ( n3489 , n3486 , n3487 );
xor ( n3490 , n3040 , n3159 );
nor ( n3491 , n3017 , n3475 );
and ( n3492 , n3490 , n3491 );
xor ( n3493 , n3490 , n3491 );
xor ( n3494 , n3049 , n3157 );
nor ( n3495 , n3026 , n3475 );
and ( n3496 , n3494 , n3495 );
xor ( n3497 , n3494 , n3495 );
xor ( n3498 , n3058 , n3155 );
nor ( n3499 , n3035 , n3475 );
and ( n3500 , n3498 , n3499 );
xor ( n3501 , n3498 , n3499 );
xor ( n3502 , n3067 , n3153 );
nor ( n3503 , n3044 , n3475 );
and ( n3504 , n3502 , n3503 );
xor ( n3505 , n3502 , n3503 );
xor ( n3506 , n3076 , n3151 );
nor ( n3507 , n3053 , n3475 );
and ( n3508 , n3506 , n3507 );
xor ( n3509 , n3506 , n3507 );
xor ( n3510 , n3085 , n3149 );
nor ( n3511 , n3062 , n3475 );
and ( n3512 , n3510 , n3511 );
xor ( n3513 , n3510 , n3511 );
xor ( n3514 , n3094 , n3147 );
nor ( n3515 , n3071 , n3475 );
and ( n3516 , n3514 , n3515 );
xor ( n3517 , n3514 , n3515 );
xor ( n3518 , n3103 , n3145 );
nor ( n3519 , n3080 , n3475 );
and ( n3520 , n3518 , n3519 );
xor ( n3521 , n3518 , n3519 );
xor ( n3522 , n3112 , n3143 );
nor ( n3523 , n3089 , n3475 );
and ( n3524 , n3522 , n3523 );
xor ( n3525 , n3522 , n3523 );
xor ( n3526 , n3121 , n3141 );
nor ( n3527 , n3098 , n3475 );
and ( n3528 , n3526 , n3527 );
xor ( n3529 , n3526 , n3527 );
xor ( n3530 , n3130 , n3139 );
nor ( n3531 , n3107 , n3475 );
and ( n3532 , n3530 , n3531 );
xor ( n3533 , n3530 , n3531 );
xor ( n3534 , n3136 , n3137 );
buf ( n3535 , n3534 );
nor ( n3536 , n3116 , n3475 );
and ( n3537 , n3535 , n3536 );
xor ( n3538 , n3535 , n3536 );
nor ( n3539 , n3134 , n3002 );
buf ( n3540 , n3539 );
nor ( n3541 , n3125 , n3475 );
and ( n3542 , n3540 , n3541 );
buf ( n3543 , n3542 );
and ( n3544 , n3538 , n3543 );
or ( n3545 , n3537 , n3544 );
and ( n3546 , n3533 , n3545 );
or ( n3547 , n3532 , n3546 );
and ( n3548 , n3529 , n3547 );
or ( n3549 , n3528 , n3548 );
and ( n3550 , n3525 , n3549 );
or ( n3551 , n3524 , n3550 );
and ( n3552 , n3521 , n3551 );
or ( n3553 , n3520 , n3552 );
and ( n3554 , n3517 , n3553 );
or ( n3555 , n3516 , n3554 );
and ( n3556 , n3513 , n3555 );
or ( n3557 , n3512 , n3556 );
and ( n3558 , n3509 , n3557 );
or ( n3559 , n3508 , n3558 );
and ( n3560 , n3505 , n3559 );
or ( n3561 , n3504 , n3560 );
and ( n3562 , n3501 , n3561 );
or ( n3563 , n3500 , n3562 );
and ( n3564 , n3497 , n3563 );
or ( n3565 , n3496 , n3564 );
and ( n3566 , n3493 , n3565 );
or ( n3567 , n3492 , n3566 );
and ( n3568 , n3489 , n3567 );
or ( n3569 , n3488 , n3568 );
and ( n3570 , n3485 , n3569 );
or ( n3571 , n3484 , n3570 );
and ( n3572 , n3481 , n3571 );
or ( n3573 , n3480 , n3572 );
xor ( n3574 , n3477 , n3573 );
and ( n3575 , n285 , n383 );
nor ( n3576 , n384 , n3575 );
nor ( n3577 , n456 , n305 );
xor ( n3578 , n3576 , n3577 );
and ( n3579 , n3170 , n3171 );
and ( n3580 , n3172 , n3175 );
or ( n3581 , n3579 , n3580 );
xor ( n3582 , n3578 , n3581 );
nor ( n3583 , n549 , n336 );
xor ( n3584 , n3582 , n3583 );
and ( n3585 , n3176 , n3177 );
and ( n3586 , n3178 , n3181 );
or ( n3587 , n3585 , n3586 );
xor ( n3588 , n3584 , n3587 );
nor ( n3589 , n663 , n386 );
xor ( n3590 , n3588 , n3589 );
and ( n3591 , n3182 , n3183 );
and ( n3592 , n3184 , n3187 );
or ( n3593 , n3591 , n3592 );
xor ( n3594 , n3590 , n3593 );
nor ( n3595 , n795 , n458 );
xor ( n3596 , n3594 , n3595 );
and ( n3597 , n3188 , n3189 );
and ( n3598 , n3190 , n3193 );
or ( n3599 , n3597 , n3598 );
xor ( n3600 , n3596 , n3599 );
nor ( n3601 , n952 , n551 );
xor ( n3602 , n3600 , n3601 );
and ( n3603 , n3194 , n3195 );
and ( n3604 , n3196 , n3199 );
or ( n3605 , n3603 , n3604 );
xor ( n3606 , n3602 , n3605 );
nor ( n3607 , n1126 , n665 );
xor ( n3608 , n3606 , n3607 );
and ( n3609 , n3200 , n3201 );
and ( n3610 , n3202 , n3205 );
or ( n3611 , n3609 , n3610 );
xor ( n3612 , n3608 , n3611 );
nor ( n3613 , n1318 , n797 );
xor ( n3614 , n3612 , n3613 );
and ( n3615 , n3206 , n3207 );
and ( n3616 , n3208 , n3211 );
or ( n3617 , n3615 , n3616 );
xor ( n3618 , n3614 , n3617 );
nor ( n3619 , n1534 , n954 );
xor ( n3620 , n3618 , n3619 );
and ( n3621 , n3212 , n3213 );
and ( n3622 , n3214 , n3217 );
or ( n3623 , n3621 , n3622 );
xor ( n3624 , n3620 , n3623 );
nor ( n3625 , n1771 , n1128 );
xor ( n3626 , n3624 , n3625 );
and ( n3627 , n3218 , n3219 );
and ( n3628 , n3220 , n3223 );
or ( n3629 , n3627 , n3628 );
xor ( n3630 , n3626 , n3629 );
nor ( n3631 , n2025 , n1320 );
xor ( n3632 , n3630 , n3631 );
and ( n3633 , n3224 , n3225 );
and ( n3634 , n3226 , n3229 );
or ( n3635 , n3633 , n3634 );
xor ( n3636 , n3632 , n3635 );
nor ( n3637 , n2300 , n1536 );
xor ( n3638 , n3636 , n3637 );
and ( n3639 , n3230 , n3231 );
and ( n3640 , n3232 , n3235 );
or ( n3641 , n3639 , n3640 );
xor ( n3642 , n3638 , n3641 );
nor ( n3643 , n2596 , n1773 );
xor ( n3644 , n3642 , n3643 );
and ( n3645 , n3236 , n3237 );
and ( n3646 , n3238 , n3241 );
or ( n3647 , n3645 , n3646 );
xor ( n3648 , n3644 , n3647 );
nor ( n3649 , n2991 , n2027 );
xor ( n3650 , n3648 , n3649 );
and ( n3651 , n3242 , n3243 );
and ( n3652 , n3244 , n3247 );
or ( n3653 , n3651 , n3652 );
xor ( n3654 , n3650 , n3653 );
nor ( n3655 , n3464 , n2302 );
xor ( n3656 , n3654 , n3655 );
and ( n3657 , n3248 , n3249 );
and ( n3658 , n3250 , n3253 );
or ( n3659 , n3657 , n3658 );
xor ( n3660 , n3656 , n3659 );
and ( n3661 , n3271 , n3275 );
and ( n3662 , n3275 , n3279 );
and ( n3663 , n3271 , n3279 );
or ( n3664 , n3661 , n3662 , n3663 );
and ( n3665 , n3267 , n3280 );
and ( n3666 , n3280 , n3450 );
and ( n3667 , n3267 , n3450 );
or ( n3668 , n3665 , n3666 , n3667 );
xor ( n3669 , n3664 , n3668 );
and ( n3670 , n3285 , n3311 );
and ( n3671 , n3311 , n3449 );
and ( n3672 , n3285 , n3449 );
or ( n3673 , n3670 , n3671 , n3672 );
and ( n3674 , n3299 , n3300 );
and ( n3675 , n3300 , n3302 );
and ( n3676 , n3299 , n3302 );
or ( n3677 , n3674 , n3675 , n3676 );
and ( n3678 , n3289 , n3293 );
and ( n3679 , n3293 , n3310 );
and ( n3680 , n3289 , n3310 );
or ( n3681 , n3678 , n3679 , n3680 );
xor ( n3682 , n3677 , n3681 );
not ( n3683 , n371 );
and ( n3684 , n2406 , n371 );
nor ( n3685 , n3683 , n3684 );
xor ( n3686 , n3682 , n3685 );
xor ( n3687 , n3673 , n3686 );
and ( n3688 , n3316 , n3331 );
and ( n3689 , n3331 , n3448 );
and ( n3690 , n3316 , n3448 );
or ( n3691 , n3688 , n3689 , n3690 );
and ( n3692 , n3298 , n3303 );
and ( n3693 , n3303 , n3309 );
and ( n3694 , n3298 , n3309 );
or ( n3695 , n3692 , n3693 , n3694 );
and ( n3696 , n3320 , n3324 );
and ( n3697 , n3324 , n3330 );
and ( n3698 , n3320 , n3330 );
or ( n3699 , n3696 , n3697 , n3698 );
xor ( n3700 , n3695 , n3699 );
and ( n3701 , n3305 , n3306 );
and ( n3702 , n3306 , n3308 );
and ( n3703 , n3305 , n3308 );
or ( n3704 , n3701 , n3702 , n3703 );
and ( n3705 , n446 , n2138 );
and ( n3706 , n533 , n1864 );
xor ( n3707 , n3705 , n3706 );
and ( n3708 , n636 , n1753 );
xor ( n3709 , n3707 , n3708 );
xor ( n3710 , n3704 , n3709 );
and ( n3711 , n782 , n1396 );
and ( n3712 , n931 , n1302 );
xor ( n3713 , n3711 , n3712 );
and ( n3714 , n1088 , n1114 );
xor ( n3715 , n3713 , n3714 );
xor ( n3716 , n3710 , n3715 );
xor ( n3717 , n3700 , n3716 );
xor ( n3718 , n3691 , n3717 );
and ( n3719 , n3336 , n3341 );
and ( n3720 , n3341 , n3447 );
and ( n3721 , n3336 , n3447 );
or ( n3722 , n3719 , n3720 , n3721 );
and ( n3723 , n3326 , n3327 );
and ( n3724 , n3327 , n3329 );
and ( n3725 , n3326 , n3329 );
or ( n3726 , n3723 , n3724 , n3725 );
and ( n3727 , n3337 , n3338 );
and ( n3728 , n3338 , n3340 );
and ( n3729 , n3337 , n3340 );
or ( n3730 , n3727 , n3728 , n3729 );
xor ( n3731 , n3726 , n3730 );
and ( n3732 , n1292 , n852 );
and ( n3733 , n1516 , n714 );
xor ( n3734 , n3732 , n3733 );
and ( n3735 , n1730 , n651 );
xor ( n3736 , n3734 , n3735 );
xor ( n3737 , n3731 , n3736 );
xor ( n3738 , n3722 , n3737 );
and ( n3739 , n3343 , n3344 );
and ( n3740 , n3344 , n3446 );
and ( n3741 , n3343 , n3446 );
or ( n3742 , n3739 , n3740 , n3741 );
and ( n3743 , n2001 , n488 );
and ( n3744 , n2286 , n411 );
xor ( n3745 , n3743 , n3744 );
and ( n3746 , n2581 , n375 );
xor ( n3747 , n3745 , n3746 );
xor ( n3748 , n3742 , n3747 );
and ( n3749 , n2972 , n312 );
and ( n3750 , n3445 , n288 );
xor ( n3751 , n3749 , n3750 );
and ( n3752 , n3362 , n3366 );
and ( n3753 , n3366 , n3370 );
and ( n3754 , n3362 , n3370 );
or ( n3755 , n3752 , n3753 , n3754 );
and ( n3756 , n3358 , n3371 );
and ( n3757 , n3371 , n3432 );
and ( n3758 , n3358 , n3432 );
or ( n3759 , n3756 , n3757 , n3758 );
xor ( n3760 , n3755 , n3759 );
and ( n3761 , n3376 , n3402 );
and ( n3762 , n3402 , n3431 );
and ( n3763 , n3376 , n3431 );
or ( n3764 , n3761 , n3762 , n3763 );
and ( n3765 , n3396 , n3397 );
and ( n3766 , n3397 , n3399 );
and ( n3767 , n3396 , n3399 );
or ( n3768 , n3765 , n3766 , n3767 );
and ( n3769 , n3380 , n3384 );
and ( n3770 , n3384 , n3401 );
and ( n3771 , n3380 , n3401 );
or ( n3772 , n3769 , n3770 , n3771 );
xor ( n3773 , n3768 , n3772 );
and ( n3774 , n2206 , n435 );
not ( n3775 , n435 );
nor ( n3776 , n3774 , n3775 );
xor ( n3777 , n3773 , n3776 );
xor ( n3778 , n3764 , n3777 );
and ( n3779 , n3407 , n3414 );
and ( n3780 , n3414 , n3430 );
and ( n3781 , n3407 , n3430 );
or ( n3782 , n3779 , n3780 , n3781 );
and ( n3783 , n3389 , n3394 );
and ( n3784 , n3394 , n3400 );
and ( n3785 , n3389 , n3400 );
or ( n3786 , n3783 , n3784 , n3785 );
and ( n3787 , n3419 , n3423 );
and ( n3788 , n3423 , n3429 );
and ( n3789 , n3419 , n3429 );
or ( n3790 , n3787 , n3788 , n3789 );
xor ( n3791 , n3786 , n3790 );
and ( n3792 , n3390 , n3391 );
and ( n3793 , n3391 , n3393 );
and ( n3794 , n3390 , n3393 );
or ( n3795 , n3792 , n3793 , n3794 );
and ( n3796 , n917 , n1261 );
and ( n3797 , n1077 , n1048 );
xor ( n3798 , n3796 , n3797 );
and ( n3799 , n1277 , n905 );
xor ( n3800 , n3798 , n3799 );
xor ( n3801 , n3795 , n3800 );
and ( n3802 , n1458 , n766 );
and ( n3803 , n1713 , n607 );
xor ( n3804 , n3802 , n3803 );
and ( n3805 , n1935 , n510 );
xor ( n3806 , n3804 , n3805 );
xor ( n3807 , n3801 , n3806 );
xor ( n3808 , n3791 , n3807 );
xor ( n3809 , n3782 , n3808 );
and ( n3810 , n3410 , n3411 );
and ( n3811 , n3411 , n3413 );
and ( n3812 , n3410 , n3413 );
or ( n3813 , n3810 , n3811 , n3812 );
and ( n3814 , n3425 , n3426 );
and ( n3815 , n3426 , n3428 );
and ( n3816 , n3425 , n3428 );
or ( n3817 , n3814 , n3815 , n3816 );
xor ( n3818 , n3813 , n3817 );
and ( n3819 , n521 , n1975 );
and ( n3820 , n625 , n1685 );
xor ( n3821 , n3819 , n3820 );
and ( n3822 , n753 , n1497 );
xor ( n3823 , n3821 , n3822 );
xor ( n3824 , n3818 , n3823 );
not ( n3825 , n361 );
and ( n3826 , n2563 , n361 );
nor ( n3827 , n3825 , n3826 );
and ( n3828 , n431 , n2271 );
xor ( n3829 , n3827 , n3828 );
xor ( n3830 , n3824 , n3829 );
xor ( n3831 , n3809 , n3830 );
xor ( n3832 , n3778 , n3831 );
xor ( n3833 , n3760 , n3832 );
and ( n3834 , n3349 , n3353 );
and ( n3835 , n3353 , n3433 );
and ( n3836 , n3349 , n3433 );
or ( n3837 , n3834 , n3835 , n3836 );
xor ( n3838 , n3833 , n3837 );
and ( n3839 , n3434 , n3438 );
and ( n3840 , n3439 , n3442 );
or ( n3841 , n3839 , n3840 );
xor ( n3842 , n3838 , n3841 );
buf ( n3843 , n3842 );
buf ( n3844 , n3843 );
and ( n3845 , n3844 , n279 );
xor ( n3846 , n3751 , n3845 );
xor ( n3847 , n3748 , n3846 );
xor ( n3848 , n3738 , n3847 );
xor ( n3849 , n3718 , n3848 );
xor ( n3850 , n3687 , n3849 );
xor ( n3851 , n3669 , n3850 );
and ( n3852 , n3258 , n3262 );
and ( n3853 , n3262 , n3451 );
and ( n3854 , n3258 , n3451 );
or ( n3855 , n3852 , n3853 , n3854 );
xor ( n3856 , n3851 , n3855 );
and ( n3857 , n3452 , n3456 );
and ( n3858 , n3457 , n3460 );
or ( n3859 , n3857 , n3858 );
xor ( n3860 , n3856 , n3859 );
buf ( n3861 , n3860 );
buf ( n3862 , n3861 );
not ( n3863 , n3862 );
nor ( n3864 , n3863 , n2598 );
xor ( n3865 , n3660 , n3864 );
and ( n3866 , n3254 , n3465 );
and ( n3867 , n3466 , n3469 );
or ( n3868 , n3866 , n3867 );
xor ( n3869 , n3865 , n3868 );
buf ( n3870 , n3869 );
buf ( n3871 , n3870 );
not ( n3872 , n3871 );
buf ( n3873 , n260 );
not ( n3874 , n3873 );
nor ( n3875 , n3872 , n3874 );
xor ( n3876 , n3574 , n3875 );
xor ( n3877 , n3481 , n3571 );
nor ( n3878 , n3473 , n3874 );
and ( n3879 , n3877 , n3878 );
xor ( n3880 , n3877 , n3878 );
xor ( n3881 , n3485 , n3569 );
nor ( n3882 , n3000 , n3874 );
and ( n3883 , n3881 , n3882 );
xor ( n3884 , n3881 , n3882 );
xor ( n3885 , n3489 , n3567 );
nor ( n3886 , n2688 , n3874 );
and ( n3887 , n3885 , n3886 );
xor ( n3888 , n3885 , n3886 );
xor ( n3889 , n3493 , n3565 );
nor ( n3890 , n3008 , n3874 );
and ( n3891 , n3889 , n3890 );
xor ( n3892 , n3889 , n3890 );
xor ( n3893 , n3497 , n3563 );
nor ( n3894 , n3017 , n3874 );
and ( n3895 , n3893 , n3894 );
xor ( n3896 , n3893 , n3894 );
xor ( n3897 , n3501 , n3561 );
nor ( n3898 , n3026 , n3874 );
and ( n3899 , n3897 , n3898 );
xor ( n3900 , n3897 , n3898 );
xor ( n3901 , n3505 , n3559 );
nor ( n3902 , n3035 , n3874 );
and ( n3903 , n3901 , n3902 );
xor ( n3904 , n3901 , n3902 );
xor ( n3905 , n3509 , n3557 );
nor ( n3906 , n3044 , n3874 );
and ( n3907 , n3905 , n3906 );
xor ( n3908 , n3905 , n3906 );
xor ( n3909 , n3513 , n3555 );
nor ( n3910 , n3053 , n3874 );
and ( n3911 , n3909 , n3910 );
xor ( n3912 , n3909 , n3910 );
xor ( n3913 , n3517 , n3553 );
nor ( n3914 , n3062 , n3874 );
and ( n3915 , n3913 , n3914 );
xor ( n3916 , n3913 , n3914 );
xor ( n3917 , n3521 , n3551 );
nor ( n3918 , n3071 , n3874 );
and ( n3919 , n3917 , n3918 );
xor ( n3920 , n3917 , n3918 );
xor ( n3921 , n3525 , n3549 );
nor ( n3922 , n3080 , n3874 );
and ( n3923 , n3921 , n3922 );
xor ( n3924 , n3921 , n3922 );
xor ( n3925 , n3529 , n3547 );
nor ( n3926 , n3089 , n3874 );
and ( n3927 , n3925 , n3926 );
xor ( n3928 , n3925 , n3926 );
xor ( n3929 , n3533 , n3545 );
nor ( n3930 , n3098 , n3874 );
and ( n3931 , n3929 , n3930 );
xor ( n3932 , n3929 , n3930 );
xor ( n3933 , n3538 , n3543 );
nor ( n3934 , n3107 , n3874 );
and ( n3935 , n3933 , n3934 );
xor ( n3936 , n3933 , n3934 );
xor ( n3937 , n3540 , n3541 );
buf ( n3938 , n3937 );
nor ( n3939 , n3116 , n3874 );
and ( n3940 , n3938 , n3939 );
xor ( n3941 , n3938 , n3939 );
nor ( n3942 , n3134 , n3475 );
buf ( n3943 , n3942 );
nor ( n3944 , n3125 , n3874 );
and ( n3945 , n3943 , n3944 );
buf ( n3946 , n3945 );
and ( n3947 , n3941 , n3946 );
or ( n3948 , n3940 , n3947 );
and ( n3949 , n3936 , n3948 );
or ( n3950 , n3935 , n3949 );
and ( n3951 , n3932 , n3950 );
or ( n3952 , n3931 , n3951 );
and ( n3953 , n3928 , n3952 );
or ( n3954 , n3927 , n3953 );
and ( n3955 , n3924 , n3954 );
or ( n3956 , n3923 , n3955 );
and ( n3957 , n3920 , n3956 );
or ( n3958 , n3919 , n3957 );
and ( n3959 , n3916 , n3958 );
or ( n3960 , n3915 , n3959 );
and ( n3961 , n3912 , n3960 );
or ( n3962 , n3911 , n3961 );
and ( n3963 , n3908 , n3962 );
or ( n3964 , n3907 , n3963 );
and ( n3965 , n3904 , n3964 );
or ( n3966 , n3903 , n3965 );
and ( n3967 , n3900 , n3966 );
or ( n3968 , n3899 , n3967 );
and ( n3969 , n3896 , n3968 );
or ( n3970 , n3895 , n3969 );
and ( n3971 , n3892 , n3970 );
or ( n3972 , n3891 , n3971 );
and ( n3973 , n3888 , n3972 );
or ( n3974 , n3887 , n3973 );
and ( n3975 , n3884 , n3974 );
or ( n3976 , n3883 , n3975 );
and ( n3977 , n3880 , n3976 );
or ( n3978 , n3879 , n3977 );
xor ( n3979 , n3876 , n3978 );
and ( n3980 , n285 , n455 );
nor ( n3981 , n456 , n3980 );
nor ( n3982 , n549 , n305 );
xor ( n3983 , n3981 , n3982 );
and ( n3984 , n3576 , n3577 );
and ( n3985 , n3578 , n3581 );
or ( n3986 , n3984 , n3985 );
xor ( n3987 , n3983 , n3986 );
nor ( n3988 , n663 , n336 );
xor ( n3989 , n3987 , n3988 );
and ( n3990 , n3582 , n3583 );
and ( n3991 , n3584 , n3587 );
or ( n3992 , n3990 , n3991 );
xor ( n3993 , n3989 , n3992 );
nor ( n3994 , n795 , n386 );
xor ( n3995 , n3993 , n3994 );
and ( n3996 , n3588 , n3589 );
and ( n3997 , n3590 , n3593 );
or ( n3998 , n3996 , n3997 );
xor ( n3999 , n3995 , n3998 );
nor ( n4000 , n952 , n458 );
xor ( n4001 , n3999 , n4000 );
and ( n4002 , n3594 , n3595 );
and ( n4003 , n3596 , n3599 );
or ( n4004 , n4002 , n4003 );
xor ( n4005 , n4001 , n4004 );
nor ( n4006 , n1126 , n551 );
xor ( n4007 , n4005 , n4006 );
and ( n4008 , n3600 , n3601 );
and ( n4009 , n3602 , n3605 );
or ( n4010 , n4008 , n4009 );
xor ( n4011 , n4007 , n4010 );
nor ( n4012 , n1318 , n665 );
xor ( n4013 , n4011 , n4012 );
and ( n4014 , n3606 , n3607 );
and ( n4015 , n3608 , n3611 );
or ( n4016 , n4014 , n4015 );
xor ( n4017 , n4013 , n4016 );
nor ( n4018 , n1534 , n797 );
xor ( n4019 , n4017 , n4018 );
and ( n4020 , n3612 , n3613 );
and ( n4021 , n3614 , n3617 );
or ( n4022 , n4020 , n4021 );
xor ( n4023 , n4019 , n4022 );
nor ( n4024 , n1771 , n954 );
xor ( n4025 , n4023 , n4024 );
and ( n4026 , n3618 , n3619 );
and ( n4027 , n3620 , n3623 );
or ( n4028 , n4026 , n4027 );
xor ( n4029 , n4025 , n4028 );
nor ( n4030 , n2025 , n1128 );
xor ( n4031 , n4029 , n4030 );
and ( n4032 , n3624 , n3625 );
and ( n4033 , n3626 , n3629 );
or ( n4034 , n4032 , n4033 );
xor ( n4035 , n4031 , n4034 );
nor ( n4036 , n2300 , n1320 );
xor ( n4037 , n4035 , n4036 );
and ( n4038 , n3630 , n3631 );
and ( n4039 , n3632 , n3635 );
or ( n4040 , n4038 , n4039 );
xor ( n4041 , n4037 , n4040 );
nor ( n4042 , n2596 , n1536 );
xor ( n4043 , n4041 , n4042 );
and ( n4044 , n3636 , n3637 );
and ( n4045 , n3638 , n3641 );
or ( n4046 , n4044 , n4045 );
xor ( n4047 , n4043 , n4046 );
nor ( n4048 , n2991 , n1773 );
xor ( n4049 , n4047 , n4048 );
and ( n4050 , n3642 , n3643 );
and ( n4051 , n3644 , n3647 );
or ( n4052 , n4050 , n4051 );
xor ( n4053 , n4049 , n4052 );
nor ( n4054 , n3464 , n2027 );
xor ( n4055 , n4053 , n4054 );
and ( n4056 , n3648 , n3649 );
and ( n4057 , n3650 , n3653 );
or ( n4058 , n4056 , n4057 );
xor ( n4059 , n4055 , n4058 );
nor ( n4060 , n3863 , n2302 );
xor ( n4061 , n4059 , n4060 );
and ( n4062 , n3654 , n3655 );
and ( n4063 , n3656 , n3659 );
or ( n4064 , n4062 , n4063 );
xor ( n4065 , n4061 , n4064 );
and ( n4066 , n3677 , n3681 );
and ( n4067 , n3681 , n3685 );
and ( n4068 , n3677 , n3685 );
or ( n4069 , n4066 , n4067 , n4068 );
and ( n4070 , n3673 , n3686 );
and ( n4071 , n3686 , n3849 );
and ( n4072 , n3673 , n3849 );
or ( n4073 , n4070 , n4071 , n4072 );
xor ( n4074 , n4069 , n4073 );
and ( n4075 , n3691 , n3717 );
and ( n4076 , n3717 , n3848 );
and ( n4077 , n3691 , n3848 );
or ( n4078 , n4075 , n4076 , n4077 );
and ( n4079 , n3705 , n3706 );
and ( n4080 , n3706 , n3708 );
and ( n4081 , n3705 , n3708 );
or ( n4082 , n4079 , n4080 , n4081 );
and ( n4083 , n3695 , n3699 );
and ( n4084 , n3699 , n3716 );
and ( n4085 , n3695 , n3716 );
or ( n4086 , n4083 , n4084 , n4085 );
xor ( n4087 , n4082 , n4086 );
not ( n4088 , n446 );
and ( n4089 , n2406 , n446 );
nor ( n4090 , n4088 , n4089 );
xor ( n4091 , n4087 , n4090 );
xor ( n4092 , n4078 , n4091 );
and ( n4093 , n3722 , n3737 );
and ( n4094 , n3737 , n3847 );
and ( n4095 , n3722 , n3847 );
or ( n4096 , n4093 , n4094 , n4095 );
and ( n4097 , n3704 , n3709 );
and ( n4098 , n3709 , n3715 );
and ( n4099 , n3704 , n3715 );
or ( n4100 , n4097 , n4098 , n4099 );
and ( n4101 , n3726 , n3730 );
and ( n4102 , n3730 , n3736 );
and ( n4103 , n3726 , n3736 );
or ( n4104 , n4101 , n4102 , n4103 );
xor ( n4105 , n4100 , n4104 );
and ( n4106 , n3711 , n3712 );
and ( n4107 , n3712 , n3714 );
and ( n4108 , n3711 , n3714 );
or ( n4109 , n4106 , n4107 , n4108 );
and ( n4110 , n533 , n2138 );
and ( n4111 , n636 , n1864 );
xor ( n4112 , n4110 , n4111 );
and ( n4113 , n782 , n1753 );
xor ( n4114 , n4112 , n4113 );
xor ( n4115 , n4109 , n4114 );
and ( n4116 , n931 , n1396 );
and ( n4117 , n1088 , n1302 );
xor ( n4118 , n4116 , n4117 );
and ( n4119 , n1292 , n1114 );
xor ( n4120 , n4118 , n4119 );
xor ( n4121 , n4115 , n4120 );
xor ( n4122 , n4105 , n4121 );
xor ( n4123 , n4096 , n4122 );
and ( n4124 , n3742 , n3747 );
and ( n4125 , n3747 , n3846 );
and ( n4126 , n3742 , n3846 );
or ( n4127 , n4124 , n4125 , n4126 );
and ( n4128 , n3732 , n3733 );
and ( n4129 , n3733 , n3735 );
and ( n4130 , n3732 , n3735 );
or ( n4131 , n4128 , n4129 , n4130 );
and ( n4132 , n3743 , n3744 );
and ( n4133 , n3744 , n3746 );
and ( n4134 , n3743 , n3746 );
or ( n4135 , n4132 , n4133 , n4134 );
xor ( n4136 , n4131 , n4135 );
and ( n4137 , n1516 , n852 );
and ( n4138 , n1730 , n714 );
xor ( n4139 , n4137 , n4138 );
and ( n4140 , n2001 , n651 );
xor ( n4141 , n4139 , n4140 );
xor ( n4142 , n4136 , n4141 );
xor ( n4143 , n4127 , n4142 );
and ( n4144 , n3749 , n3750 );
and ( n4145 , n3750 , n3845 );
and ( n4146 , n3749 , n3845 );
or ( n4147 , n4144 , n4145 , n4146 );
and ( n4148 , n2286 , n488 );
and ( n4149 , n2581 , n411 );
xor ( n4150 , n4148 , n4149 );
and ( n4151 , n2972 , n375 );
xor ( n4152 , n4150 , n4151 );
xor ( n4153 , n4147 , n4152 );
and ( n4154 , n3445 , n312 );
and ( n4155 , n3844 , n288 );
xor ( n4156 , n4154 , n4155 );
and ( n4157 , n3768 , n3772 );
and ( n4158 , n3772 , n3776 );
and ( n4159 , n3768 , n3776 );
or ( n4160 , n4157 , n4158 , n4159 );
and ( n4161 , n3764 , n3777 );
and ( n4162 , n3777 , n3831 );
and ( n4163 , n3764 , n3831 );
or ( n4164 , n4161 , n4162 , n4163 );
xor ( n4165 , n4160 , n4164 );
and ( n4166 , n3782 , n3808 );
and ( n4167 , n3808 , n3830 );
and ( n4168 , n3782 , n3830 );
or ( n4169 , n4166 , n4167 , n4168 );
and ( n4170 , n3802 , n3803 );
and ( n4171 , n3803 , n3805 );
and ( n4172 , n3802 , n3805 );
or ( n4173 , n4170 , n4171 , n4172 );
and ( n4174 , n3786 , n3790 );
and ( n4175 , n3790 , n3807 );
and ( n4176 , n3786 , n3807 );
or ( n4177 , n4174 , n4175 , n4176 );
xor ( n4178 , n4173 , n4177 );
and ( n4179 , n2206 , n510 );
not ( n4180 , n510 );
nor ( n4181 , n4179 , n4180 );
xor ( n4182 , n4178 , n4181 );
xor ( n4183 , n4169 , n4182 );
and ( n4184 , n3824 , n3829 );
and ( n4185 , n3813 , n3817 );
and ( n4186 , n3817 , n3823 );
and ( n4187 , n3813 , n3823 );
or ( n4188 , n4185 , n4186 , n4187 );
and ( n4189 , n3795 , n3800 );
and ( n4190 , n3800 , n3806 );
and ( n4191 , n3795 , n3806 );
or ( n4192 , n4189 , n4190 , n4191 );
xor ( n4193 , n4188 , n4192 );
and ( n4194 , n3796 , n3797 );
and ( n4195 , n3797 , n3799 );
and ( n4196 , n3796 , n3799 );
or ( n4197 , n4194 , n4195 , n4196 );
and ( n4198 , n917 , n1497 );
and ( n4199 , n1077 , n1261 );
xor ( n4200 , n4198 , n4199 );
and ( n4201 , n1277 , n1048 );
xor ( n4202 , n4200 , n4201 );
xor ( n4203 , n4197 , n4202 );
and ( n4204 , n1458 , n905 );
and ( n4205 , n1713 , n766 );
xor ( n4206 , n4204 , n4205 );
and ( n4207 , n1935 , n607 );
xor ( n4208 , n4206 , n4207 );
xor ( n4209 , n4203 , n4208 );
xor ( n4210 , n4193 , n4209 );
xor ( n4211 , n4184 , n4210 );
not ( n4212 , n431 );
and ( n4213 , n2563 , n431 );
nor ( n4214 , n4212 , n4213 );
and ( n4215 , n3819 , n3820 );
and ( n4216 , n3820 , n3822 );
and ( n4217 , n3819 , n3822 );
or ( n4218 , n4215 , n4216 , n4217 );
and ( n4219 , n3827 , n3828 );
xor ( n4220 , n4218 , n4219 );
and ( n4221 , n521 , n2271 );
and ( n4222 , n625 , n1975 );
xor ( n4223 , n4221 , n4222 );
and ( n4224 , n753 , n1685 );
xor ( n4225 , n4223 , n4224 );
xor ( n4226 , n4220 , n4225 );
xor ( n4227 , n4214 , n4226 );
xor ( n4228 , n4211 , n4227 );
xor ( n4229 , n4183 , n4228 );
xor ( n4230 , n4165 , n4229 );
and ( n4231 , n3755 , n3759 );
and ( n4232 , n3759 , n3832 );
and ( n4233 , n3755 , n3832 );
or ( n4234 , n4231 , n4232 , n4233 );
xor ( n4235 , n4230 , n4234 );
and ( n4236 , n3833 , n3837 );
and ( n4237 , n3838 , n3841 );
or ( n4238 , n4236 , n4237 );
xor ( n4239 , n4235 , n4238 );
buf ( n4240 , n4239 );
buf ( n4241 , n4240 );
and ( n4242 , n4241 , n279 );
xor ( n4243 , n4156 , n4242 );
xor ( n4244 , n4153 , n4243 );
xor ( n4245 , n4143 , n4244 );
xor ( n4246 , n4123 , n4245 );
xor ( n4247 , n4092 , n4246 );
xor ( n4248 , n4074 , n4247 );
and ( n4249 , n3664 , n3668 );
and ( n4250 , n3668 , n3850 );
and ( n4251 , n3664 , n3850 );
or ( n4252 , n4249 , n4250 , n4251 );
xor ( n4253 , n4248 , n4252 );
and ( n4254 , n3851 , n3855 );
and ( n4255 , n3856 , n3859 );
or ( n4256 , n4254 , n4255 );
xor ( n4257 , n4253 , n4256 );
buf ( n4258 , n4257 );
buf ( n4259 , n4258 );
not ( n4260 , n4259 );
nor ( n4261 , n4260 , n2598 );
xor ( n4262 , n4065 , n4261 );
and ( n4263 , n3660 , n3864 );
and ( n4264 , n3865 , n3868 );
or ( n4265 , n4263 , n4264 );
xor ( n4266 , n4262 , n4265 );
buf ( n4267 , n4266 );
buf ( n4268 , n4267 );
not ( n4269 , n4268 );
buf ( n4270 , n261 );
not ( n4271 , n4270 );
nor ( n4272 , n4269 , n4271 );
xor ( n4273 , n3979 , n4272 );
xor ( n4274 , n3880 , n3976 );
nor ( n4275 , n3872 , n4271 );
and ( n4276 , n4274 , n4275 );
xor ( n4277 , n4274 , n4275 );
xor ( n4278 , n3884 , n3974 );
nor ( n4279 , n3473 , n4271 );
and ( n4280 , n4278 , n4279 );
xor ( n4281 , n4278 , n4279 );
xor ( n4282 , n3888 , n3972 );
nor ( n4283 , n3000 , n4271 );
and ( n4284 , n4282 , n4283 );
xor ( n4285 , n4282 , n4283 );
xor ( n4286 , n3892 , n3970 );
nor ( n4287 , n2688 , n4271 );
and ( n4288 , n4286 , n4287 );
xor ( n4289 , n4286 , n4287 );
xor ( n4290 , n3896 , n3968 );
nor ( n4291 , n3008 , n4271 );
and ( n4292 , n4290 , n4291 );
xor ( n4293 , n4290 , n4291 );
xor ( n4294 , n3900 , n3966 );
nor ( n4295 , n3017 , n4271 );
and ( n4296 , n4294 , n4295 );
xor ( n4297 , n4294 , n4295 );
xor ( n4298 , n3904 , n3964 );
nor ( n4299 , n3026 , n4271 );
and ( n4300 , n4298 , n4299 );
xor ( n4301 , n4298 , n4299 );
xor ( n4302 , n3908 , n3962 );
nor ( n4303 , n3035 , n4271 );
and ( n4304 , n4302 , n4303 );
xor ( n4305 , n4302 , n4303 );
xor ( n4306 , n3912 , n3960 );
nor ( n4307 , n3044 , n4271 );
and ( n4308 , n4306 , n4307 );
xor ( n4309 , n4306 , n4307 );
xor ( n4310 , n3916 , n3958 );
nor ( n4311 , n3053 , n4271 );
and ( n4312 , n4310 , n4311 );
xor ( n4313 , n4310 , n4311 );
xor ( n4314 , n3920 , n3956 );
nor ( n4315 , n3062 , n4271 );
and ( n4316 , n4314 , n4315 );
xor ( n4317 , n4314 , n4315 );
xor ( n4318 , n3924 , n3954 );
nor ( n4319 , n3071 , n4271 );
and ( n4320 , n4318 , n4319 );
xor ( n4321 , n4318 , n4319 );
xor ( n4322 , n3928 , n3952 );
nor ( n4323 , n3080 , n4271 );
and ( n4324 , n4322 , n4323 );
xor ( n4325 , n4322 , n4323 );
xor ( n4326 , n3932 , n3950 );
nor ( n4327 , n3089 , n4271 );
and ( n4328 , n4326 , n4327 );
xor ( n4329 , n4326 , n4327 );
xor ( n4330 , n3936 , n3948 );
nor ( n4331 , n3098 , n4271 );
and ( n4332 , n4330 , n4331 );
xor ( n4333 , n4330 , n4331 );
xor ( n4334 , n3941 , n3946 );
nor ( n4335 , n3107 , n4271 );
and ( n4336 , n4334 , n4335 );
xor ( n4337 , n4334 , n4335 );
xor ( n4338 , n3943 , n3944 );
buf ( n4339 , n4338 );
nor ( n4340 , n3116 , n4271 );
and ( n4341 , n4339 , n4340 );
xor ( n4342 , n4339 , n4340 );
nor ( n4343 , n3134 , n3874 );
buf ( n4344 , n4343 );
nor ( n4345 , n3125 , n4271 );
and ( n4346 , n4344 , n4345 );
buf ( n4347 , n4346 );
and ( n4348 , n4342 , n4347 );
or ( n4349 , n4341 , n4348 );
and ( n4350 , n4337 , n4349 );
or ( n4351 , n4336 , n4350 );
and ( n4352 , n4333 , n4351 );
or ( n4353 , n4332 , n4352 );
and ( n4354 , n4329 , n4353 );
or ( n4355 , n4328 , n4354 );
and ( n4356 , n4325 , n4355 );
or ( n4357 , n4324 , n4356 );
and ( n4358 , n4321 , n4357 );
or ( n4359 , n4320 , n4358 );
and ( n4360 , n4317 , n4359 );
or ( n4361 , n4316 , n4360 );
and ( n4362 , n4313 , n4361 );
or ( n4363 , n4312 , n4362 );
and ( n4364 , n4309 , n4363 );
or ( n4365 , n4308 , n4364 );
and ( n4366 , n4305 , n4365 );
or ( n4367 , n4304 , n4366 );
and ( n4368 , n4301 , n4367 );
or ( n4369 , n4300 , n4368 );
and ( n4370 , n4297 , n4369 );
or ( n4371 , n4296 , n4370 );
and ( n4372 , n4293 , n4371 );
or ( n4373 , n4292 , n4372 );
and ( n4374 , n4289 , n4373 );
or ( n4375 , n4288 , n4374 );
and ( n4376 , n4285 , n4375 );
or ( n4377 , n4284 , n4376 );
and ( n4378 , n4281 , n4377 );
or ( n4379 , n4280 , n4378 );
and ( n4380 , n4277 , n4379 );
or ( n4381 , n4276 , n4380 );
xor ( n4382 , n4273 , n4381 );
and ( n4383 , n285 , n548 );
nor ( n4384 , n549 , n4383 );
nor ( n4385 , n663 , n305 );
xor ( n4386 , n4384 , n4385 );
and ( n4387 , n3981 , n3982 );
and ( n4388 , n3983 , n3986 );
or ( n4389 , n4387 , n4388 );
xor ( n4390 , n4386 , n4389 );
nor ( n4391 , n795 , n336 );
xor ( n4392 , n4390 , n4391 );
and ( n4393 , n3987 , n3988 );
and ( n4394 , n3989 , n3992 );
or ( n4395 , n4393 , n4394 );
xor ( n4396 , n4392 , n4395 );
nor ( n4397 , n952 , n386 );
xor ( n4398 , n4396 , n4397 );
and ( n4399 , n3993 , n3994 );
and ( n4400 , n3995 , n3998 );
or ( n4401 , n4399 , n4400 );
xor ( n4402 , n4398 , n4401 );
nor ( n4403 , n1126 , n458 );
xor ( n4404 , n4402 , n4403 );
and ( n4405 , n3999 , n4000 );
and ( n4406 , n4001 , n4004 );
or ( n4407 , n4405 , n4406 );
xor ( n4408 , n4404 , n4407 );
nor ( n4409 , n1318 , n551 );
xor ( n4410 , n4408 , n4409 );
and ( n4411 , n4005 , n4006 );
and ( n4412 , n4007 , n4010 );
or ( n4413 , n4411 , n4412 );
xor ( n4414 , n4410 , n4413 );
nor ( n4415 , n1534 , n665 );
xor ( n4416 , n4414 , n4415 );
and ( n4417 , n4011 , n4012 );
and ( n4418 , n4013 , n4016 );
or ( n4419 , n4417 , n4418 );
xor ( n4420 , n4416 , n4419 );
nor ( n4421 , n1771 , n797 );
xor ( n4422 , n4420 , n4421 );
and ( n4423 , n4017 , n4018 );
and ( n4424 , n4019 , n4022 );
or ( n4425 , n4423 , n4424 );
xor ( n4426 , n4422 , n4425 );
nor ( n4427 , n2025 , n954 );
xor ( n4428 , n4426 , n4427 );
and ( n4429 , n4023 , n4024 );
and ( n4430 , n4025 , n4028 );
or ( n4431 , n4429 , n4430 );
xor ( n4432 , n4428 , n4431 );
nor ( n4433 , n2300 , n1128 );
xor ( n4434 , n4432 , n4433 );
and ( n4435 , n4029 , n4030 );
and ( n4436 , n4031 , n4034 );
or ( n4437 , n4435 , n4436 );
xor ( n4438 , n4434 , n4437 );
nor ( n4439 , n2596 , n1320 );
xor ( n4440 , n4438 , n4439 );
and ( n4441 , n4035 , n4036 );
and ( n4442 , n4037 , n4040 );
or ( n4443 , n4441 , n4442 );
xor ( n4444 , n4440 , n4443 );
nor ( n4445 , n2991 , n1536 );
xor ( n4446 , n4444 , n4445 );
and ( n4447 , n4041 , n4042 );
and ( n4448 , n4043 , n4046 );
or ( n4449 , n4447 , n4448 );
xor ( n4450 , n4446 , n4449 );
nor ( n4451 , n3464 , n1773 );
xor ( n4452 , n4450 , n4451 );
and ( n4453 , n4047 , n4048 );
and ( n4454 , n4049 , n4052 );
or ( n4455 , n4453 , n4454 );
xor ( n4456 , n4452 , n4455 );
nor ( n4457 , n3863 , n2027 );
xor ( n4458 , n4456 , n4457 );
and ( n4459 , n4053 , n4054 );
and ( n4460 , n4055 , n4058 );
or ( n4461 , n4459 , n4460 );
xor ( n4462 , n4458 , n4461 );
nor ( n4463 , n4260 , n2302 );
xor ( n4464 , n4462 , n4463 );
and ( n4465 , n4059 , n4060 );
and ( n4466 , n4061 , n4064 );
or ( n4467 , n4465 , n4466 );
xor ( n4468 , n4464 , n4467 );
and ( n4469 , n4082 , n4086 );
and ( n4470 , n4086 , n4090 );
and ( n4471 , n4082 , n4090 );
or ( n4472 , n4469 , n4470 , n4471 );
and ( n4473 , n4078 , n4091 );
and ( n4474 , n4091 , n4246 );
and ( n4475 , n4078 , n4246 );
or ( n4476 , n4473 , n4474 , n4475 );
xor ( n4477 , n4472 , n4476 );
and ( n4478 , n4096 , n4122 );
and ( n4479 , n4122 , n4245 );
and ( n4480 , n4096 , n4245 );
or ( n4481 , n4478 , n4479 , n4480 );
and ( n4482 , n4110 , n4111 );
and ( n4483 , n4111 , n4113 );
and ( n4484 , n4110 , n4113 );
or ( n4485 , n4482 , n4483 , n4484 );
and ( n4486 , n4100 , n4104 );
and ( n4487 , n4104 , n4121 );
and ( n4488 , n4100 , n4121 );
or ( n4489 , n4486 , n4487 , n4488 );
xor ( n4490 , n4485 , n4489 );
not ( n4491 , n533 );
and ( n4492 , n2406 , n533 );
nor ( n4493 , n4491 , n4492 );
xor ( n4494 , n4490 , n4493 );
xor ( n4495 , n4481 , n4494 );
and ( n4496 , n4127 , n4142 );
and ( n4497 , n4142 , n4244 );
and ( n4498 , n4127 , n4244 );
or ( n4499 , n4496 , n4497 , n4498 );
and ( n4500 , n4109 , n4114 );
and ( n4501 , n4114 , n4120 );
and ( n4502 , n4109 , n4120 );
or ( n4503 , n4500 , n4501 , n4502 );
and ( n4504 , n4131 , n4135 );
and ( n4505 , n4135 , n4141 );
and ( n4506 , n4131 , n4141 );
or ( n4507 , n4504 , n4505 , n4506 );
xor ( n4508 , n4503 , n4507 );
and ( n4509 , n4116 , n4117 );
and ( n4510 , n4117 , n4119 );
and ( n4511 , n4116 , n4119 );
or ( n4512 , n4509 , n4510 , n4511 );
and ( n4513 , n636 , n2138 );
and ( n4514 , n782 , n1864 );
xor ( n4515 , n4513 , n4514 );
and ( n4516 , n931 , n1753 );
xor ( n4517 , n4515 , n4516 );
xor ( n4518 , n4512 , n4517 );
and ( n4519 , n1088 , n1396 );
and ( n4520 , n1292 , n1302 );
xor ( n4521 , n4519 , n4520 );
and ( n4522 , n1516 , n1114 );
xor ( n4523 , n4521 , n4522 );
xor ( n4524 , n4518 , n4523 );
xor ( n4525 , n4508 , n4524 );
xor ( n4526 , n4499 , n4525 );
and ( n4527 , n4147 , n4152 );
and ( n4528 , n4152 , n4243 );
and ( n4529 , n4147 , n4243 );
or ( n4530 , n4527 , n4528 , n4529 );
and ( n4531 , n4137 , n4138 );
and ( n4532 , n4138 , n4140 );
and ( n4533 , n4137 , n4140 );
or ( n4534 , n4531 , n4532 , n4533 );
and ( n4535 , n4148 , n4149 );
and ( n4536 , n4149 , n4151 );
and ( n4537 , n4148 , n4151 );
or ( n4538 , n4535 , n4536 , n4537 );
xor ( n4539 , n4534 , n4538 );
and ( n4540 , n1730 , n852 );
and ( n4541 , n2001 , n714 );
xor ( n4542 , n4540 , n4541 );
and ( n4543 , n2286 , n651 );
xor ( n4544 , n4542 , n4543 );
xor ( n4545 , n4539 , n4544 );
xor ( n4546 , n4530 , n4545 );
and ( n4547 , n4154 , n4155 );
and ( n4548 , n4155 , n4242 );
and ( n4549 , n4154 , n4242 );
or ( n4550 , n4547 , n4548 , n4549 );
and ( n4551 , n2581 , n488 );
and ( n4552 , n2972 , n411 );
xor ( n4553 , n4551 , n4552 );
and ( n4554 , n3445 , n375 );
xor ( n4555 , n4553 , n4554 );
xor ( n4556 , n4550 , n4555 );
and ( n4557 , n3844 , n312 );
and ( n4558 , n4241 , n288 );
xor ( n4559 , n4557 , n4558 );
and ( n4560 , n4173 , n4177 );
and ( n4561 , n4177 , n4181 );
and ( n4562 , n4173 , n4181 );
or ( n4563 , n4560 , n4561 , n4562 );
and ( n4564 , n4169 , n4182 );
and ( n4565 , n4182 , n4228 );
and ( n4566 , n4169 , n4228 );
or ( n4567 , n4564 , n4565 , n4566 );
xor ( n4568 , n4563 , n4567 );
and ( n4569 , n4184 , n4210 );
and ( n4570 , n4210 , n4227 );
and ( n4571 , n4184 , n4227 );
or ( n4572 , n4569 , n4570 , n4571 );
and ( n4573 , n4204 , n4205 );
and ( n4574 , n4205 , n4207 );
and ( n4575 , n4204 , n4207 );
or ( n4576 , n4573 , n4574 , n4575 );
and ( n4577 , n4188 , n4192 );
and ( n4578 , n4192 , n4209 );
and ( n4579 , n4188 , n4209 );
or ( n4580 , n4577 , n4578 , n4579 );
xor ( n4581 , n4576 , n4580 );
and ( n4582 , n2206 , n607 );
not ( n4583 , n607 );
nor ( n4584 , n4582 , n4583 );
xor ( n4585 , n4581 , n4584 );
xor ( n4586 , n4572 , n4585 );
and ( n4587 , n4214 , n4226 );
and ( n4588 , n4218 , n4219 );
and ( n4589 , n4219 , n4225 );
and ( n4590 , n4218 , n4225 );
or ( n4591 , n4588 , n4589 , n4590 );
and ( n4592 , n4197 , n4202 );
and ( n4593 , n4202 , n4208 );
and ( n4594 , n4197 , n4208 );
or ( n4595 , n4592 , n4593 , n4594 );
xor ( n4596 , n4591 , n4595 );
and ( n4597 , n4198 , n4199 );
and ( n4598 , n4199 , n4201 );
and ( n4599 , n4198 , n4201 );
or ( n4600 , n4597 , n4598 , n4599 );
and ( n4601 , n1458 , n1048 );
and ( n4602 , n1713 , n905 );
xor ( n4603 , n4601 , n4602 );
and ( n4604 , n1935 , n766 );
xor ( n4605 , n4603 , n4604 );
xor ( n4606 , n4600 , n4605 );
and ( n4607 , n917 , n1685 );
and ( n4608 , n1077 , n1497 );
xor ( n4609 , n4607 , n4608 );
and ( n4610 , n1277 , n1261 );
xor ( n4611 , n4609 , n4610 );
xor ( n4612 , n4606 , n4611 );
xor ( n4613 , n4596 , n4612 );
xor ( n4614 , n4587 , n4613 );
and ( n4615 , n4221 , n4222 );
and ( n4616 , n4222 , n4224 );
and ( n4617 , n4221 , n4224 );
or ( n4618 , n4615 , n4616 , n4617 );
not ( n4619 , n521 );
and ( n4620 , n2563 , n521 );
nor ( n4621 , n4619 , n4620 );
and ( n4622 , n625 , n2271 );
xor ( n4623 , n4621 , n4622 );
and ( n4624 , n753 , n1975 );
xor ( n4625 , n4623 , n4624 );
xor ( n4626 , n4618 , n4625 );
xor ( n4627 , n4614 , n4626 );
xor ( n4628 , n4586 , n4627 );
xor ( n4629 , n4568 , n4628 );
and ( n4630 , n4160 , n4164 );
and ( n4631 , n4164 , n4229 );
and ( n4632 , n4160 , n4229 );
or ( n4633 , n4630 , n4631 , n4632 );
xor ( n4634 , n4629 , n4633 );
and ( n4635 , n4230 , n4234 );
and ( n4636 , n4235 , n4238 );
or ( n4637 , n4635 , n4636 );
xor ( n4638 , n4634 , n4637 );
buf ( n4639 , n4638 );
buf ( n4640 , n4639 );
and ( n4641 , n4640 , n279 );
xor ( n4642 , n4559 , n4641 );
xor ( n4643 , n4556 , n4642 );
xor ( n4644 , n4546 , n4643 );
xor ( n4645 , n4526 , n4644 );
xor ( n4646 , n4495 , n4645 );
xor ( n4647 , n4477 , n4646 );
and ( n4648 , n4069 , n4073 );
and ( n4649 , n4073 , n4247 );
and ( n4650 , n4069 , n4247 );
or ( n4651 , n4648 , n4649 , n4650 );
xor ( n4652 , n4647 , n4651 );
and ( n4653 , n4248 , n4252 );
and ( n4654 , n4253 , n4256 );
or ( n4655 , n4653 , n4654 );
xor ( n4656 , n4652 , n4655 );
buf ( n4657 , n4656 );
buf ( n4658 , n4657 );
not ( n4659 , n4658 );
nor ( n4660 , n4659 , n2598 );
xor ( n4661 , n4468 , n4660 );
and ( n4662 , n4065 , n4261 );
and ( n4663 , n4262 , n4265 );
or ( n4664 , n4662 , n4663 );
xor ( n4665 , n4661 , n4664 );
buf ( n4666 , n4665 );
buf ( n4667 , n4666 );
not ( n4668 , n4667 );
buf ( n4669 , n262 );
not ( n4670 , n4669 );
nor ( n4671 , n4668 , n4670 );
xor ( n4672 , n4382 , n4671 );
xor ( n4673 , n4277 , n4379 );
nor ( n4674 , n4269 , n4670 );
and ( n4675 , n4673 , n4674 );
xor ( n4676 , n4673 , n4674 );
xor ( n4677 , n4281 , n4377 );
nor ( n4678 , n3872 , n4670 );
and ( n4679 , n4677 , n4678 );
xor ( n4680 , n4677 , n4678 );
xor ( n4681 , n4285 , n4375 );
nor ( n4682 , n3473 , n4670 );
and ( n4683 , n4681 , n4682 );
xor ( n4684 , n4681 , n4682 );
xor ( n4685 , n4289 , n4373 );
nor ( n4686 , n3000 , n4670 );
and ( n4687 , n4685 , n4686 );
xor ( n4688 , n4685 , n4686 );
xor ( n4689 , n4293 , n4371 );
nor ( n4690 , n2688 , n4670 );
and ( n4691 , n4689 , n4690 );
xor ( n4692 , n4689 , n4690 );
xor ( n4693 , n4297 , n4369 );
nor ( n4694 , n3008 , n4670 );
and ( n4695 , n4693 , n4694 );
xor ( n4696 , n4693 , n4694 );
xor ( n4697 , n4301 , n4367 );
nor ( n4698 , n3017 , n4670 );
and ( n4699 , n4697 , n4698 );
xor ( n4700 , n4697 , n4698 );
xor ( n4701 , n4305 , n4365 );
nor ( n4702 , n3026 , n4670 );
and ( n4703 , n4701 , n4702 );
xor ( n4704 , n4701 , n4702 );
xor ( n4705 , n4309 , n4363 );
nor ( n4706 , n3035 , n4670 );
and ( n4707 , n4705 , n4706 );
xor ( n4708 , n4705 , n4706 );
xor ( n4709 , n4313 , n4361 );
nor ( n4710 , n3044 , n4670 );
and ( n4711 , n4709 , n4710 );
xor ( n4712 , n4709 , n4710 );
xor ( n4713 , n4317 , n4359 );
nor ( n4714 , n3053 , n4670 );
and ( n4715 , n4713 , n4714 );
xor ( n4716 , n4713 , n4714 );
xor ( n4717 , n4321 , n4357 );
nor ( n4718 , n3062 , n4670 );
and ( n4719 , n4717 , n4718 );
xor ( n4720 , n4717 , n4718 );
xor ( n4721 , n4325 , n4355 );
nor ( n4722 , n3071 , n4670 );
and ( n4723 , n4721 , n4722 );
xor ( n4724 , n4721 , n4722 );
xor ( n4725 , n4329 , n4353 );
nor ( n4726 , n3080 , n4670 );
and ( n4727 , n4725 , n4726 );
xor ( n4728 , n4725 , n4726 );
xor ( n4729 , n4333 , n4351 );
nor ( n4730 , n3089 , n4670 );
and ( n4731 , n4729 , n4730 );
xor ( n4732 , n4729 , n4730 );
xor ( n4733 , n4337 , n4349 );
nor ( n4734 , n3098 , n4670 );
and ( n4735 , n4733 , n4734 );
xor ( n4736 , n4733 , n4734 );
xor ( n4737 , n4342 , n4347 );
nor ( n4738 , n3107 , n4670 );
and ( n4739 , n4737 , n4738 );
xor ( n4740 , n4737 , n4738 );
xor ( n4741 , n4344 , n4345 );
buf ( n4742 , n4741 );
nor ( n4743 , n3116 , n4670 );
and ( n4744 , n4742 , n4743 );
xor ( n4745 , n4742 , n4743 );
nor ( n4746 , n3134 , n4271 );
buf ( n4747 , n4746 );
nor ( n4748 , n3125 , n4670 );
and ( n4749 , n4747 , n4748 );
buf ( n4750 , n4749 );
and ( n4751 , n4745 , n4750 );
or ( n4752 , n4744 , n4751 );
and ( n4753 , n4740 , n4752 );
or ( n4754 , n4739 , n4753 );
and ( n4755 , n4736 , n4754 );
or ( n4756 , n4735 , n4755 );
and ( n4757 , n4732 , n4756 );
or ( n4758 , n4731 , n4757 );
and ( n4759 , n4728 , n4758 );
or ( n4760 , n4727 , n4759 );
and ( n4761 , n4724 , n4760 );
or ( n4762 , n4723 , n4761 );
and ( n4763 , n4720 , n4762 );
or ( n4764 , n4719 , n4763 );
and ( n4765 , n4716 , n4764 );
or ( n4766 , n4715 , n4765 );
and ( n4767 , n4712 , n4766 );
or ( n4768 , n4711 , n4767 );
and ( n4769 , n4708 , n4768 );
or ( n4770 , n4707 , n4769 );
and ( n4771 , n4704 , n4770 );
or ( n4772 , n4703 , n4771 );
and ( n4773 , n4700 , n4772 );
or ( n4774 , n4699 , n4773 );
and ( n4775 , n4696 , n4774 );
or ( n4776 , n4695 , n4775 );
and ( n4777 , n4692 , n4776 );
or ( n4778 , n4691 , n4777 );
and ( n4779 , n4688 , n4778 );
or ( n4780 , n4687 , n4779 );
and ( n4781 , n4684 , n4780 );
or ( n4782 , n4683 , n4781 );
and ( n4783 , n4680 , n4782 );
or ( n4784 , n4679 , n4783 );
and ( n4785 , n4676 , n4784 );
or ( n4786 , n4675 , n4785 );
xor ( n4787 , n4672 , n4786 );
and ( n4788 , n285 , n662 );
nor ( n4789 , n663 , n4788 );
nor ( n4790 , n795 , n305 );
xor ( n4791 , n4789 , n4790 );
and ( n4792 , n4384 , n4385 );
and ( n4793 , n4386 , n4389 );
or ( n4794 , n4792 , n4793 );
xor ( n4795 , n4791 , n4794 );
nor ( n4796 , n952 , n336 );
xor ( n4797 , n4795 , n4796 );
and ( n4798 , n4390 , n4391 );
and ( n4799 , n4392 , n4395 );
or ( n4800 , n4798 , n4799 );
xor ( n4801 , n4797 , n4800 );
nor ( n4802 , n1126 , n386 );
xor ( n4803 , n4801 , n4802 );
and ( n4804 , n4396 , n4397 );
and ( n4805 , n4398 , n4401 );
or ( n4806 , n4804 , n4805 );
xor ( n4807 , n4803 , n4806 );
nor ( n4808 , n1318 , n458 );
xor ( n4809 , n4807 , n4808 );
and ( n4810 , n4402 , n4403 );
and ( n4811 , n4404 , n4407 );
or ( n4812 , n4810 , n4811 );
xor ( n4813 , n4809 , n4812 );
nor ( n4814 , n1534 , n551 );
xor ( n4815 , n4813 , n4814 );
and ( n4816 , n4408 , n4409 );
and ( n4817 , n4410 , n4413 );
or ( n4818 , n4816 , n4817 );
xor ( n4819 , n4815 , n4818 );
nor ( n4820 , n1771 , n665 );
xor ( n4821 , n4819 , n4820 );
and ( n4822 , n4414 , n4415 );
and ( n4823 , n4416 , n4419 );
or ( n4824 , n4822 , n4823 );
xor ( n4825 , n4821 , n4824 );
nor ( n4826 , n2025 , n797 );
xor ( n4827 , n4825 , n4826 );
and ( n4828 , n4420 , n4421 );
and ( n4829 , n4422 , n4425 );
or ( n4830 , n4828 , n4829 );
xor ( n4831 , n4827 , n4830 );
nor ( n4832 , n2300 , n954 );
xor ( n4833 , n4831 , n4832 );
and ( n4834 , n4426 , n4427 );
and ( n4835 , n4428 , n4431 );
or ( n4836 , n4834 , n4835 );
xor ( n4837 , n4833 , n4836 );
nor ( n4838 , n2596 , n1128 );
xor ( n4839 , n4837 , n4838 );
and ( n4840 , n4432 , n4433 );
and ( n4841 , n4434 , n4437 );
or ( n4842 , n4840 , n4841 );
xor ( n4843 , n4839 , n4842 );
nor ( n4844 , n2991 , n1320 );
xor ( n4845 , n4843 , n4844 );
and ( n4846 , n4438 , n4439 );
and ( n4847 , n4440 , n4443 );
or ( n4848 , n4846 , n4847 );
xor ( n4849 , n4845 , n4848 );
nor ( n4850 , n3464 , n1536 );
xor ( n4851 , n4849 , n4850 );
and ( n4852 , n4444 , n4445 );
and ( n4853 , n4446 , n4449 );
or ( n4854 , n4852 , n4853 );
xor ( n4855 , n4851 , n4854 );
nor ( n4856 , n3863 , n1773 );
xor ( n4857 , n4855 , n4856 );
and ( n4858 , n4450 , n4451 );
and ( n4859 , n4452 , n4455 );
or ( n4860 , n4858 , n4859 );
xor ( n4861 , n4857 , n4860 );
nor ( n4862 , n4260 , n2027 );
xor ( n4863 , n4861 , n4862 );
and ( n4864 , n4456 , n4457 );
and ( n4865 , n4458 , n4461 );
or ( n4866 , n4864 , n4865 );
xor ( n4867 , n4863 , n4866 );
nor ( n4868 , n4659 , n2302 );
xor ( n4869 , n4867 , n4868 );
and ( n4870 , n4462 , n4463 );
and ( n4871 , n4464 , n4467 );
or ( n4872 , n4870 , n4871 );
xor ( n4873 , n4869 , n4872 );
and ( n4874 , n4485 , n4489 );
and ( n4875 , n4489 , n4493 );
and ( n4876 , n4485 , n4493 );
or ( n4877 , n4874 , n4875 , n4876 );
and ( n4878 , n4481 , n4494 );
and ( n4879 , n4494 , n4645 );
and ( n4880 , n4481 , n4645 );
or ( n4881 , n4878 , n4879 , n4880 );
xor ( n4882 , n4877 , n4881 );
and ( n4883 , n4499 , n4525 );
and ( n4884 , n4525 , n4644 );
and ( n4885 , n4499 , n4644 );
or ( n4886 , n4883 , n4884 , n4885 );
and ( n4887 , n4513 , n4514 );
and ( n4888 , n4514 , n4516 );
and ( n4889 , n4513 , n4516 );
or ( n4890 , n4887 , n4888 , n4889 );
and ( n4891 , n4503 , n4507 );
and ( n4892 , n4507 , n4524 );
and ( n4893 , n4503 , n4524 );
or ( n4894 , n4891 , n4892 , n4893 );
xor ( n4895 , n4890 , n4894 );
not ( n4896 , n636 );
and ( n4897 , n2406 , n636 );
nor ( n4898 , n4896 , n4897 );
xor ( n4899 , n4895 , n4898 );
xor ( n4900 , n4886 , n4899 );
and ( n4901 , n4530 , n4545 );
and ( n4902 , n4545 , n4643 );
and ( n4903 , n4530 , n4643 );
or ( n4904 , n4901 , n4902 , n4903 );
and ( n4905 , n4512 , n4517 );
and ( n4906 , n4517 , n4523 );
and ( n4907 , n4512 , n4523 );
or ( n4908 , n4905 , n4906 , n4907 );
and ( n4909 , n4534 , n4538 );
and ( n4910 , n4538 , n4544 );
and ( n4911 , n4534 , n4544 );
or ( n4912 , n4909 , n4910 , n4911 );
xor ( n4913 , n4908 , n4912 );
and ( n4914 , n4519 , n4520 );
and ( n4915 , n4520 , n4522 );
and ( n4916 , n4519 , n4522 );
or ( n4917 , n4914 , n4915 , n4916 );
and ( n4918 , n782 , n2138 );
and ( n4919 , n931 , n1864 );
xor ( n4920 , n4918 , n4919 );
and ( n4921 , n1088 , n1753 );
xor ( n4922 , n4920 , n4921 );
xor ( n4923 , n4917 , n4922 );
and ( n4924 , n1292 , n1396 );
and ( n4925 , n1516 , n1302 );
xor ( n4926 , n4924 , n4925 );
and ( n4927 , n1730 , n1114 );
xor ( n4928 , n4926 , n4927 );
xor ( n4929 , n4923 , n4928 );
xor ( n4930 , n4913 , n4929 );
xor ( n4931 , n4904 , n4930 );
and ( n4932 , n4550 , n4555 );
and ( n4933 , n4555 , n4642 );
and ( n4934 , n4550 , n4642 );
or ( n4935 , n4932 , n4933 , n4934 );
and ( n4936 , n4540 , n4541 );
and ( n4937 , n4541 , n4543 );
and ( n4938 , n4540 , n4543 );
or ( n4939 , n4936 , n4937 , n4938 );
and ( n4940 , n4551 , n4552 );
and ( n4941 , n4552 , n4554 );
and ( n4942 , n4551 , n4554 );
or ( n4943 , n4940 , n4941 , n4942 );
xor ( n4944 , n4939 , n4943 );
and ( n4945 , n2001 , n852 );
and ( n4946 , n2286 , n714 );
xor ( n4947 , n4945 , n4946 );
and ( n4948 , n2581 , n651 );
xor ( n4949 , n4947 , n4948 );
xor ( n4950 , n4944 , n4949 );
xor ( n4951 , n4935 , n4950 );
and ( n4952 , n4557 , n4558 );
and ( n4953 , n4558 , n4641 );
and ( n4954 , n4557 , n4641 );
or ( n4955 , n4952 , n4953 , n4954 );
and ( n4956 , n2972 , n488 );
and ( n4957 , n3445 , n411 );
xor ( n4958 , n4956 , n4957 );
and ( n4959 , n3844 , n375 );
xor ( n4960 , n4958 , n4959 );
xor ( n4961 , n4955 , n4960 );
and ( n4962 , n4241 , n312 );
and ( n4963 , n4640 , n288 );
xor ( n4964 , n4962 , n4963 );
and ( n4965 , n4576 , n4580 );
and ( n4966 , n4580 , n4584 );
and ( n4967 , n4576 , n4584 );
or ( n4968 , n4965 , n4966 , n4967 );
and ( n4969 , n4572 , n4585 );
and ( n4970 , n4585 , n4627 );
and ( n4971 , n4572 , n4627 );
or ( n4972 , n4969 , n4970 , n4971 );
xor ( n4973 , n4968 , n4972 );
and ( n4974 , n4587 , n4613 );
and ( n4975 , n4613 , n4626 );
and ( n4976 , n4587 , n4626 );
or ( n4977 , n4974 , n4975 , n4976 );
and ( n4978 , n4601 , n4602 );
and ( n4979 , n4602 , n4604 );
and ( n4980 , n4601 , n4604 );
or ( n4981 , n4978 , n4979 , n4980 );
and ( n4982 , n4591 , n4595 );
and ( n4983 , n4595 , n4612 );
and ( n4984 , n4591 , n4612 );
or ( n4985 , n4982 , n4983 , n4984 );
xor ( n4986 , n4981 , n4985 );
and ( n4987 , n2206 , n766 );
not ( n4988 , n766 );
nor ( n4989 , n4987 , n4988 );
xor ( n4990 , n4986 , n4989 );
xor ( n4991 , n4977 , n4990 );
and ( n4992 , n4600 , n4605 );
and ( n4993 , n4605 , n4611 );
and ( n4994 , n4600 , n4611 );
or ( n4995 , n4992 , n4993 , n4994 );
and ( n4996 , n4618 , n4625 );
xor ( n4997 , n4995 , n4996 );
and ( n4998 , n4607 , n4608 );
and ( n4999 , n4608 , n4610 );
and ( n5000 , n4607 , n4610 );
or ( n5001 , n4998 , n4999 , n5000 );
and ( n5002 , n917 , n1975 );
and ( n5003 , n1077 , n1685 );
xor ( n5004 , n5002 , n5003 );
and ( n5005 , n1277 , n1497 );
xor ( n5006 , n5004 , n5005 );
xor ( n5007 , n5001 , n5006 );
and ( n5008 , n1458 , n1261 );
and ( n5009 , n1713 , n1048 );
xor ( n5010 , n5008 , n5009 );
and ( n5011 , n1935 , n905 );
xor ( n5012 , n5010 , n5011 );
xor ( n5013 , n5007 , n5012 );
xor ( n5014 , n4997 , n5013 );
and ( n5015 , n4621 , n4622 );
and ( n5016 , n4622 , n4624 );
and ( n5017 , n4621 , n4624 );
or ( n5018 , n5015 , n5016 , n5017 );
not ( n5019 , n625 );
and ( n5020 , n2563 , n625 );
nor ( n5021 , n5019 , n5020 );
and ( n5022 , n753 , n2271 );
xor ( n5023 , n5021 , n5022 );
xor ( n5024 , n5018 , n5023 );
xor ( n5025 , n5014 , n5024 );
xor ( n5026 , n4991 , n5025 );
xor ( n5027 , n4973 , n5026 );
and ( n5028 , n4563 , n4567 );
and ( n5029 , n4567 , n4628 );
and ( n5030 , n4563 , n4628 );
or ( n5031 , n5028 , n5029 , n5030 );
xor ( n5032 , n5027 , n5031 );
and ( n5033 , n4629 , n4633 );
and ( n5034 , n4634 , n4637 );
or ( n5035 , n5033 , n5034 );
xor ( n5036 , n5032 , n5035 );
buf ( n5037 , n5036 );
buf ( n5038 , n5037 );
and ( n5039 , n5038 , n279 );
xor ( n5040 , n4964 , n5039 );
xor ( n5041 , n4961 , n5040 );
xor ( n5042 , n4951 , n5041 );
xor ( n5043 , n4931 , n5042 );
xor ( n5044 , n4900 , n5043 );
xor ( n5045 , n4882 , n5044 );
and ( n5046 , n4472 , n4476 );
and ( n5047 , n4476 , n4646 );
and ( n5048 , n4472 , n4646 );
or ( n5049 , n5046 , n5047 , n5048 );
xor ( n5050 , n5045 , n5049 );
and ( n5051 , n4647 , n4651 );
and ( n5052 , n4652 , n4655 );
or ( n5053 , n5051 , n5052 );
xor ( n5054 , n5050 , n5053 );
buf ( n5055 , n5054 );
buf ( n5056 , n5055 );
not ( n5057 , n5056 );
nor ( n5058 , n5057 , n2598 );
xor ( n5059 , n4873 , n5058 );
and ( n5060 , n4468 , n4660 );
and ( n5061 , n4661 , n4664 );
or ( n5062 , n5060 , n5061 );
xor ( n5063 , n5059 , n5062 );
buf ( n5064 , n5063 );
buf ( n5065 , n5064 );
not ( n5066 , n5065 );
buf ( n5067 , n263 );
not ( n5068 , n5067 );
nor ( n5069 , n5066 , n5068 );
xor ( n5070 , n4787 , n5069 );
xor ( n5071 , n4676 , n4784 );
nor ( n5072 , n4668 , n5068 );
and ( n5073 , n5071 , n5072 );
xor ( n5074 , n5071 , n5072 );
xor ( n5075 , n4680 , n4782 );
nor ( n5076 , n4269 , n5068 );
and ( n5077 , n5075 , n5076 );
xor ( n5078 , n5075 , n5076 );
xor ( n5079 , n4684 , n4780 );
nor ( n5080 , n3872 , n5068 );
and ( n5081 , n5079 , n5080 );
xor ( n5082 , n5079 , n5080 );
xor ( n5083 , n4688 , n4778 );
nor ( n5084 , n3473 , n5068 );
and ( n5085 , n5083 , n5084 );
xor ( n5086 , n5083 , n5084 );
xor ( n5087 , n4692 , n4776 );
nor ( n5088 , n3000 , n5068 );
and ( n5089 , n5087 , n5088 );
xor ( n5090 , n5087 , n5088 );
xor ( n5091 , n4696 , n4774 );
nor ( n5092 , n2688 , n5068 );
and ( n5093 , n5091 , n5092 );
xor ( n5094 , n5091 , n5092 );
xor ( n5095 , n4700 , n4772 );
nor ( n5096 , n3008 , n5068 );
and ( n5097 , n5095 , n5096 );
xor ( n5098 , n5095 , n5096 );
xor ( n5099 , n4704 , n4770 );
nor ( n5100 , n3017 , n5068 );
and ( n5101 , n5099 , n5100 );
xor ( n5102 , n5099 , n5100 );
xor ( n5103 , n4708 , n4768 );
nor ( n5104 , n3026 , n5068 );
and ( n5105 , n5103 , n5104 );
xor ( n5106 , n5103 , n5104 );
xor ( n5107 , n4712 , n4766 );
nor ( n5108 , n3035 , n5068 );
and ( n5109 , n5107 , n5108 );
xor ( n5110 , n5107 , n5108 );
xor ( n5111 , n4716 , n4764 );
nor ( n5112 , n3044 , n5068 );
and ( n5113 , n5111 , n5112 );
xor ( n5114 , n5111 , n5112 );
xor ( n5115 , n4720 , n4762 );
nor ( n5116 , n3053 , n5068 );
and ( n5117 , n5115 , n5116 );
xor ( n5118 , n5115 , n5116 );
xor ( n5119 , n4724 , n4760 );
nor ( n5120 , n3062 , n5068 );
and ( n5121 , n5119 , n5120 );
xor ( n5122 , n5119 , n5120 );
xor ( n5123 , n4728 , n4758 );
nor ( n5124 , n3071 , n5068 );
and ( n5125 , n5123 , n5124 );
xor ( n5126 , n5123 , n5124 );
xor ( n5127 , n4732 , n4756 );
nor ( n5128 , n3080 , n5068 );
and ( n5129 , n5127 , n5128 );
xor ( n5130 , n5127 , n5128 );
xor ( n5131 , n4736 , n4754 );
nor ( n5132 , n3089 , n5068 );
and ( n5133 , n5131 , n5132 );
xor ( n5134 , n5131 , n5132 );
xor ( n5135 , n4740 , n4752 );
nor ( n5136 , n3098 , n5068 );
and ( n5137 , n5135 , n5136 );
xor ( n5138 , n5135 , n5136 );
xor ( n5139 , n4745 , n4750 );
nor ( n5140 , n3107 , n5068 );
and ( n5141 , n5139 , n5140 );
xor ( n5142 , n5139 , n5140 );
xor ( n5143 , n4747 , n4748 );
buf ( n5144 , n5143 );
nor ( n5145 , n3116 , n5068 );
and ( n5146 , n5144 , n5145 );
xor ( n5147 , n5144 , n5145 );
nor ( n5148 , n3134 , n4670 );
buf ( n5149 , n5148 );
nor ( n5150 , n3125 , n5068 );
and ( n5151 , n5149 , n5150 );
buf ( n5152 , n5151 );
and ( n5153 , n5147 , n5152 );
or ( n5154 , n5146 , n5153 );
and ( n5155 , n5142 , n5154 );
or ( n5156 , n5141 , n5155 );
and ( n5157 , n5138 , n5156 );
or ( n5158 , n5137 , n5157 );
and ( n5159 , n5134 , n5158 );
or ( n5160 , n5133 , n5159 );
and ( n5161 , n5130 , n5160 );
or ( n5162 , n5129 , n5161 );
and ( n5163 , n5126 , n5162 );
or ( n5164 , n5125 , n5163 );
and ( n5165 , n5122 , n5164 );
or ( n5166 , n5121 , n5165 );
and ( n5167 , n5118 , n5166 );
or ( n5168 , n5117 , n5167 );
and ( n5169 , n5114 , n5168 );
or ( n5170 , n5113 , n5169 );
and ( n5171 , n5110 , n5170 );
or ( n5172 , n5109 , n5171 );
and ( n5173 , n5106 , n5172 );
or ( n5174 , n5105 , n5173 );
and ( n5175 , n5102 , n5174 );
or ( n5176 , n5101 , n5175 );
and ( n5177 , n5098 , n5176 );
or ( n5178 , n5097 , n5177 );
and ( n5179 , n5094 , n5178 );
or ( n5180 , n5093 , n5179 );
and ( n5181 , n5090 , n5180 );
or ( n5182 , n5089 , n5181 );
and ( n5183 , n5086 , n5182 );
or ( n5184 , n5085 , n5183 );
and ( n5185 , n5082 , n5184 );
or ( n5186 , n5081 , n5185 );
and ( n5187 , n5078 , n5186 );
or ( n5188 , n5077 , n5187 );
and ( n5189 , n5074 , n5188 );
or ( n5190 , n5073 , n5189 );
xor ( n5191 , n5070 , n5190 );
and ( n5192 , n285 , n794 );
nor ( n5193 , n795 , n5192 );
nor ( n5194 , n952 , n305 );
xor ( n5195 , n5193 , n5194 );
and ( n5196 , n4789 , n4790 );
and ( n5197 , n4791 , n4794 );
or ( n5198 , n5196 , n5197 );
xor ( n5199 , n5195 , n5198 );
nor ( n5200 , n1126 , n336 );
xor ( n5201 , n5199 , n5200 );
and ( n5202 , n4795 , n4796 );
and ( n5203 , n4797 , n4800 );
or ( n5204 , n5202 , n5203 );
xor ( n5205 , n5201 , n5204 );
nor ( n5206 , n1318 , n386 );
xor ( n5207 , n5205 , n5206 );
and ( n5208 , n4801 , n4802 );
and ( n5209 , n4803 , n4806 );
or ( n5210 , n5208 , n5209 );
xor ( n5211 , n5207 , n5210 );
nor ( n5212 , n1534 , n458 );
xor ( n5213 , n5211 , n5212 );
and ( n5214 , n4807 , n4808 );
and ( n5215 , n4809 , n4812 );
or ( n5216 , n5214 , n5215 );
xor ( n5217 , n5213 , n5216 );
nor ( n5218 , n1771 , n551 );
xor ( n5219 , n5217 , n5218 );
and ( n5220 , n4813 , n4814 );
and ( n5221 , n4815 , n4818 );
or ( n5222 , n5220 , n5221 );
xor ( n5223 , n5219 , n5222 );
nor ( n5224 , n2025 , n665 );
xor ( n5225 , n5223 , n5224 );
and ( n5226 , n4819 , n4820 );
and ( n5227 , n4821 , n4824 );
or ( n5228 , n5226 , n5227 );
xor ( n5229 , n5225 , n5228 );
nor ( n5230 , n2300 , n797 );
xor ( n5231 , n5229 , n5230 );
and ( n5232 , n4825 , n4826 );
and ( n5233 , n4827 , n4830 );
or ( n5234 , n5232 , n5233 );
xor ( n5235 , n5231 , n5234 );
nor ( n5236 , n2596 , n954 );
xor ( n5237 , n5235 , n5236 );
and ( n5238 , n4831 , n4832 );
and ( n5239 , n4833 , n4836 );
or ( n5240 , n5238 , n5239 );
xor ( n5241 , n5237 , n5240 );
nor ( n5242 , n2991 , n1128 );
xor ( n5243 , n5241 , n5242 );
and ( n5244 , n4837 , n4838 );
and ( n5245 , n4839 , n4842 );
or ( n5246 , n5244 , n5245 );
xor ( n5247 , n5243 , n5246 );
nor ( n5248 , n3464 , n1320 );
xor ( n5249 , n5247 , n5248 );
and ( n5250 , n4843 , n4844 );
and ( n5251 , n4845 , n4848 );
or ( n5252 , n5250 , n5251 );
xor ( n5253 , n5249 , n5252 );
nor ( n5254 , n3863 , n1536 );
xor ( n5255 , n5253 , n5254 );
and ( n5256 , n4849 , n4850 );
and ( n5257 , n4851 , n4854 );
or ( n5258 , n5256 , n5257 );
xor ( n5259 , n5255 , n5258 );
nor ( n5260 , n4260 , n1773 );
xor ( n5261 , n5259 , n5260 );
and ( n5262 , n4855 , n4856 );
and ( n5263 , n4857 , n4860 );
or ( n5264 , n5262 , n5263 );
xor ( n5265 , n5261 , n5264 );
nor ( n5266 , n4659 , n2027 );
xor ( n5267 , n5265 , n5266 );
and ( n5268 , n4861 , n4862 );
and ( n5269 , n4863 , n4866 );
or ( n5270 , n5268 , n5269 );
xor ( n5271 , n5267 , n5270 );
nor ( n5272 , n5057 , n2302 );
xor ( n5273 , n5271 , n5272 );
and ( n5274 , n4867 , n4868 );
and ( n5275 , n4869 , n4872 );
or ( n5276 , n5274 , n5275 );
xor ( n5277 , n5273 , n5276 );
and ( n5278 , n4890 , n4894 );
and ( n5279 , n4894 , n4898 );
and ( n5280 , n4890 , n4898 );
or ( n5281 , n5278 , n5279 , n5280 );
and ( n5282 , n4886 , n4899 );
and ( n5283 , n4899 , n5043 );
and ( n5284 , n4886 , n5043 );
or ( n5285 , n5282 , n5283 , n5284 );
xor ( n5286 , n5281 , n5285 );
and ( n5287 , n4904 , n4930 );
and ( n5288 , n4930 , n5042 );
and ( n5289 , n4904 , n5042 );
or ( n5290 , n5287 , n5288 , n5289 );
and ( n5291 , n4918 , n4919 );
and ( n5292 , n4919 , n4921 );
and ( n5293 , n4918 , n4921 );
or ( n5294 , n5291 , n5292 , n5293 );
and ( n5295 , n4908 , n4912 );
and ( n5296 , n4912 , n4929 );
and ( n5297 , n4908 , n4929 );
or ( n5298 , n5295 , n5296 , n5297 );
xor ( n5299 , n5294 , n5298 );
not ( n5300 , n782 );
and ( n5301 , n2406 , n782 );
nor ( n5302 , n5300 , n5301 );
xor ( n5303 , n5299 , n5302 );
xor ( n5304 , n5290 , n5303 );
and ( n5305 , n4935 , n4950 );
and ( n5306 , n4950 , n5041 );
and ( n5307 , n4935 , n5041 );
or ( n5308 , n5305 , n5306 , n5307 );
and ( n5309 , n4917 , n4922 );
and ( n5310 , n4922 , n4928 );
and ( n5311 , n4917 , n4928 );
or ( n5312 , n5309 , n5310 , n5311 );
and ( n5313 , n4939 , n4943 );
and ( n5314 , n4943 , n4949 );
and ( n5315 , n4939 , n4949 );
or ( n5316 , n5313 , n5314 , n5315 );
xor ( n5317 , n5312 , n5316 );
and ( n5318 , n4924 , n4925 );
and ( n5319 , n4925 , n4927 );
and ( n5320 , n4924 , n4927 );
or ( n5321 , n5318 , n5319 , n5320 );
and ( n5322 , n931 , n2138 );
and ( n5323 , n1088 , n1864 );
xor ( n5324 , n5322 , n5323 );
and ( n5325 , n1292 , n1753 );
xor ( n5326 , n5324 , n5325 );
xor ( n5327 , n5321 , n5326 );
and ( n5328 , n1516 , n1396 );
and ( n5329 , n1730 , n1302 );
xor ( n5330 , n5328 , n5329 );
and ( n5331 , n2001 , n1114 );
xor ( n5332 , n5330 , n5331 );
xor ( n5333 , n5327 , n5332 );
xor ( n5334 , n5317 , n5333 );
xor ( n5335 , n5308 , n5334 );
and ( n5336 , n4955 , n4960 );
and ( n5337 , n4960 , n5040 );
and ( n5338 , n4955 , n5040 );
or ( n5339 , n5336 , n5337 , n5338 );
and ( n5340 , n4945 , n4946 );
and ( n5341 , n4946 , n4948 );
and ( n5342 , n4945 , n4948 );
or ( n5343 , n5340 , n5341 , n5342 );
and ( n5344 , n4956 , n4957 );
and ( n5345 , n4957 , n4959 );
and ( n5346 , n4956 , n4959 );
or ( n5347 , n5344 , n5345 , n5346 );
xor ( n5348 , n5343 , n5347 );
and ( n5349 , n2286 , n852 );
and ( n5350 , n2581 , n714 );
xor ( n5351 , n5349 , n5350 );
and ( n5352 , n2972 , n651 );
xor ( n5353 , n5351 , n5352 );
xor ( n5354 , n5348 , n5353 );
xor ( n5355 , n5339 , n5354 );
and ( n5356 , n4962 , n4963 );
and ( n5357 , n4963 , n5039 );
and ( n5358 , n4962 , n5039 );
or ( n5359 , n5356 , n5357 , n5358 );
and ( n5360 , n3445 , n488 );
and ( n5361 , n3844 , n411 );
xor ( n5362 , n5360 , n5361 );
and ( n5363 , n4241 , n375 );
xor ( n5364 , n5362 , n5363 );
xor ( n5365 , n5359 , n5364 );
and ( n5366 , n4640 , n312 );
and ( n5367 , n5038 , n288 );
xor ( n5368 , n5366 , n5367 );
and ( n5369 , n4981 , n4985 );
and ( n5370 , n4985 , n4989 );
and ( n5371 , n4981 , n4989 );
or ( n5372 , n5369 , n5370 , n5371 );
and ( n5373 , n4977 , n4990 );
and ( n5374 , n4990 , n5025 );
and ( n5375 , n4977 , n5025 );
or ( n5376 , n5373 , n5374 , n5375 );
xor ( n5377 , n5372 , n5376 );
and ( n5378 , n5014 , n5024 );
and ( n5379 , n5008 , n5009 );
and ( n5380 , n5009 , n5011 );
and ( n5381 , n5008 , n5011 );
or ( n5382 , n5379 , n5380 , n5381 );
and ( n5383 , n4995 , n4996 );
and ( n5384 , n4996 , n5013 );
and ( n5385 , n4995 , n5013 );
or ( n5386 , n5383 , n5384 , n5385 );
xor ( n5387 , n5382 , n5386 );
and ( n5388 , n2206 , n905 );
not ( n5389 , n905 );
nor ( n5390 , n5388 , n5389 );
xor ( n5391 , n5387 , n5390 );
xor ( n5392 , n5378 , n5391 );
and ( n5393 , n5001 , n5006 );
and ( n5394 , n5006 , n5012 );
and ( n5395 , n5001 , n5012 );
or ( n5396 , n5393 , n5394 , n5395 );
and ( n5397 , n5018 , n5023 );
xor ( n5398 , n5396 , n5397 );
and ( n5399 , n5002 , n5003 );
and ( n5400 , n5003 , n5005 );
and ( n5401 , n5002 , n5005 );
or ( n5402 , n5399 , n5400 , n5401 );
and ( n5403 , n1458 , n1497 );
and ( n5404 , n1713 , n1261 );
xor ( n5405 , n5403 , n5404 );
and ( n5406 , n1935 , n1048 );
xor ( n5407 , n5405 , n5406 );
xor ( n5408 , n5402 , n5407 );
and ( n5409 , n917 , n2271 );
and ( n5410 , n1077 , n1975 );
xor ( n5411 , n5409 , n5410 );
and ( n5412 , n1277 , n1685 );
xor ( n5413 , n5411 , n5412 );
xor ( n5414 , n5408 , n5413 );
xor ( n5415 , n5398 , n5414 );
and ( n5416 , n5021 , n5022 );
not ( n5417 , n753 );
and ( n5418 , n2563 , n753 );
nor ( n5419 , n5417 , n5418 );
xor ( n5420 , n5416 , n5419 );
xor ( n5421 , n5415 , n5420 );
xor ( n5422 , n5392 , n5421 );
xor ( n5423 , n5377 , n5422 );
and ( n5424 , n4968 , n4972 );
and ( n5425 , n4972 , n5026 );
and ( n5426 , n4968 , n5026 );
or ( n5427 , n5424 , n5425 , n5426 );
xor ( n5428 , n5423 , n5427 );
and ( n5429 , n5027 , n5031 );
and ( n5430 , n5032 , n5035 );
or ( n5431 , n5429 , n5430 );
xor ( n5432 , n5428 , n5431 );
buf ( n5433 , n5432 );
buf ( n5434 , n5433 );
and ( n5435 , n5434 , n279 );
xor ( n5436 , n5368 , n5435 );
xor ( n5437 , n5365 , n5436 );
xor ( n5438 , n5355 , n5437 );
xor ( n5439 , n5335 , n5438 );
xor ( n5440 , n5304 , n5439 );
xor ( n5441 , n5286 , n5440 );
and ( n5442 , n4877 , n4881 );
and ( n5443 , n4881 , n5044 );
and ( n5444 , n4877 , n5044 );
or ( n5445 , n5442 , n5443 , n5444 );
xor ( n5446 , n5441 , n5445 );
and ( n5447 , n5045 , n5049 );
and ( n5448 , n5050 , n5053 );
or ( n5449 , n5447 , n5448 );
xor ( n5450 , n5446 , n5449 );
buf ( n5451 , n5450 );
buf ( n5452 , n5451 );
not ( n5453 , n5452 );
nor ( n5454 , n5453 , n2598 );
xor ( n5455 , n5277 , n5454 );
and ( n5456 , n4873 , n5058 );
and ( n5457 , n5059 , n5062 );
or ( n5458 , n5456 , n5457 );
xor ( n5459 , n5455 , n5458 );
buf ( n5460 , n5459 );
buf ( n5461 , n5460 );
not ( n5462 , n5461 );
buf ( n5463 , n264 );
not ( n5464 , n5463 );
nor ( n5465 , n5462 , n5464 );
xor ( n5466 , n5191 , n5465 );
xor ( n5467 , n5074 , n5188 );
nor ( n5468 , n5066 , n5464 );
and ( n5469 , n5467 , n5468 );
xor ( n5470 , n5467 , n5468 );
xor ( n5471 , n5078 , n5186 );
nor ( n5472 , n4668 , n5464 );
and ( n5473 , n5471 , n5472 );
xor ( n5474 , n5471 , n5472 );
xor ( n5475 , n5082 , n5184 );
nor ( n5476 , n4269 , n5464 );
and ( n5477 , n5475 , n5476 );
xor ( n5478 , n5475 , n5476 );
xor ( n5479 , n5086 , n5182 );
nor ( n5480 , n3872 , n5464 );
and ( n5481 , n5479 , n5480 );
xor ( n5482 , n5479 , n5480 );
xor ( n5483 , n5090 , n5180 );
nor ( n5484 , n3473 , n5464 );
and ( n5485 , n5483 , n5484 );
xor ( n5486 , n5483 , n5484 );
xor ( n5487 , n5094 , n5178 );
nor ( n5488 , n3000 , n5464 );
and ( n5489 , n5487 , n5488 );
xor ( n5490 , n5487 , n5488 );
xor ( n5491 , n5098 , n5176 );
nor ( n5492 , n2688 , n5464 );
and ( n5493 , n5491 , n5492 );
xor ( n5494 , n5491 , n5492 );
xor ( n5495 , n5102 , n5174 );
nor ( n5496 , n3008 , n5464 );
and ( n5497 , n5495 , n5496 );
xor ( n5498 , n5495 , n5496 );
xor ( n5499 , n5106 , n5172 );
nor ( n5500 , n3017 , n5464 );
and ( n5501 , n5499 , n5500 );
xor ( n5502 , n5499 , n5500 );
xor ( n5503 , n5110 , n5170 );
nor ( n5504 , n3026 , n5464 );
and ( n5505 , n5503 , n5504 );
xor ( n5506 , n5503 , n5504 );
xor ( n5507 , n5114 , n5168 );
nor ( n5508 , n3035 , n5464 );
and ( n5509 , n5507 , n5508 );
xor ( n5510 , n5507 , n5508 );
xor ( n5511 , n5118 , n5166 );
nor ( n5512 , n3044 , n5464 );
and ( n5513 , n5511 , n5512 );
xor ( n5514 , n5511 , n5512 );
xor ( n5515 , n5122 , n5164 );
nor ( n5516 , n3053 , n5464 );
and ( n5517 , n5515 , n5516 );
xor ( n5518 , n5515 , n5516 );
xor ( n5519 , n5126 , n5162 );
nor ( n5520 , n3062 , n5464 );
and ( n5521 , n5519 , n5520 );
xor ( n5522 , n5519 , n5520 );
xor ( n5523 , n5130 , n5160 );
nor ( n5524 , n3071 , n5464 );
and ( n5525 , n5523 , n5524 );
xor ( n5526 , n5523 , n5524 );
xor ( n5527 , n5134 , n5158 );
nor ( n5528 , n3080 , n5464 );
and ( n5529 , n5527 , n5528 );
xor ( n5530 , n5527 , n5528 );
xor ( n5531 , n5138 , n5156 );
nor ( n5532 , n3089 , n5464 );
and ( n5533 , n5531 , n5532 );
xor ( n5534 , n5531 , n5532 );
xor ( n5535 , n5142 , n5154 );
nor ( n5536 , n3098 , n5464 );
and ( n5537 , n5535 , n5536 );
xor ( n5538 , n5535 , n5536 );
xor ( n5539 , n5147 , n5152 );
nor ( n5540 , n3107 , n5464 );
and ( n5541 , n5539 , n5540 );
xor ( n5542 , n5539 , n5540 );
xor ( n5543 , n5149 , n5150 );
buf ( n5544 , n5543 );
nor ( n5545 , n3116 , n5464 );
and ( n5546 , n5544 , n5545 );
xor ( n5547 , n5544 , n5545 );
nor ( n5548 , n3134 , n5068 );
buf ( n5549 , n5548 );
nor ( n5550 , n3125 , n5464 );
and ( n5551 , n5549 , n5550 );
buf ( n5552 , n5551 );
and ( n5553 , n5547 , n5552 );
or ( n5554 , n5546 , n5553 );
and ( n5555 , n5542 , n5554 );
or ( n5556 , n5541 , n5555 );
and ( n5557 , n5538 , n5556 );
or ( n5558 , n5537 , n5557 );
and ( n5559 , n5534 , n5558 );
or ( n5560 , n5533 , n5559 );
and ( n5561 , n5530 , n5560 );
or ( n5562 , n5529 , n5561 );
and ( n5563 , n5526 , n5562 );
or ( n5564 , n5525 , n5563 );
and ( n5565 , n5522 , n5564 );
or ( n5566 , n5521 , n5565 );
and ( n5567 , n5518 , n5566 );
or ( n5568 , n5517 , n5567 );
and ( n5569 , n5514 , n5568 );
or ( n5570 , n5513 , n5569 );
and ( n5571 , n5510 , n5570 );
or ( n5572 , n5509 , n5571 );
and ( n5573 , n5506 , n5572 );
or ( n5574 , n5505 , n5573 );
and ( n5575 , n5502 , n5574 );
or ( n5576 , n5501 , n5575 );
and ( n5577 , n5498 , n5576 );
or ( n5578 , n5497 , n5577 );
and ( n5579 , n5494 , n5578 );
or ( n5580 , n5493 , n5579 );
and ( n5581 , n5490 , n5580 );
or ( n5582 , n5489 , n5581 );
and ( n5583 , n5486 , n5582 );
or ( n5584 , n5485 , n5583 );
and ( n5585 , n5482 , n5584 );
or ( n5586 , n5481 , n5585 );
and ( n5587 , n5478 , n5586 );
or ( n5588 , n5477 , n5587 );
and ( n5589 , n5474 , n5588 );
or ( n5590 , n5473 , n5589 );
and ( n5591 , n5470 , n5590 );
or ( n5592 , n5469 , n5591 );
xor ( n5593 , n5466 , n5592 );
and ( n5594 , n285 , n951 );
nor ( n5595 , n952 , n5594 );
nor ( n5596 , n1126 , n305 );
xor ( n5597 , n5595 , n5596 );
and ( n5598 , n5193 , n5194 );
and ( n5599 , n5195 , n5198 );
or ( n5600 , n5598 , n5599 );
xor ( n5601 , n5597 , n5600 );
nor ( n5602 , n1318 , n336 );
xor ( n5603 , n5601 , n5602 );
and ( n5604 , n5199 , n5200 );
and ( n5605 , n5201 , n5204 );
or ( n5606 , n5604 , n5605 );
xor ( n5607 , n5603 , n5606 );
nor ( n5608 , n1534 , n386 );
xor ( n5609 , n5607 , n5608 );
and ( n5610 , n5205 , n5206 );
and ( n5611 , n5207 , n5210 );
or ( n5612 , n5610 , n5611 );
xor ( n5613 , n5609 , n5612 );
nor ( n5614 , n1771 , n458 );
xor ( n5615 , n5613 , n5614 );
and ( n5616 , n5211 , n5212 );
and ( n5617 , n5213 , n5216 );
or ( n5618 , n5616 , n5617 );
xor ( n5619 , n5615 , n5618 );
nor ( n5620 , n2025 , n551 );
xor ( n5621 , n5619 , n5620 );
and ( n5622 , n5217 , n5218 );
and ( n5623 , n5219 , n5222 );
or ( n5624 , n5622 , n5623 );
xor ( n5625 , n5621 , n5624 );
nor ( n5626 , n2300 , n665 );
xor ( n5627 , n5625 , n5626 );
and ( n5628 , n5223 , n5224 );
and ( n5629 , n5225 , n5228 );
or ( n5630 , n5628 , n5629 );
xor ( n5631 , n5627 , n5630 );
nor ( n5632 , n2596 , n797 );
xor ( n5633 , n5631 , n5632 );
and ( n5634 , n5229 , n5230 );
and ( n5635 , n5231 , n5234 );
or ( n5636 , n5634 , n5635 );
xor ( n5637 , n5633 , n5636 );
nor ( n5638 , n2991 , n954 );
xor ( n5639 , n5637 , n5638 );
and ( n5640 , n5235 , n5236 );
and ( n5641 , n5237 , n5240 );
or ( n5642 , n5640 , n5641 );
xor ( n5643 , n5639 , n5642 );
nor ( n5644 , n3464 , n1128 );
xor ( n5645 , n5643 , n5644 );
and ( n5646 , n5241 , n5242 );
and ( n5647 , n5243 , n5246 );
or ( n5648 , n5646 , n5647 );
xor ( n5649 , n5645 , n5648 );
nor ( n5650 , n3863 , n1320 );
xor ( n5651 , n5649 , n5650 );
and ( n5652 , n5247 , n5248 );
and ( n5653 , n5249 , n5252 );
or ( n5654 , n5652 , n5653 );
xor ( n5655 , n5651 , n5654 );
nor ( n5656 , n4260 , n1536 );
xor ( n5657 , n5655 , n5656 );
and ( n5658 , n5253 , n5254 );
and ( n5659 , n5255 , n5258 );
or ( n5660 , n5658 , n5659 );
xor ( n5661 , n5657 , n5660 );
nor ( n5662 , n4659 , n1773 );
xor ( n5663 , n5661 , n5662 );
and ( n5664 , n5259 , n5260 );
and ( n5665 , n5261 , n5264 );
or ( n5666 , n5664 , n5665 );
xor ( n5667 , n5663 , n5666 );
nor ( n5668 , n5057 , n2027 );
xor ( n5669 , n5667 , n5668 );
and ( n5670 , n5265 , n5266 );
and ( n5671 , n5267 , n5270 );
or ( n5672 , n5670 , n5671 );
xor ( n5673 , n5669 , n5672 );
nor ( n5674 , n5453 , n2302 );
xor ( n5675 , n5673 , n5674 );
and ( n5676 , n5271 , n5272 );
and ( n5677 , n5273 , n5276 );
or ( n5678 , n5676 , n5677 );
xor ( n5679 , n5675 , n5678 );
and ( n5680 , n5294 , n5298 );
and ( n5681 , n5298 , n5302 );
and ( n5682 , n5294 , n5302 );
or ( n5683 , n5680 , n5681 , n5682 );
and ( n5684 , n5290 , n5303 );
and ( n5685 , n5303 , n5439 );
and ( n5686 , n5290 , n5439 );
or ( n5687 , n5684 , n5685 , n5686 );
xor ( n5688 , n5683 , n5687 );
and ( n5689 , n5308 , n5334 );
and ( n5690 , n5334 , n5438 );
and ( n5691 , n5308 , n5438 );
or ( n5692 , n5689 , n5690 , n5691 );
and ( n5693 , n5322 , n5323 );
and ( n5694 , n5323 , n5325 );
and ( n5695 , n5322 , n5325 );
or ( n5696 , n5693 , n5694 , n5695 );
and ( n5697 , n5312 , n5316 );
and ( n5698 , n5316 , n5333 );
and ( n5699 , n5312 , n5333 );
or ( n5700 , n5697 , n5698 , n5699 );
xor ( n5701 , n5696 , n5700 );
not ( n5702 , n931 );
and ( n5703 , n2406 , n931 );
nor ( n5704 , n5702 , n5703 );
xor ( n5705 , n5701 , n5704 );
xor ( n5706 , n5692 , n5705 );
and ( n5707 , n5339 , n5354 );
and ( n5708 , n5354 , n5437 );
and ( n5709 , n5339 , n5437 );
or ( n5710 , n5707 , n5708 , n5709 );
and ( n5711 , n5321 , n5326 );
and ( n5712 , n5326 , n5332 );
and ( n5713 , n5321 , n5332 );
or ( n5714 , n5711 , n5712 , n5713 );
and ( n5715 , n5343 , n5347 );
and ( n5716 , n5347 , n5353 );
and ( n5717 , n5343 , n5353 );
or ( n5718 , n5715 , n5716 , n5717 );
xor ( n5719 , n5714 , n5718 );
and ( n5720 , n5328 , n5329 );
and ( n5721 , n5329 , n5331 );
and ( n5722 , n5328 , n5331 );
or ( n5723 , n5720 , n5721 , n5722 );
and ( n5724 , n1088 , n2138 );
and ( n5725 , n1292 , n1864 );
xor ( n5726 , n5724 , n5725 );
and ( n5727 , n1516 , n1753 );
xor ( n5728 , n5726 , n5727 );
xor ( n5729 , n5723 , n5728 );
and ( n5730 , n1730 , n1396 );
and ( n5731 , n2001 , n1302 );
xor ( n5732 , n5730 , n5731 );
and ( n5733 , n2286 , n1114 );
xor ( n5734 , n5732 , n5733 );
xor ( n5735 , n5729 , n5734 );
xor ( n5736 , n5719 , n5735 );
xor ( n5737 , n5710 , n5736 );
and ( n5738 , n5359 , n5364 );
and ( n5739 , n5364 , n5436 );
and ( n5740 , n5359 , n5436 );
or ( n5741 , n5738 , n5739 , n5740 );
and ( n5742 , n5349 , n5350 );
and ( n5743 , n5350 , n5352 );
and ( n5744 , n5349 , n5352 );
or ( n5745 , n5742 , n5743 , n5744 );
and ( n5746 , n5360 , n5361 );
and ( n5747 , n5361 , n5363 );
and ( n5748 , n5360 , n5363 );
or ( n5749 , n5746 , n5747 , n5748 );
xor ( n5750 , n5745 , n5749 );
and ( n5751 , n2581 , n852 );
and ( n5752 , n2972 , n714 );
xor ( n5753 , n5751 , n5752 );
and ( n5754 , n3445 , n651 );
xor ( n5755 , n5753 , n5754 );
xor ( n5756 , n5750 , n5755 );
xor ( n5757 , n5741 , n5756 );
and ( n5758 , n5366 , n5367 );
and ( n5759 , n5367 , n5435 );
and ( n5760 , n5366 , n5435 );
or ( n5761 , n5758 , n5759 , n5760 );
and ( n5762 , n3844 , n488 );
and ( n5763 , n4241 , n411 );
xor ( n5764 , n5762 , n5763 );
and ( n5765 , n4640 , n375 );
xor ( n5766 , n5764 , n5765 );
xor ( n5767 , n5761 , n5766 );
and ( n5768 , n5038 , n312 );
and ( n5769 , n5434 , n288 );
xor ( n5770 , n5768 , n5769 );
and ( n5771 , n5382 , n5386 );
and ( n5772 , n5386 , n5390 );
and ( n5773 , n5382 , n5390 );
or ( n5774 , n5771 , n5772 , n5773 );
and ( n5775 , n5378 , n5391 );
and ( n5776 , n5391 , n5421 );
and ( n5777 , n5378 , n5421 );
or ( n5778 , n5775 , n5776 , n5777 );
xor ( n5779 , n5774 , n5778 );
and ( n5780 , n5415 , n5420 );
and ( n5781 , n5403 , n5404 );
and ( n5782 , n5404 , n5406 );
and ( n5783 , n5403 , n5406 );
or ( n5784 , n5781 , n5782 , n5783 );
and ( n5785 , n5396 , n5397 );
and ( n5786 , n5397 , n5414 );
and ( n5787 , n5396 , n5414 );
or ( n5788 , n5785 , n5786 , n5787 );
xor ( n5789 , n5784 , n5788 );
and ( n5790 , n2206 , n1048 );
not ( n5791 , n1048 );
nor ( n5792 , n5790 , n5791 );
xor ( n5793 , n5789 , n5792 );
xor ( n5794 , n5780 , n5793 );
and ( n5795 , n5402 , n5407 );
and ( n5796 , n5407 , n5413 );
and ( n5797 , n5402 , n5413 );
or ( n5798 , n5795 , n5796 , n5797 );
and ( n5799 , n5416 , n5419 );
xor ( n5800 , n5798 , n5799 );
and ( n5801 , n5409 , n5410 );
and ( n5802 , n5410 , n5412 );
and ( n5803 , n5409 , n5412 );
or ( n5804 , n5801 , n5802 , n5803 );
and ( n5805 , n1458 , n1685 );
and ( n5806 , n1713 , n1497 );
xor ( n5807 , n5805 , n5806 );
and ( n5808 , n1935 , n1261 );
xor ( n5809 , n5807 , n5808 );
xor ( n5810 , n5804 , n5809 );
not ( n5811 , n917 );
and ( n5812 , n2563 , n917 );
nor ( n5813 , n5811 , n5812 );
and ( n5814 , n1077 , n2271 );
xor ( n5815 , n5813 , n5814 );
and ( n5816 , n1277 , n1975 );
xor ( n5817 , n5815 , n5816 );
xor ( n5818 , n5810 , n5817 );
xor ( n5819 , n5800 , n5818 );
xor ( n5820 , n5794 , n5819 );
xor ( n5821 , n5779 , n5820 );
and ( n5822 , n5372 , n5376 );
and ( n5823 , n5376 , n5422 );
and ( n5824 , n5372 , n5422 );
or ( n5825 , n5822 , n5823 , n5824 );
xor ( n5826 , n5821 , n5825 );
and ( n5827 , n5423 , n5427 );
and ( n5828 , n5428 , n5431 );
or ( n5829 , n5827 , n5828 );
xor ( n5830 , n5826 , n5829 );
buf ( n5831 , n5830 );
buf ( n5832 , n5831 );
and ( n5833 , n5832 , n279 );
xor ( n5834 , n5770 , n5833 );
xor ( n5835 , n5767 , n5834 );
xor ( n5836 , n5757 , n5835 );
xor ( n5837 , n5737 , n5836 );
xor ( n5838 , n5706 , n5837 );
xor ( n5839 , n5688 , n5838 );
and ( n5840 , n5281 , n5285 );
and ( n5841 , n5285 , n5440 );
and ( n5842 , n5281 , n5440 );
or ( n5843 , n5840 , n5841 , n5842 );
xor ( n5844 , n5839 , n5843 );
and ( n5845 , n5441 , n5445 );
and ( n5846 , n5446 , n5449 );
or ( n5847 , n5845 , n5846 );
xor ( n5848 , n5844 , n5847 );
buf ( n5849 , n5848 );
buf ( n5850 , n5849 );
not ( n5851 , n5850 );
nor ( n5852 , n5851 , n2598 );
xor ( n5853 , n5679 , n5852 );
and ( n5854 , n5277 , n5454 );
and ( n5855 , n5455 , n5458 );
or ( n5856 , n5854 , n5855 );
xor ( n5857 , n5853 , n5856 );
buf ( n5858 , n5857 );
buf ( n5859 , n5858 );
not ( n5860 , n5859 );
buf ( n5861 , n265 );
not ( n5862 , n5861 );
nor ( n5863 , n5860 , n5862 );
xor ( n5864 , n5593 , n5863 );
xor ( n5865 , n5470 , n5590 );
nor ( n5866 , n5462 , n5862 );
and ( n5867 , n5865 , n5866 );
xor ( n5868 , n5865 , n5866 );
xor ( n5869 , n5474 , n5588 );
nor ( n5870 , n5066 , n5862 );
and ( n5871 , n5869 , n5870 );
xor ( n5872 , n5869 , n5870 );
xor ( n5873 , n5478 , n5586 );
nor ( n5874 , n4668 , n5862 );
and ( n5875 , n5873 , n5874 );
xor ( n5876 , n5873 , n5874 );
xor ( n5877 , n5482 , n5584 );
nor ( n5878 , n4269 , n5862 );
and ( n5879 , n5877 , n5878 );
xor ( n5880 , n5877 , n5878 );
xor ( n5881 , n5486 , n5582 );
nor ( n5882 , n3872 , n5862 );
and ( n5883 , n5881 , n5882 );
xor ( n5884 , n5881 , n5882 );
xor ( n5885 , n5490 , n5580 );
nor ( n5886 , n3473 , n5862 );
and ( n5887 , n5885 , n5886 );
xor ( n5888 , n5885 , n5886 );
xor ( n5889 , n5494 , n5578 );
nor ( n5890 , n3000 , n5862 );
and ( n5891 , n5889 , n5890 );
xor ( n5892 , n5889 , n5890 );
xor ( n5893 , n5498 , n5576 );
nor ( n5894 , n2688 , n5862 );
and ( n5895 , n5893 , n5894 );
xor ( n5896 , n5893 , n5894 );
xor ( n5897 , n5502 , n5574 );
nor ( n5898 , n3008 , n5862 );
and ( n5899 , n5897 , n5898 );
xor ( n5900 , n5897 , n5898 );
xor ( n5901 , n5506 , n5572 );
nor ( n5902 , n3017 , n5862 );
and ( n5903 , n5901 , n5902 );
xor ( n5904 , n5901 , n5902 );
xor ( n5905 , n5510 , n5570 );
nor ( n5906 , n3026 , n5862 );
and ( n5907 , n5905 , n5906 );
xor ( n5908 , n5905 , n5906 );
xor ( n5909 , n5514 , n5568 );
nor ( n5910 , n3035 , n5862 );
and ( n5911 , n5909 , n5910 );
xor ( n5912 , n5909 , n5910 );
xor ( n5913 , n5518 , n5566 );
nor ( n5914 , n3044 , n5862 );
and ( n5915 , n5913 , n5914 );
xor ( n5916 , n5913 , n5914 );
xor ( n5917 , n5522 , n5564 );
nor ( n5918 , n3053 , n5862 );
and ( n5919 , n5917 , n5918 );
xor ( n5920 , n5917 , n5918 );
xor ( n5921 , n5526 , n5562 );
nor ( n5922 , n3062 , n5862 );
and ( n5923 , n5921 , n5922 );
xor ( n5924 , n5921 , n5922 );
xor ( n5925 , n5530 , n5560 );
nor ( n5926 , n3071 , n5862 );
and ( n5927 , n5925 , n5926 );
xor ( n5928 , n5925 , n5926 );
xor ( n5929 , n5534 , n5558 );
nor ( n5930 , n3080 , n5862 );
and ( n5931 , n5929 , n5930 );
xor ( n5932 , n5929 , n5930 );
xor ( n5933 , n5538 , n5556 );
nor ( n5934 , n3089 , n5862 );
and ( n5935 , n5933 , n5934 );
xor ( n5936 , n5933 , n5934 );
xor ( n5937 , n5542 , n5554 );
nor ( n5938 , n3098 , n5862 );
and ( n5939 , n5937 , n5938 );
xor ( n5940 , n5937 , n5938 );
xor ( n5941 , n5547 , n5552 );
nor ( n5942 , n3107 , n5862 );
and ( n5943 , n5941 , n5942 );
xor ( n5944 , n5941 , n5942 );
xor ( n5945 , n5549 , n5550 );
buf ( n5946 , n5945 );
nor ( n5947 , n3116 , n5862 );
and ( n5948 , n5946 , n5947 );
xor ( n5949 , n5946 , n5947 );
nor ( n5950 , n3134 , n5464 );
buf ( n5951 , n5950 );
nor ( n5952 , n3125 , n5862 );
and ( n5953 , n5951 , n5952 );
buf ( n5954 , n5953 );
and ( n5955 , n5949 , n5954 );
or ( n5956 , n5948 , n5955 );
and ( n5957 , n5944 , n5956 );
or ( n5958 , n5943 , n5957 );
and ( n5959 , n5940 , n5958 );
or ( n5960 , n5939 , n5959 );
and ( n5961 , n5936 , n5960 );
or ( n5962 , n5935 , n5961 );
and ( n5963 , n5932 , n5962 );
or ( n5964 , n5931 , n5963 );
and ( n5965 , n5928 , n5964 );
or ( n5966 , n5927 , n5965 );
and ( n5967 , n5924 , n5966 );
or ( n5968 , n5923 , n5967 );
and ( n5969 , n5920 , n5968 );
or ( n5970 , n5919 , n5969 );
and ( n5971 , n5916 , n5970 );
or ( n5972 , n5915 , n5971 );
and ( n5973 , n5912 , n5972 );
or ( n5974 , n5911 , n5973 );
and ( n5975 , n5908 , n5974 );
or ( n5976 , n5907 , n5975 );
and ( n5977 , n5904 , n5976 );
or ( n5978 , n5903 , n5977 );
and ( n5979 , n5900 , n5978 );
or ( n5980 , n5899 , n5979 );
and ( n5981 , n5896 , n5980 );
or ( n5982 , n5895 , n5981 );
and ( n5983 , n5892 , n5982 );
or ( n5984 , n5891 , n5983 );
and ( n5985 , n5888 , n5984 );
or ( n5986 , n5887 , n5985 );
and ( n5987 , n5884 , n5986 );
or ( n5988 , n5883 , n5987 );
and ( n5989 , n5880 , n5988 );
or ( n5990 , n5879 , n5989 );
and ( n5991 , n5876 , n5990 );
or ( n5992 , n5875 , n5991 );
and ( n5993 , n5872 , n5992 );
or ( n5994 , n5871 , n5993 );
and ( n5995 , n5868 , n5994 );
or ( n5996 , n5867 , n5995 );
xor ( n5997 , n5864 , n5996 );
and ( n5998 , n285 , n1125 );
nor ( n5999 , n1126 , n5998 );
nor ( n6000 , n1318 , n305 );
xor ( n6001 , n5999 , n6000 );
and ( n6002 , n5595 , n5596 );
and ( n6003 , n5597 , n5600 );
or ( n6004 , n6002 , n6003 );
xor ( n6005 , n6001 , n6004 );
nor ( n6006 , n1534 , n336 );
xor ( n6007 , n6005 , n6006 );
and ( n6008 , n5601 , n5602 );
and ( n6009 , n5603 , n5606 );
or ( n6010 , n6008 , n6009 );
xor ( n6011 , n6007 , n6010 );
nor ( n6012 , n1771 , n386 );
xor ( n6013 , n6011 , n6012 );
and ( n6014 , n5607 , n5608 );
and ( n6015 , n5609 , n5612 );
or ( n6016 , n6014 , n6015 );
xor ( n6017 , n6013 , n6016 );
nor ( n6018 , n2025 , n458 );
xor ( n6019 , n6017 , n6018 );
and ( n6020 , n5613 , n5614 );
and ( n6021 , n5615 , n5618 );
or ( n6022 , n6020 , n6021 );
xor ( n6023 , n6019 , n6022 );
nor ( n6024 , n2300 , n551 );
xor ( n6025 , n6023 , n6024 );
and ( n6026 , n5619 , n5620 );
and ( n6027 , n5621 , n5624 );
or ( n6028 , n6026 , n6027 );
xor ( n6029 , n6025 , n6028 );
nor ( n6030 , n2596 , n665 );
xor ( n6031 , n6029 , n6030 );
and ( n6032 , n5625 , n5626 );
and ( n6033 , n5627 , n5630 );
or ( n6034 , n6032 , n6033 );
xor ( n6035 , n6031 , n6034 );
nor ( n6036 , n2991 , n797 );
xor ( n6037 , n6035 , n6036 );
and ( n6038 , n5631 , n5632 );
and ( n6039 , n5633 , n5636 );
or ( n6040 , n6038 , n6039 );
xor ( n6041 , n6037 , n6040 );
nor ( n6042 , n3464 , n954 );
xor ( n6043 , n6041 , n6042 );
and ( n6044 , n5637 , n5638 );
and ( n6045 , n5639 , n5642 );
or ( n6046 , n6044 , n6045 );
xor ( n6047 , n6043 , n6046 );
nor ( n6048 , n3863 , n1128 );
xor ( n6049 , n6047 , n6048 );
and ( n6050 , n5643 , n5644 );
and ( n6051 , n5645 , n5648 );
or ( n6052 , n6050 , n6051 );
xor ( n6053 , n6049 , n6052 );
nor ( n6054 , n4260 , n1320 );
xor ( n6055 , n6053 , n6054 );
and ( n6056 , n5649 , n5650 );
and ( n6057 , n5651 , n5654 );
or ( n6058 , n6056 , n6057 );
xor ( n6059 , n6055 , n6058 );
nor ( n6060 , n4659 , n1536 );
xor ( n6061 , n6059 , n6060 );
and ( n6062 , n5655 , n5656 );
and ( n6063 , n5657 , n5660 );
or ( n6064 , n6062 , n6063 );
xor ( n6065 , n6061 , n6064 );
nor ( n6066 , n5057 , n1773 );
xor ( n6067 , n6065 , n6066 );
and ( n6068 , n5661 , n5662 );
and ( n6069 , n5663 , n5666 );
or ( n6070 , n6068 , n6069 );
xor ( n6071 , n6067 , n6070 );
nor ( n6072 , n5453 , n2027 );
xor ( n6073 , n6071 , n6072 );
and ( n6074 , n5667 , n5668 );
and ( n6075 , n5669 , n5672 );
or ( n6076 , n6074 , n6075 );
xor ( n6077 , n6073 , n6076 );
nor ( n6078 , n5851 , n2302 );
xor ( n6079 , n6077 , n6078 );
and ( n6080 , n5673 , n5674 );
and ( n6081 , n5675 , n5678 );
or ( n6082 , n6080 , n6081 );
xor ( n6083 , n6079 , n6082 );
and ( n6084 , n5696 , n5700 );
and ( n6085 , n5700 , n5704 );
and ( n6086 , n5696 , n5704 );
or ( n6087 , n6084 , n6085 , n6086 );
and ( n6088 , n5692 , n5705 );
and ( n6089 , n5705 , n5837 );
and ( n6090 , n5692 , n5837 );
or ( n6091 , n6088 , n6089 , n6090 );
xor ( n6092 , n6087 , n6091 );
and ( n6093 , n5710 , n5736 );
and ( n6094 , n5736 , n5836 );
and ( n6095 , n5710 , n5836 );
or ( n6096 , n6093 , n6094 , n6095 );
and ( n6097 , n5724 , n5725 );
and ( n6098 , n5725 , n5727 );
and ( n6099 , n5724 , n5727 );
or ( n6100 , n6097 , n6098 , n6099 );
and ( n6101 , n5714 , n5718 );
and ( n6102 , n5718 , n5735 );
and ( n6103 , n5714 , n5735 );
or ( n6104 , n6101 , n6102 , n6103 );
xor ( n6105 , n6100 , n6104 );
not ( n6106 , n1088 );
and ( n6107 , n2406 , n1088 );
nor ( n6108 , n6106 , n6107 );
xor ( n6109 , n6105 , n6108 );
xor ( n6110 , n6096 , n6109 );
and ( n6111 , n5741 , n5756 );
and ( n6112 , n5756 , n5835 );
and ( n6113 , n5741 , n5835 );
or ( n6114 , n6111 , n6112 , n6113 );
and ( n6115 , n5723 , n5728 );
and ( n6116 , n5728 , n5734 );
and ( n6117 , n5723 , n5734 );
or ( n6118 , n6115 , n6116 , n6117 );
and ( n6119 , n5745 , n5749 );
and ( n6120 , n5749 , n5755 );
and ( n6121 , n5745 , n5755 );
or ( n6122 , n6119 , n6120 , n6121 );
xor ( n6123 , n6118 , n6122 );
and ( n6124 , n5730 , n5731 );
and ( n6125 , n5731 , n5733 );
and ( n6126 , n5730 , n5733 );
or ( n6127 , n6124 , n6125 , n6126 );
and ( n6128 , n1292 , n2138 );
and ( n6129 , n1516 , n1864 );
xor ( n6130 , n6128 , n6129 );
and ( n6131 , n1730 , n1753 );
xor ( n6132 , n6130 , n6131 );
xor ( n6133 , n6127 , n6132 );
and ( n6134 , n2001 , n1396 );
and ( n6135 , n2286 , n1302 );
xor ( n6136 , n6134 , n6135 );
and ( n6137 , n2581 , n1114 );
xor ( n6138 , n6136 , n6137 );
xor ( n6139 , n6133 , n6138 );
xor ( n6140 , n6123 , n6139 );
xor ( n6141 , n6114 , n6140 );
and ( n6142 , n5761 , n5766 );
and ( n6143 , n5766 , n5834 );
and ( n6144 , n5761 , n5834 );
or ( n6145 , n6142 , n6143 , n6144 );
and ( n6146 , n5751 , n5752 );
and ( n6147 , n5752 , n5754 );
and ( n6148 , n5751 , n5754 );
or ( n6149 , n6146 , n6147 , n6148 );
and ( n6150 , n5762 , n5763 );
and ( n6151 , n5763 , n5765 );
and ( n6152 , n5762 , n5765 );
or ( n6153 , n6150 , n6151 , n6152 );
xor ( n6154 , n6149 , n6153 );
and ( n6155 , n2972 , n852 );
and ( n6156 , n3445 , n714 );
xor ( n6157 , n6155 , n6156 );
and ( n6158 , n3844 , n651 );
xor ( n6159 , n6157 , n6158 );
xor ( n6160 , n6154 , n6159 );
xor ( n6161 , n6145 , n6160 );
and ( n6162 , n5768 , n5769 );
and ( n6163 , n5769 , n5833 );
and ( n6164 , n5768 , n5833 );
or ( n6165 , n6162 , n6163 , n6164 );
and ( n6166 , n4241 , n488 );
and ( n6167 , n4640 , n411 );
xor ( n6168 , n6166 , n6167 );
and ( n6169 , n5038 , n375 );
xor ( n6170 , n6168 , n6169 );
xor ( n6171 , n6165 , n6170 );
and ( n6172 , n5434 , n312 );
and ( n6173 , n5832 , n288 );
xor ( n6174 , n6172 , n6173 );
and ( n6175 , n5784 , n5788 );
and ( n6176 , n5788 , n5792 );
and ( n6177 , n5784 , n5792 );
or ( n6178 , n6175 , n6176 , n6177 );
and ( n6179 , n5780 , n5793 );
and ( n6180 , n5793 , n5819 );
and ( n6181 , n5780 , n5819 );
or ( n6182 , n6179 , n6180 , n6181 );
xor ( n6183 , n6178 , n6182 );
and ( n6184 , n5805 , n5806 );
and ( n6185 , n5806 , n5808 );
and ( n6186 , n5805 , n5808 );
or ( n6187 , n6184 , n6185 , n6186 );
and ( n6188 , n5798 , n5799 );
and ( n6189 , n5799 , n5818 );
and ( n6190 , n5798 , n5818 );
or ( n6191 , n6188 , n6189 , n6190 );
xor ( n6192 , n6187 , n6191 );
and ( n6193 , n2206 , n1261 );
not ( n6194 , n1261 );
nor ( n6195 , n6193 , n6194 );
xor ( n6196 , n6192 , n6195 );
and ( n6197 , n5804 , n5809 );
and ( n6198 , n5809 , n5817 );
and ( n6199 , n5804 , n5817 );
or ( n6200 , n6197 , n6198 , n6199 );
and ( n6201 , n5813 , n5814 );
and ( n6202 , n5814 , n5816 );
and ( n6203 , n5813 , n5816 );
or ( n6204 , n6201 , n6202 , n6203 );
and ( n6205 , n1458 , n1975 );
and ( n6206 , n1713 , n1685 );
xor ( n6207 , n6205 , n6206 );
and ( n6208 , n1935 , n1497 );
xor ( n6209 , n6207 , n6208 );
xor ( n6210 , n6204 , n6209 );
not ( n6211 , n1077 );
and ( n6212 , n2563 , n1077 );
nor ( n6213 , n6211 , n6212 );
and ( n6214 , n1277 , n2271 );
xor ( n6215 , n6213 , n6214 );
xor ( n6216 , n6210 , n6215 );
xor ( n6217 , n6200 , n6216 );
xor ( n6218 , n6196 , n6217 );
xor ( n6219 , n6183 , n6218 );
and ( n6220 , n5774 , n5778 );
and ( n6221 , n5778 , n5820 );
and ( n6222 , n5774 , n5820 );
or ( n6223 , n6220 , n6221 , n6222 );
xor ( n6224 , n6219 , n6223 );
and ( n6225 , n5821 , n5825 );
and ( n6226 , n5826 , n5829 );
or ( n6227 , n6225 , n6226 );
xor ( n6228 , n6224 , n6227 );
buf ( n6229 , n6228 );
buf ( n6230 , n6229 );
and ( n6231 , n6230 , n279 );
xor ( n6232 , n6174 , n6231 );
xor ( n6233 , n6171 , n6232 );
xor ( n6234 , n6161 , n6233 );
xor ( n6235 , n6141 , n6234 );
xor ( n6236 , n6110 , n6235 );
xor ( n6237 , n6092 , n6236 );
and ( n6238 , n5683 , n5687 );
and ( n6239 , n5687 , n5838 );
and ( n6240 , n5683 , n5838 );
or ( n6241 , n6238 , n6239 , n6240 );
xor ( n6242 , n6237 , n6241 );
and ( n6243 , n5839 , n5843 );
and ( n6244 , n5844 , n5847 );
or ( n6245 , n6243 , n6244 );
xor ( n6246 , n6242 , n6245 );
buf ( n6247 , n6246 );
buf ( n6248 , n6247 );
not ( n6249 , n6248 );
nor ( n6250 , n6249 , n2598 );
xor ( n6251 , n6083 , n6250 );
and ( n6252 , n5679 , n5852 );
and ( n6253 , n5853 , n5856 );
or ( n6254 , n6252 , n6253 );
xor ( n6255 , n6251 , n6254 );
buf ( n6256 , n6255 );
buf ( n6257 , n6256 );
not ( n6258 , n6257 );
buf ( n6259 , n266 );
not ( n6260 , n6259 );
nor ( n6261 , n6258 , n6260 );
xor ( n6262 , n5997 , n6261 );
xor ( n6263 , n5868 , n5994 );
nor ( n6264 , n5860 , n6260 );
and ( n6265 , n6263 , n6264 );
xor ( n6266 , n6263 , n6264 );
xor ( n6267 , n5872 , n5992 );
nor ( n6268 , n5462 , n6260 );
and ( n6269 , n6267 , n6268 );
xor ( n6270 , n6267 , n6268 );
xor ( n6271 , n5876 , n5990 );
nor ( n6272 , n5066 , n6260 );
and ( n6273 , n6271 , n6272 );
xor ( n6274 , n6271 , n6272 );
xor ( n6275 , n5880 , n5988 );
nor ( n6276 , n4668 , n6260 );
and ( n6277 , n6275 , n6276 );
xor ( n6278 , n6275 , n6276 );
xor ( n6279 , n5884 , n5986 );
nor ( n6280 , n4269 , n6260 );
and ( n6281 , n6279 , n6280 );
xor ( n6282 , n6279 , n6280 );
xor ( n6283 , n5888 , n5984 );
nor ( n6284 , n3872 , n6260 );
and ( n6285 , n6283 , n6284 );
xor ( n6286 , n6283 , n6284 );
xor ( n6287 , n5892 , n5982 );
nor ( n6288 , n3473 , n6260 );
and ( n6289 , n6287 , n6288 );
xor ( n6290 , n6287 , n6288 );
xor ( n6291 , n5896 , n5980 );
nor ( n6292 , n3000 , n6260 );
and ( n6293 , n6291 , n6292 );
xor ( n6294 , n6291 , n6292 );
xor ( n6295 , n5900 , n5978 );
nor ( n6296 , n2688 , n6260 );
and ( n6297 , n6295 , n6296 );
xor ( n6298 , n6295 , n6296 );
xor ( n6299 , n5904 , n5976 );
nor ( n6300 , n3008 , n6260 );
and ( n6301 , n6299 , n6300 );
xor ( n6302 , n6299 , n6300 );
xor ( n6303 , n5908 , n5974 );
nor ( n6304 , n3017 , n6260 );
and ( n6305 , n6303 , n6304 );
xor ( n6306 , n6303 , n6304 );
xor ( n6307 , n5912 , n5972 );
nor ( n6308 , n3026 , n6260 );
and ( n6309 , n6307 , n6308 );
xor ( n6310 , n6307 , n6308 );
xor ( n6311 , n5916 , n5970 );
nor ( n6312 , n3035 , n6260 );
and ( n6313 , n6311 , n6312 );
xor ( n6314 , n6311 , n6312 );
xor ( n6315 , n5920 , n5968 );
nor ( n6316 , n3044 , n6260 );
and ( n6317 , n6315 , n6316 );
xor ( n6318 , n6315 , n6316 );
xor ( n6319 , n5924 , n5966 );
nor ( n6320 , n3053 , n6260 );
and ( n6321 , n6319 , n6320 );
xor ( n6322 , n6319 , n6320 );
xor ( n6323 , n5928 , n5964 );
nor ( n6324 , n3062 , n6260 );
and ( n6325 , n6323 , n6324 );
xor ( n6326 , n6323 , n6324 );
xor ( n6327 , n5932 , n5962 );
nor ( n6328 , n3071 , n6260 );
and ( n6329 , n6327 , n6328 );
xor ( n6330 , n6327 , n6328 );
xor ( n6331 , n5936 , n5960 );
nor ( n6332 , n3080 , n6260 );
and ( n6333 , n6331 , n6332 );
xor ( n6334 , n6331 , n6332 );
xor ( n6335 , n5940 , n5958 );
nor ( n6336 , n3089 , n6260 );
and ( n6337 , n6335 , n6336 );
xor ( n6338 , n6335 , n6336 );
xor ( n6339 , n5944 , n5956 );
nor ( n6340 , n3098 , n6260 );
and ( n6341 , n6339 , n6340 );
xor ( n6342 , n6339 , n6340 );
xor ( n6343 , n5949 , n5954 );
nor ( n6344 , n3107 , n6260 );
and ( n6345 , n6343 , n6344 );
xor ( n6346 , n6343 , n6344 );
xor ( n6347 , n5951 , n5952 );
buf ( n6348 , n6347 );
nor ( n6349 , n3116 , n6260 );
and ( n6350 , n6348 , n6349 );
xor ( n6351 , n6348 , n6349 );
nor ( n6352 , n3134 , n5862 );
buf ( n6353 , n6352 );
nor ( n6354 , n3125 , n6260 );
and ( n6355 , n6353 , n6354 );
buf ( n6356 , n6355 );
and ( n6357 , n6351 , n6356 );
or ( n6358 , n6350 , n6357 );
and ( n6359 , n6346 , n6358 );
or ( n6360 , n6345 , n6359 );
and ( n6361 , n6342 , n6360 );
or ( n6362 , n6341 , n6361 );
and ( n6363 , n6338 , n6362 );
or ( n6364 , n6337 , n6363 );
and ( n6365 , n6334 , n6364 );
or ( n6366 , n6333 , n6365 );
and ( n6367 , n6330 , n6366 );
or ( n6368 , n6329 , n6367 );
and ( n6369 , n6326 , n6368 );
or ( n6370 , n6325 , n6369 );
and ( n6371 , n6322 , n6370 );
or ( n6372 , n6321 , n6371 );
and ( n6373 , n6318 , n6372 );
or ( n6374 , n6317 , n6373 );
and ( n6375 , n6314 , n6374 );
or ( n6376 , n6313 , n6375 );
and ( n6377 , n6310 , n6376 );
or ( n6378 , n6309 , n6377 );
and ( n6379 , n6306 , n6378 );
or ( n6380 , n6305 , n6379 );
and ( n6381 , n6302 , n6380 );
or ( n6382 , n6301 , n6381 );
and ( n6383 , n6298 , n6382 );
or ( n6384 , n6297 , n6383 );
and ( n6385 , n6294 , n6384 );
or ( n6386 , n6293 , n6385 );
and ( n6387 , n6290 , n6386 );
or ( n6388 , n6289 , n6387 );
and ( n6389 , n6286 , n6388 );
or ( n6390 , n6285 , n6389 );
and ( n6391 , n6282 , n6390 );
or ( n6392 , n6281 , n6391 );
and ( n6393 , n6278 , n6392 );
or ( n6394 , n6277 , n6393 );
and ( n6395 , n6274 , n6394 );
or ( n6396 , n6273 , n6395 );
and ( n6397 , n6270 , n6396 );
or ( n6398 , n6269 , n6397 );
and ( n6399 , n6266 , n6398 );
or ( n6400 , n6265 , n6399 );
xor ( n6401 , n6262 , n6400 );
and ( n6402 , n285 , n1317 );
nor ( n6403 , n1318 , n6402 );
nor ( n6404 , n1534 , n305 );
xor ( n6405 , n6403 , n6404 );
and ( n6406 , n5999 , n6000 );
and ( n6407 , n6001 , n6004 );
or ( n6408 , n6406 , n6407 );
xor ( n6409 , n6405 , n6408 );
nor ( n6410 , n1771 , n336 );
xor ( n6411 , n6409 , n6410 );
and ( n6412 , n6005 , n6006 );
and ( n6413 , n6007 , n6010 );
or ( n6414 , n6412 , n6413 );
xor ( n6415 , n6411 , n6414 );
nor ( n6416 , n2025 , n386 );
xor ( n6417 , n6415 , n6416 );
and ( n6418 , n6011 , n6012 );
and ( n6419 , n6013 , n6016 );
or ( n6420 , n6418 , n6419 );
xor ( n6421 , n6417 , n6420 );
nor ( n6422 , n2300 , n458 );
xor ( n6423 , n6421 , n6422 );
and ( n6424 , n6017 , n6018 );
and ( n6425 , n6019 , n6022 );
or ( n6426 , n6424 , n6425 );
xor ( n6427 , n6423 , n6426 );
nor ( n6428 , n2596 , n551 );
xor ( n6429 , n6427 , n6428 );
and ( n6430 , n6023 , n6024 );
and ( n6431 , n6025 , n6028 );
or ( n6432 , n6430 , n6431 );
xor ( n6433 , n6429 , n6432 );
nor ( n6434 , n2991 , n665 );
xor ( n6435 , n6433 , n6434 );
and ( n6436 , n6029 , n6030 );
and ( n6437 , n6031 , n6034 );
or ( n6438 , n6436 , n6437 );
xor ( n6439 , n6435 , n6438 );
nor ( n6440 , n3464 , n797 );
xor ( n6441 , n6439 , n6440 );
and ( n6442 , n6035 , n6036 );
and ( n6443 , n6037 , n6040 );
or ( n6444 , n6442 , n6443 );
xor ( n6445 , n6441 , n6444 );
nor ( n6446 , n3863 , n954 );
xor ( n6447 , n6445 , n6446 );
and ( n6448 , n6041 , n6042 );
and ( n6449 , n6043 , n6046 );
or ( n6450 , n6448 , n6449 );
xor ( n6451 , n6447 , n6450 );
nor ( n6452 , n4260 , n1128 );
xor ( n6453 , n6451 , n6452 );
and ( n6454 , n6047 , n6048 );
and ( n6455 , n6049 , n6052 );
or ( n6456 , n6454 , n6455 );
xor ( n6457 , n6453 , n6456 );
nor ( n6458 , n4659 , n1320 );
xor ( n6459 , n6457 , n6458 );
and ( n6460 , n6053 , n6054 );
and ( n6461 , n6055 , n6058 );
or ( n6462 , n6460 , n6461 );
xor ( n6463 , n6459 , n6462 );
nor ( n6464 , n5057 , n1536 );
xor ( n6465 , n6463 , n6464 );
and ( n6466 , n6059 , n6060 );
and ( n6467 , n6061 , n6064 );
or ( n6468 , n6466 , n6467 );
xor ( n6469 , n6465 , n6468 );
nor ( n6470 , n5453 , n1773 );
xor ( n6471 , n6469 , n6470 );
and ( n6472 , n6065 , n6066 );
and ( n6473 , n6067 , n6070 );
or ( n6474 , n6472 , n6473 );
xor ( n6475 , n6471 , n6474 );
nor ( n6476 , n5851 , n2027 );
xor ( n6477 , n6475 , n6476 );
and ( n6478 , n6071 , n6072 );
and ( n6479 , n6073 , n6076 );
or ( n6480 , n6478 , n6479 );
xor ( n6481 , n6477 , n6480 );
nor ( n6482 , n6249 , n2302 );
xor ( n6483 , n6481 , n6482 );
and ( n6484 , n6077 , n6078 );
and ( n6485 , n6079 , n6082 );
or ( n6486 , n6484 , n6485 );
xor ( n6487 , n6483 , n6486 );
and ( n6488 , n6100 , n6104 );
and ( n6489 , n6104 , n6108 );
and ( n6490 , n6100 , n6108 );
or ( n6491 , n6488 , n6489 , n6490 );
and ( n6492 , n6096 , n6109 );
and ( n6493 , n6109 , n6235 );
and ( n6494 , n6096 , n6235 );
or ( n6495 , n6492 , n6493 , n6494 );
xor ( n6496 , n6491 , n6495 );
and ( n6497 , n6114 , n6140 );
and ( n6498 , n6140 , n6234 );
and ( n6499 , n6114 , n6234 );
or ( n6500 , n6497 , n6498 , n6499 );
and ( n6501 , n6128 , n6129 );
and ( n6502 , n6129 , n6131 );
and ( n6503 , n6128 , n6131 );
or ( n6504 , n6501 , n6502 , n6503 );
and ( n6505 , n6118 , n6122 );
and ( n6506 , n6122 , n6139 );
and ( n6507 , n6118 , n6139 );
or ( n6508 , n6505 , n6506 , n6507 );
xor ( n6509 , n6504 , n6508 );
not ( n6510 , n1292 );
and ( n6511 , n2406 , n1292 );
nor ( n6512 , n6510 , n6511 );
xor ( n6513 , n6509 , n6512 );
xor ( n6514 , n6500 , n6513 );
and ( n6515 , n6145 , n6160 );
and ( n6516 , n6160 , n6233 );
and ( n6517 , n6145 , n6233 );
or ( n6518 , n6515 , n6516 , n6517 );
and ( n6519 , n6127 , n6132 );
and ( n6520 , n6132 , n6138 );
and ( n6521 , n6127 , n6138 );
or ( n6522 , n6519 , n6520 , n6521 );
and ( n6523 , n6149 , n6153 );
and ( n6524 , n6153 , n6159 );
and ( n6525 , n6149 , n6159 );
or ( n6526 , n6523 , n6524 , n6525 );
xor ( n6527 , n6522 , n6526 );
and ( n6528 , n6134 , n6135 );
and ( n6529 , n6135 , n6137 );
and ( n6530 , n6134 , n6137 );
or ( n6531 , n6528 , n6529 , n6530 );
and ( n6532 , n1516 , n2138 );
and ( n6533 , n1730 , n1864 );
xor ( n6534 , n6532 , n6533 );
and ( n6535 , n2001 , n1753 );
xor ( n6536 , n6534 , n6535 );
xor ( n6537 , n6531 , n6536 );
and ( n6538 , n2286 , n1396 );
and ( n6539 , n2581 , n1302 );
xor ( n6540 , n6538 , n6539 );
and ( n6541 , n2972 , n1114 );
xor ( n6542 , n6540 , n6541 );
xor ( n6543 , n6537 , n6542 );
xor ( n6544 , n6527 , n6543 );
xor ( n6545 , n6518 , n6544 );
and ( n6546 , n6165 , n6170 );
and ( n6547 , n6170 , n6232 );
and ( n6548 , n6165 , n6232 );
or ( n6549 , n6546 , n6547 , n6548 );
and ( n6550 , n6155 , n6156 );
and ( n6551 , n6156 , n6158 );
and ( n6552 , n6155 , n6158 );
or ( n6553 , n6550 , n6551 , n6552 );
and ( n6554 , n6166 , n6167 );
and ( n6555 , n6167 , n6169 );
and ( n6556 , n6166 , n6169 );
or ( n6557 , n6554 , n6555 , n6556 );
xor ( n6558 , n6553 , n6557 );
and ( n6559 , n3445 , n852 );
and ( n6560 , n3844 , n714 );
xor ( n6561 , n6559 , n6560 );
and ( n6562 , n4241 , n651 );
xor ( n6563 , n6561 , n6562 );
xor ( n6564 , n6558 , n6563 );
xor ( n6565 , n6549 , n6564 );
and ( n6566 , n6172 , n6173 );
and ( n6567 , n6173 , n6231 );
and ( n6568 , n6172 , n6231 );
or ( n6569 , n6566 , n6567 , n6568 );
and ( n6570 , n4640 , n488 );
and ( n6571 , n5038 , n411 );
xor ( n6572 , n6570 , n6571 );
and ( n6573 , n5434 , n375 );
xor ( n6574 , n6572 , n6573 );
xor ( n6575 , n6569 , n6574 );
and ( n6576 , n5832 , n312 );
and ( n6577 , n6230 , n288 );
xor ( n6578 , n6576 , n6577 );
and ( n6579 , n6187 , n6191 );
and ( n6580 , n6191 , n6195 );
and ( n6581 , n6187 , n6195 );
or ( n6582 , n6579 , n6580 , n6581 );
and ( n6583 , n6196 , n6217 );
xor ( n6584 , n6582 , n6583 );
and ( n6585 , n6205 , n6206 );
and ( n6586 , n6206 , n6208 );
and ( n6587 , n6205 , n6208 );
or ( n6588 , n6585 , n6586 , n6587 );
and ( n6589 , n6200 , n6216 );
xor ( n6590 , n6588 , n6589 );
and ( n6591 , n2206 , n1497 );
not ( n6592 , n1497 );
nor ( n6593 , n6591 , n6592 );
xor ( n6594 , n6590 , n6593 );
and ( n6595 , n6204 , n6209 );
and ( n6596 , n6209 , n6215 );
and ( n6597 , n6204 , n6215 );
or ( n6598 , n6595 , n6596 , n6597 );
and ( n6599 , n6213 , n6214 );
not ( n6600 , n1277 );
and ( n6601 , n2563 , n1277 );
nor ( n6602 , n6600 , n6601 );
xor ( n6603 , n6599 , n6602 );
and ( n6604 , n1458 , n2271 );
and ( n6605 , n1713 , n1975 );
xor ( n6606 , n6604 , n6605 );
and ( n6607 , n1935 , n1685 );
xor ( n6608 , n6606 , n6607 );
xor ( n6609 , n6603 , n6608 );
xor ( n6610 , n6598 , n6609 );
xor ( n6611 , n6594 , n6610 );
xor ( n6612 , n6584 , n6611 );
and ( n6613 , n6178 , n6182 );
and ( n6614 , n6182 , n6218 );
and ( n6615 , n6178 , n6218 );
or ( n6616 , n6613 , n6614 , n6615 );
xor ( n6617 , n6612 , n6616 );
and ( n6618 , n6219 , n6223 );
and ( n6619 , n6224 , n6227 );
or ( n6620 , n6618 , n6619 );
xor ( n6621 , n6617 , n6620 );
buf ( n6622 , n6621 );
buf ( n6623 , n6622 );
and ( n6624 , n6623 , n279 );
xor ( n6625 , n6578 , n6624 );
xor ( n6626 , n6575 , n6625 );
xor ( n6627 , n6565 , n6626 );
xor ( n6628 , n6545 , n6627 );
xor ( n6629 , n6514 , n6628 );
xor ( n6630 , n6496 , n6629 );
and ( n6631 , n6087 , n6091 );
and ( n6632 , n6091 , n6236 );
and ( n6633 , n6087 , n6236 );
or ( n6634 , n6631 , n6632 , n6633 );
xor ( n6635 , n6630 , n6634 );
and ( n6636 , n6237 , n6241 );
and ( n6637 , n6242 , n6245 );
or ( n6638 , n6636 , n6637 );
xor ( n6639 , n6635 , n6638 );
buf ( n6640 , n6639 );
buf ( n6641 , n6640 );
not ( n6642 , n6641 );
nor ( n6643 , n6642 , n2598 );
xor ( n6644 , n6487 , n6643 );
and ( n6645 , n6083 , n6250 );
and ( n6646 , n6251 , n6254 );
or ( n6647 , n6645 , n6646 );
xor ( n6648 , n6644 , n6647 );
buf ( n6649 , n6648 );
buf ( n6650 , n6649 );
not ( n6651 , n6650 );
buf ( n6652 , n267 );
not ( n6653 , n6652 );
nor ( n6654 , n6651 , n6653 );
xor ( n6655 , n6401 , n6654 );
xor ( n6656 , n6266 , n6398 );
nor ( n6657 , n6258 , n6653 );
and ( n6658 , n6656 , n6657 );
xor ( n6659 , n6656 , n6657 );
xor ( n6660 , n6270 , n6396 );
nor ( n6661 , n5860 , n6653 );
and ( n6662 , n6660 , n6661 );
xor ( n6663 , n6660 , n6661 );
xor ( n6664 , n6274 , n6394 );
nor ( n6665 , n5462 , n6653 );
and ( n6666 , n6664 , n6665 );
xor ( n6667 , n6664 , n6665 );
xor ( n6668 , n6278 , n6392 );
nor ( n6669 , n5066 , n6653 );
and ( n6670 , n6668 , n6669 );
xor ( n6671 , n6668 , n6669 );
xor ( n6672 , n6282 , n6390 );
nor ( n6673 , n4668 , n6653 );
and ( n6674 , n6672 , n6673 );
xor ( n6675 , n6672 , n6673 );
xor ( n6676 , n6286 , n6388 );
nor ( n6677 , n4269 , n6653 );
and ( n6678 , n6676 , n6677 );
xor ( n6679 , n6676 , n6677 );
xor ( n6680 , n6290 , n6386 );
nor ( n6681 , n3872 , n6653 );
and ( n6682 , n6680 , n6681 );
xor ( n6683 , n6680 , n6681 );
xor ( n6684 , n6294 , n6384 );
nor ( n6685 , n3473 , n6653 );
and ( n6686 , n6684 , n6685 );
xor ( n6687 , n6684 , n6685 );
xor ( n6688 , n6298 , n6382 );
nor ( n6689 , n3000 , n6653 );
and ( n6690 , n6688 , n6689 );
xor ( n6691 , n6688 , n6689 );
xor ( n6692 , n6302 , n6380 );
nor ( n6693 , n2688 , n6653 );
and ( n6694 , n6692 , n6693 );
xor ( n6695 , n6692 , n6693 );
xor ( n6696 , n6306 , n6378 );
nor ( n6697 , n3008 , n6653 );
and ( n6698 , n6696 , n6697 );
xor ( n6699 , n6696 , n6697 );
xor ( n6700 , n6310 , n6376 );
nor ( n6701 , n3017 , n6653 );
and ( n6702 , n6700 , n6701 );
xor ( n6703 , n6700 , n6701 );
xor ( n6704 , n6314 , n6374 );
nor ( n6705 , n3026 , n6653 );
and ( n6706 , n6704 , n6705 );
xor ( n6707 , n6704 , n6705 );
xor ( n6708 , n6318 , n6372 );
nor ( n6709 , n3035 , n6653 );
and ( n6710 , n6708 , n6709 );
xor ( n6711 , n6708 , n6709 );
xor ( n6712 , n6322 , n6370 );
nor ( n6713 , n3044 , n6653 );
and ( n6714 , n6712 , n6713 );
xor ( n6715 , n6712 , n6713 );
xor ( n6716 , n6326 , n6368 );
nor ( n6717 , n3053 , n6653 );
and ( n6718 , n6716 , n6717 );
xor ( n6719 , n6716 , n6717 );
xor ( n6720 , n6330 , n6366 );
nor ( n6721 , n3062 , n6653 );
and ( n6722 , n6720 , n6721 );
xor ( n6723 , n6720 , n6721 );
xor ( n6724 , n6334 , n6364 );
nor ( n6725 , n3071 , n6653 );
and ( n6726 , n6724 , n6725 );
xor ( n6727 , n6724 , n6725 );
xor ( n6728 , n6338 , n6362 );
nor ( n6729 , n3080 , n6653 );
and ( n6730 , n6728 , n6729 );
xor ( n6731 , n6728 , n6729 );
xor ( n6732 , n6342 , n6360 );
nor ( n6733 , n3089 , n6653 );
and ( n6734 , n6732 , n6733 );
xor ( n6735 , n6732 , n6733 );
xor ( n6736 , n6346 , n6358 );
nor ( n6737 , n3098 , n6653 );
and ( n6738 , n6736 , n6737 );
xor ( n6739 , n6736 , n6737 );
xor ( n6740 , n6351 , n6356 );
nor ( n6741 , n3107 , n6653 );
and ( n6742 , n6740 , n6741 );
xor ( n6743 , n6740 , n6741 );
xor ( n6744 , n6353 , n6354 );
buf ( n6745 , n6744 );
nor ( n6746 , n3116 , n6653 );
and ( n6747 , n6745 , n6746 );
xor ( n6748 , n6745 , n6746 );
nor ( n6749 , n3134 , n6260 );
buf ( n6750 , n6749 );
nor ( n6751 , n3125 , n6653 );
and ( n6752 , n6750 , n6751 );
buf ( n6753 , n6752 );
and ( n6754 , n6748 , n6753 );
or ( n6755 , n6747 , n6754 );
and ( n6756 , n6743 , n6755 );
or ( n6757 , n6742 , n6756 );
and ( n6758 , n6739 , n6757 );
or ( n6759 , n6738 , n6758 );
and ( n6760 , n6735 , n6759 );
or ( n6761 , n6734 , n6760 );
and ( n6762 , n6731 , n6761 );
or ( n6763 , n6730 , n6762 );
and ( n6764 , n6727 , n6763 );
or ( n6765 , n6726 , n6764 );
and ( n6766 , n6723 , n6765 );
or ( n6767 , n6722 , n6766 );
and ( n6768 , n6719 , n6767 );
or ( n6769 , n6718 , n6768 );
and ( n6770 , n6715 , n6769 );
or ( n6771 , n6714 , n6770 );
and ( n6772 , n6711 , n6771 );
or ( n6773 , n6710 , n6772 );
and ( n6774 , n6707 , n6773 );
or ( n6775 , n6706 , n6774 );
and ( n6776 , n6703 , n6775 );
or ( n6777 , n6702 , n6776 );
and ( n6778 , n6699 , n6777 );
or ( n6779 , n6698 , n6778 );
and ( n6780 , n6695 , n6779 );
or ( n6781 , n6694 , n6780 );
and ( n6782 , n6691 , n6781 );
or ( n6783 , n6690 , n6782 );
and ( n6784 , n6687 , n6783 );
or ( n6785 , n6686 , n6784 );
and ( n6786 , n6683 , n6785 );
or ( n6787 , n6682 , n6786 );
and ( n6788 , n6679 , n6787 );
or ( n6789 , n6678 , n6788 );
and ( n6790 , n6675 , n6789 );
or ( n6791 , n6674 , n6790 );
and ( n6792 , n6671 , n6791 );
or ( n6793 , n6670 , n6792 );
and ( n6794 , n6667 , n6793 );
or ( n6795 , n6666 , n6794 );
and ( n6796 , n6663 , n6795 );
or ( n6797 , n6662 , n6796 );
and ( n6798 , n6659 , n6797 );
or ( n6799 , n6658 , n6798 );
xor ( n6800 , n6655 , n6799 );
and ( n6801 , n285 , n1533 );
nor ( n6802 , n1534 , n6801 );
nor ( n6803 , n1771 , n305 );
xor ( n6804 , n6802 , n6803 );
and ( n6805 , n6403 , n6404 );
and ( n6806 , n6405 , n6408 );
or ( n6807 , n6805 , n6806 );
xor ( n6808 , n6804 , n6807 );
nor ( n6809 , n2025 , n336 );
xor ( n6810 , n6808 , n6809 );
and ( n6811 , n6409 , n6410 );
and ( n6812 , n6411 , n6414 );
or ( n6813 , n6811 , n6812 );
xor ( n6814 , n6810 , n6813 );
nor ( n6815 , n2300 , n386 );
xor ( n6816 , n6814 , n6815 );
and ( n6817 , n6415 , n6416 );
and ( n6818 , n6417 , n6420 );
or ( n6819 , n6817 , n6818 );
xor ( n6820 , n6816 , n6819 );
nor ( n6821 , n2596 , n458 );
xor ( n6822 , n6820 , n6821 );
and ( n6823 , n6421 , n6422 );
and ( n6824 , n6423 , n6426 );
or ( n6825 , n6823 , n6824 );
xor ( n6826 , n6822 , n6825 );
nor ( n6827 , n2991 , n551 );
xor ( n6828 , n6826 , n6827 );
and ( n6829 , n6427 , n6428 );
and ( n6830 , n6429 , n6432 );
or ( n6831 , n6829 , n6830 );
xor ( n6832 , n6828 , n6831 );
nor ( n6833 , n3464 , n665 );
xor ( n6834 , n6832 , n6833 );
and ( n6835 , n6433 , n6434 );
and ( n6836 , n6435 , n6438 );
or ( n6837 , n6835 , n6836 );
xor ( n6838 , n6834 , n6837 );
nor ( n6839 , n3863 , n797 );
xor ( n6840 , n6838 , n6839 );
and ( n6841 , n6439 , n6440 );
and ( n6842 , n6441 , n6444 );
or ( n6843 , n6841 , n6842 );
xor ( n6844 , n6840 , n6843 );
nor ( n6845 , n4260 , n954 );
xor ( n6846 , n6844 , n6845 );
and ( n6847 , n6445 , n6446 );
and ( n6848 , n6447 , n6450 );
or ( n6849 , n6847 , n6848 );
xor ( n6850 , n6846 , n6849 );
nor ( n6851 , n4659 , n1128 );
xor ( n6852 , n6850 , n6851 );
and ( n6853 , n6451 , n6452 );
and ( n6854 , n6453 , n6456 );
or ( n6855 , n6853 , n6854 );
xor ( n6856 , n6852 , n6855 );
nor ( n6857 , n5057 , n1320 );
xor ( n6858 , n6856 , n6857 );
and ( n6859 , n6457 , n6458 );
and ( n6860 , n6459 , n6462 );
or ( n6861 , n6859 , n6860 );
xor ( n6862 , n6858 , n6861 );
nor ( n6863 , n5453 , n1536 );
xor ( n6864 , n6862 , n6863 );
and ( n6865 , n6463 , n6464 );
and ( n6866 , n6465 , n6468 );
or ( n6867 , n6865 , n6866 );
xor ( n6868 , n6864 , n6867 );
nor ( n6869 , n5851 , n1773 );
xor ( n6870 , n6868 , n6869 );
and ( n6871 , n6469 , n6470 );
and ( n6872 , n6471 , n6474 );
or ( n6873 , n6871 , n6872 );
xor ( n6874 , n6870 , n6873 );
nor ( n6875 , n6249 , n2027 );
xor ( n6876 , n6874 , n6875 );
and ( n6877 , n6475 , n6476 );
and ( n6878 , n6477 , n6480 );
or ( n6879 , n6877 , n6878 );
xor ( n6880 , n6876 , n6879 );
nor ( n6881 , n6642 , n2302 );
xor ( n6882 , n6880 , n6881 );
and ( n6883 , n6481 , n6482 );
and ( n6884 , n6483 , n6486 );
or ( n6885 , n6883 , n6884 );
xor ( n6886 , n6882 , n6885 );
and ( n6887 , n6504 , n6508 );
and ( n6888 , n6508 , n6512 );
and ( n6889 , n6504 , n6512 );
or ( n6890 , n6887 , n6888 , n6889 );
and ( n6891 , n6500 , n6513 );
and ( n6892 , n6513 , n6628 );
and ( n6893 , n6500 , n6628 );
or ( n6894 , n6891 , n6892 , n6893 );
xor ( n6895 , n6890 , n6894 );
and ( n6896 , n6518 , n6544 );
and ( n6897 , n6544 , n6627 );
and ( n6898 , n6518 , n6627 );
or ( n6899 , n6896 , n6897 , n6898 );
and ( n6900 , n6532 , n6533 );
and ( n6901 , n6533 , n6535 );
and ( n6902 , n6532 , n6535 );
or ( n6903 , n6900 , n6901 , n6902 );
and ( n6904 , n6522 , n6526 );
and ( n6905 , n6526 , n6543 );
and ( n6906 , n6522 , n6543 );
or ( n6907 , n6904 , n6905 , n6906 );
xor ( n6908 , n6903 , n6907 );
not ( n6909 , n1516 );
and ( n6910 , n2406 , n1516 );
nor ( n6911 , n6909 , n6910 );
xor ( n6912 , n6908 , n6911 );
xor ( n6913 , n6899 , n6912 );
and ( n6914 , n6549 , n6564 );
and ( n6915 , n6564 , n6626 );
and ( n6916 , n6549 , n6626 );
or ( n6917 , n6914 , n6915 , n6916 );
and ( n6918 , n6531 , n6536 );
and ( n6919 , n6536 , n6542 );
and ( n6920 , n6531 , n6542 );
or ( n6921 , n6918 , n6919 , n6920 );
and ( n6922 , n6553 , n6557 );
and ( n6923 , n6557 , n6563 );
and ( n6924 , n6553 , n6563 );
or ( n6925 , n6922 , n6923 , n6924 );
xor ( n6926 , n6921 , n6925 );
and ( n6927 , n6538 , n6539 );
and ( n6928 , n6539 , n6541 );
and ( n6929 , n6538 , n6541 );
or ( n6930 , n6927 , n6928 , n6929 );
and ( n6931 , n1730 , n2138 );
and ( n6932 , n2001 , n1864 );
xor ( n6933 , n6931 , n6932 );
and ( n6934 , n2286 , n1753 );
xor ( n6935 , n6933 , n6934 );
xor ( n6936 , n6930 , n6935 );
and ( n6937 , n2581 , n1396 );
and ( n6938 , n2972 , n1302 );
xor ( n6939 , n6937 , n6938 );
and ( n6940 , n3445 , n1114 );
xor ( n6941 , n6939 , n6940 );
xor ( n6942 , n6936 , n6941 );
xor ( n6943 , n6926 , n6942 );
xor ( n6944 , n6917 , n6943 );
and ( n6945 , n6569 , n6574 );
and ( n6946 , n6574 , n6625 );
and ( n6947 , n6569 , n6625 );
or ( n6948 , n6945 , n6946 , n6947 );
and ( n6949 , n6559 , n6560 );
and ( n6950 , n6560 , n6562 );
and ( n6951 , n6559 , n6562 );
or ( n6952 , n6949 , n6950 , n6951 );
and ( n6953 , n6570 , n6571 );
and ( n6954 , n6571 , n6573 );
and ( n6955 , n6570 , n6573 );
or ( n6956 , n6953 , n6954 , n6955 );
xor ( n6957 , n6952 , n6956 );
and ( n6958 , n3844 , n852 );
and ( n6959 , n4241 , n714 );
xor ( n6960 , n6958 , n6959 );
and ( n6961 , n4640 , n651 );
xor ( n6962 , n6960 , n6961 );
xor ( n6963 , n6957 , n6962 );
xor ( n6964 , n6948 , n6963 );
and ( n6965 , n6576 , n6577 );
and ( n6966 , n6577 , n6624 );
and ( n6967 , n6576 , n6624 );
or ( n6968 , n6965 , n6966 , n6967 );
and ( n6969 , n5038 , n488 );
and ( n6970 , n5434 , n411 );
xor ( n6971 , n6969 , n6970 );
and ( n6972 , n5832 , n375 );
xor ( n6973 , n6971 , n6972 );
xor ( n6974 , n6968 , n6973 );
and ( n6975 , n6230 , n312 );
and ( n6976 , n6623 , n288 );
xor ( n6977 , n6975 , n6976 );
and ( n6978 , n6588 , n6589 );
and ( n6979 , n6589 , n6593 );
and ( n6980 , n6588 , n6593 );
or ( n6981 , n6978 , n6979 , n6980 );
and ( n6982 , n6594 , n6610 );
xor ( n6983 , n6981 , n6982 );
and ( n6984 , n6604 , n6605 );
and ( n6985 , n6605 , n6607 );
and ( n6986 , n6604 , n6607 );
or ( n6987 , n6984 , n6985 , n6986 );
and ( n6988 , n6598 , n6609 );
xor ( n6989 , n6987 , n6988 );
and ( n6990 , n2206 , n1685 );
not ( n6991 , n1685 );
nor ( n6992 , n6990 , n6991 );
xor ( n6993 , n6989 , n6992 );
and ( n6994 , n6599 , n6602 );
and ( n6995 , n6602 , n6608 );
and ( n6996 , n6599 , n6608 );
or ( n6997 , n6994 , n6995 , n6996 );
not ( n6998 , n1458 );
and ( n6999 , n2563 , n1458 );
nor ( n7000 , n6998 , n6999 );
and ( n7001 , n1713 , n2271 );
xor ( n7002 , n7000 , n7001 );
and ( n7003 , n1935 , n1975 );
xor ( n7004 , n7002 , n7003 );
xor ( n7005 , n6997 , n7004 );
xor ( n7006 , n6993 , n7005 );
xor ( n7007 , n6983 , n7006 );
and ( n7008 , n6582 , n6583 );
and ( n7009 , n6583 , n6611 );
and ( n7010 , n6582 , n6611 );
or ( n7011 , n7008 , n7009 , n7010 );
xor ( n7012 , n7007 , n7011 );
and ( n7013 , n6612 , n6616 );
and ( n7014 , n6617 , n6620 );
or ( n7015 , n7013 , n7014 );
xor ( n7016 , n7012 , n7015 );
buf ( n7017 , n7016 );
buf ( n7018 , n7017 );
and ( n7019 , n7018 , n279 );
xor ( n7020 , n6977 , n7019 );
xor ( n7021 , n6974 , n7020 );
xor ( n7022 , n6964 , n7021 );
xor ( n7023 , n6944 , n7022 );
xor ( n7024 , n6913 , n7023 );
xor ( n7025 , n6895 , n7024 );
and ( n7026 , n6491 , n6495 );
and ( n7027 , n6495 , n6629 );
and ( n7028 , n6491 , n6629 );
or ( n7029 , n7026 , n7027 , n7028 );
xor ( n7030 , n7025 , n7029 );
and ( n7031 , n6630 , n6634 );
and ( n7032 , n6635 , n6638 );
or ( n7033 , n7031 , n7032 );
xor ( n7034 , n7030 , n7033 );
buf ( n7035 , n7034 );
buf ( n7036 , n7035 );
not ( n7037 , n7036 );
nor ( n7038 , n7037 , n2598 );
xor ( n7039 , n6886 , n7038 );
and ( n7040 , n6487 , n6643 );
and ( n7041 , n6644 , n6647 );
or ( n7042 , n7040 , n7041 );
xor ( n7043 , n7039 , n7042 );
buf ( n7044 , n7043 );
buf ( n7045 , n7044 );
not ( n7046 , n7045 );
buf ( n7047 , n268 );
not ( n7048 , n7047 );
nor ( n7049 , n7046 , n7048 );
xor ( n7050 , n6800 , n7049 );
xor ( n7051 , n6659 , n6797 );
nor ( n7052 , n6651 , n7048 );
and ( n7053 , n7051 , n7052 );
xor ( n7054 , n7051 , n7052 );
xor ( n7055 , n6663 , n6795 );
nor ( n7056 , n6258 , n7048 );
and ( n7057 , n7055 , n7056 );
xor ( n7058 , n7055 , n7056 );
xor ( n7059 , n6667 , n6793 );
nor ( n7060 , n5860 , n7048 );
and ( n7061 , n7059 , n7060 );
xor ( n7062 , n7059 , n7060 );
xor ( n7063 , n6671 , n6791 );
nor ( n7064 , n5462 , n7048 );
and ( n7065 , n7063 , n7064 );
xor ( n7066 , n7063 , n7064 );
xor ( n7067 , n6675 , n6789 );
nor ( n7068 , n5066 , n7048 );
and ( n7069 , n7067 , n7068 );
xor ( n7070 , n7067 , n7068 );
xor ( n7071 , n6679 , n6787 );
nor ( n7072 , n4668 , n7048 );
and ( n7073 , n7071 , n7072 );
xor ( n7074 , n7071 , n7072 );
xor ( n7075 , n6683 , n6785 );
nor ( n7076 , n4269 , n7048 );
and ( n7077 , n7075 , n7076 );
xor ( n7078 , n7075 , n7076 );
xor ( n7079 , n6687 , n6783 );
nor ( n7080 , n3872 , n7048 );
and ( n7081 , n7079 , n7080 );
xor ( n7082 , n7079 , n7080 );
xor ( n7083 , n6691 , n6781 );
nor ( n7084 , n3473 , n7048 );
and ( n7085 , n7083 , n7084 );
xor ( n7086 , n7083 , n7084 );
xor ( n7087 , n6695 , n6779 );
nor ( n7088 , n3000 , n7048 );
and ( n7089 , n7087 , n7088 );
xor ( n7090 , n7087 , n7088 );
xor ( n7091 , n6699 , n6777 );
nor ( n7092 , n2688 , n7048 );
and ( n7093 , n7091 , n7092 );
xor ( n7094 , n7091 , n7092 );
xor ( n7095 , n6703 , n6775 );
nor ( n7096 , n3008 , n7048 );
and ( n7097 , n7095 , n7096 );
xor ( n7098 , n7095 , n7096 );
xor ( n7099 , n6707 , n6773 );
nor ( n7100 , n3017 , n7048 );
and ( n7101 , n7099 , n7100 );
xor ( n7102 , n7099 , n7100 );
xor ( n7103 , n6711 , n6771 );
nor ( n7104 , n3026 , n7048 );
and ( n7105 , n7103 , n7104 );
xor ( n7106 , n7103 , n7104 );
xor ( n7107 , n6715 , n6769 );
nor ( n7108 , n3035 , n7048 );
and ( n7109 , n7107 , n7108 );
xor ( n7110 , n7107 , n7108 );
xor ( n7111 , n6719 , n6767 );
nor ( n7112 , n3044 , n7048 );
and ( n7113 , n7111 , n7112 );
xor ( n7114 , n7111 , n7112 );
xor ( n7115 , n6723 , n6765 );
nor ( n7116 , n3053 , n7048 );
and ( n7117 , n7115 , n7116 );
xor ( n7118 , n7115 , n7116 );
xor ( n7119 , n6727 , n6763 );
nor ( n7120 , n3062 , n7048 );
and ( n7121 , n7119 , n7120 );
xor ( n7122 , n7119 , n7120 );
xor ( n7123 , n6731 , n6761 );
nor ( n7124 , n3071 , n7048 );
and ( n7125 , n7123 , n7124 );
xor ( n7126 , n7123 , n7124 );
xor ( n7127 , n6735 , n6759 );
nor ( n7128 , n3080 , n7048 );
and ( n7129 , n7127 , n7128 );
xor ( n7130 , n7127 , n7128 );
xor ( n7131 , n6739 , n6757 );
nor ( n7132 , n3089 , n7048 );
and ( n7133 , n7131 , n7132 );
xor ( n7134 , n7131 , n7132 );
xor ( n7135 , n6743 , n6755 );
nor ( n7136 , n3098 , n7048 );
and ( n7137 , n7135 , n7136 );
xor ( n7138 , n7135 , n7136 );
xor ( n7139 , n6748 , n6753 );
nor ( n7140 , n3107 , n7048 );
and ( n7141 , n7139 , n7140 );
xor ( n7142 , n7139 , n7140 );
xor ( n7143 , n6750 , n6751 );
buf ( n7144 , n7143 );
nor ( n7145 , n3116 , n7048 );
and ( n7146 , n7144 , n7145 );
xor ( n7147 , n7144 , n7145 );
nor ( n7148 , n3134 , n6653 );
buf ( n7149 , n7148 );
nor ( n7150 , n3125 , n7048 );
and ( n7151 , n7149 , n7150 );
buf ( n7152 , n7151 );
and ( n7153 , n7147 , n7152 );
or ( n7154 , n7146 , n7153 );
and ( n7155 , n7142 , n7154 );
or ( n7156 , n7141 , n7155 );
and ( n7157 , n7138 , n7156 );
or ( n7158 , n7137 , n7157 );
and ( n7159 , n7134 , n7158 );
or ( n7160 , n7133 , n7159 );
and ( n7161 , n7130 , n7160 );
or ( n7162 , n7129 , n7161 );
and ( n7163 , n7126 , n7162 );
or ( n7164 , n7125 , n7163 );
and ( n7165 , n7122 , n7164 );
or ( n7166 , n7121 , n7165 );
and ( n7167 , n7118 , n7166 );
or ( n7168 , n7117 , n7167 );
and ( n7169 , n7114 , n7168 );
or ( n7170 , n7113 , n7169 );
and ( n7171 , n7110 , n7170 );
or ( n7172 , n7109 , n7171 );
and ( n7173 , n7106 , n7172 );
or ( n7174 , n7105 , n7173 );
and ( n7175 , n7102 , n7174 );
or ( n7176 , n7101 , n7175 );
and ( n7177 , n7098 , n7176 );
or ( n7178 , n7097 , n7177 );
and ( n7179 , n7094 , n7178 );
or ( n7180 , n7093 , n7179 );
and ( n7181 , n7090 , n7180 );
or ( n7182 , n7089 , n7181 );
and ( n7183 , n7086 , n7182 );
or ( n7184 , n7085 , n7183 );
and ( n7185 , n7082 , n7184 );
or ( n7186 , n7081 , n7185 );
and ( n7187 , n7078 , n7186 );
or ( n7188 , n7077 , n7187 );
and ( n7189 , n7074 , n7188 );
or ( n7190 , n7073 , n7189 );
and ( n7191 , n7070 , n7190 );
or ( n7192 , n7069 , n7191 );
and ( n7193 , n7066 , n7192 );
or ( n7194 , n7065 , n7193 );
and ( n7195 , n7062 , n7194 );
or ( n7196 , n7061 , n7195 );
and ( n7197 , n7058 , n7196 );
or ( n7198 , n7057 , n7197 );
and ( n7199 , n7054 , n7198 );
or ( n7200 , n7053 , n7199 );
xor ( n7201 , n7050 , n7200 );
and ( n7202 , n285 , n1770 );
nor ( n7203 , n1771 , n7202 );
nor ( n7204 , n2025 , n305 );
xor ( n7205 , n7203 , n7204 );
and ( n7206 , n6802 , n6803 );
and ( n7207 , n6804 , n6807 );
or ( n7208 , n7206 , n7207 );
xor ( n7209 , n7205 , n7208 );
nor ( n7210 , n2300 , n336 );
xor ( n7211 , n7209 , n7210 );
and ( n7212 , n6808 , n6809 );
and ( n7213 , n6810 , n6813 );
or ( n7214 , n7212 , n7213 );
xor ( n7215 , n7211 , n7214 );
nor ( n7216 , n2596 , n386 );
xor ( n7217 , n7215 , n7216 );
and ( n7218 , n6814 , n6815 );
and ( n7219 , n6816 , n6819 );
or ( n7220 , n7218 , n7219 );
xor ( n7221 , n7217 , n7220 );
nor ( n7222 , n2991 , n458 );
xor ( n7223 , n7221 , n7222 );
and ( n7224 , n6820 , n6821 );
and ( n7225 , n6822 , n6825 );
or ( n7226 , n7224 , n7225 );
xor ( n7227 , n7223 , n7226 );
nor ( n7228 , n3464 , n551 );
xor ( n7229 , n7227 , n7228 );
and ( n7230 , n6826 , n6827 );
and ( n7231 , n6828 , n6831 );
or ( n7232 , n7230 , n7231 );
xor ( n7233 , n7229 , n7232 );
nor ( n7234 , n3863 , n665 );
xor ( n7235 , n7233 , n7234 );
and ( n7236 , n6832 , n6833 );
and ( n7237 , n6834 , n6837 );
or ( n7238 , n7236 , n7237 );
xor ( n7239 , n7235 , n7238 );
nor ( n7240 , n4260 , n797 );
xor ( n7241 , n7239 , n7240 );
and ( n7242 , n6838 , n6839 );
and ( n7243 , n6840 , n6843 );
or ( n7244 , n7242 , n7243 );
xor ( n7245 , n7241 , n7244 );
nor ( n7246 , n4659 , n954 );
xor ( n7247 , n7245 , n7246 );
and ( n7248 , n6844 , n6845 );
and ( n7249 , n6846 , n6849 );
or ( n7250 , n7248 , n7249 );
xor ( n7251 , n7247 , n7250 );
nor ( n7252 , n5057 , n1128 );
xor ( n7253 , n7251 , n7252 );
and ( n7254 , n6850 , n6851 );
and ( n7255 , n6852 , n6855 );
or ( n7256 , n7254 , n7255 );
xor ( n7257 , n7253 , n7256 );
nor ( n7258 , n5453 , n1320 );
xor ( n7259 , n7257 , n7258 );
and ( n7260 , n6856 , n6857 );
and ( n7261 , n6858 , n6861 );
or ( n7262 , n7260 , n7261 );
xor ( n7263 , n7259 , n7262 );
nor ( n7264 , n5851 , n1536 );
xor ( n7265 , n7263 , n7264 );
and ( n7266 , n6862 , n6863 );
and ( n7267 , n6864 , n6867 );
or ( n7268 , n7266 , n7267 );
xor ( n7269 , n7265 , n7268 );
nor ( n7270 , n6249 , n1773 );
xor ( n7271 , n7269 , n7270 );
and ( n7272 , n6868 , n6869 );
and ( n7273 , n6870 , n6873 );
or ( n7274 , n7272 , n7273 );
xor ( n7275 , n7271 , n7274 );
nor ( n7276 , n6642 , n2027 );
xor ( n7277 , n7275 , n7276 );
and ( n7278 , n6874 , n6875 );
and ( n7279 , n6876 , n6879 );
or ( n7280 , n7278 , n7279 );
xor ( n7281 , n7277 , n7280 );
nor ( n7282 , n7037 , n2302 );
xor ( n7283 , n7281 , n7282 );
and ( n7284 , n6880 , n6881 );
and ( n7285 , n6882 , n6885 );
or ( n7286 , n7284 , n7285 );
xor ( n7287 , n7283 , n7286 );
and ( n7288 , n6903 , n6907 );
and ( n7289 , n6907 , n6911 );
and ( n7290 , n6903 , n6911 );
or ( n7291 , n7288 , n7289 , n7290 );
and ( n7292 , n6899 , n6912 );
and ( n7293 , n6912 , n7023 );
and ( n7294 , n6899 , n7023 );
or ( n7295 , n7292 , n7293 , n7294 );
xor ( n7296 , n7291 , n7295 );
and ( n7297 , n6917 , n6943 );
and ( n7298 , n6943 , n7022 );
and ( n7299 , n6917 , n7022 );
or ( n7300 , n7297 , n7298 , n7299 );
and ( n7301 , n6931 , n6932 );
and ( n7302 , n6932 , n6934 );
and ( n7303 , n6931 , n6934 );
or ( n7304 , n7301 , n7302 , n7303 );
and ( n7305 , n6921 , n6925 );
and ( n7306 , n6925 , n6942 );
and ( n7307 , n6921 , n6942 );
or ( n7308 , n7305 , n7306 , n7307 );
xor ( n7309 , n7304 , n7308 );
not ( n7310 , n1730 );
and ( n7311 , n2406 , n1730 );
nor ( n7312 , n7310 , n7311 );
xor ( n7313 , n7309 , n7312 );
xor ( n7314 , n7300 , n7313 );
and ( n7315 , n6948 , n6963 );
and ( n7316 , n6963 , n7021 );
and ( n7317 , n6948 , n7021 );
or ( n7318 , n7315 , n7316 , n7317 );
and ( n7319 , n6930 , n6935 );
and ( n7320 , n6935 , n6941 );
and ( n7321 , n6930 , n6941 );
or ( n7322 , n7319 , n7320 , n7321 );
and ( n7323 , n6952 , n6956 );
and ( n7324 , n6956 , n6962 );
and ( n7325 , n6952 , n6962 );
or ( n7326 , n7323 , n7324 , n7325 );
xor ( n7327 , n7322 , n7326 );
and ( n7328 , n6937 , n6938 );
and ( n7329 , n6938 , n6940 );
and ( n7330 , n6937 , n6940 );
or ( n7331 , n7328 , n7329 , n7330 );
and ( n7332 , n2001 , n2138 );
and ( n7333 , n2286 , n1864 );
xor ( n7334 , n7332 , n7333 );
and ( n7335 , n2581 , n1753 );
xor ( n7336 , n7334 , n7335 );
xor ( n7337 , n7331 , n7336 );
and ( n7338 , n2972 , n1396 );
and ( n7339 , n3445 , n1302 );
xor ( n7340 , n7338 , n7339 );
and ( n7341 , n3844 , n1114 );
xor ( n7342 , n7340 , n7341 );
xor ( n7343 , n7337 , n7342 );
xor ( n7344 , n7327 , n7343 );
xor ( n7345 , n7318 , n7344 );
and ( n7346 , n6968 , n6973 );
and ( n7347 , n6973 , n7020 );
and ( n7348 , n6968 , n7020 );
or ( n7349 , n7346 , n7347 , n7348 );
and ( n7350 , n6958 , n6959 );
and ( n7351 , n6959 , n6961 );
and ( n7352 , n6958 , n6961 );
or ( n7353 , n7350 , n7351 , n7352 );
and ( n7354 , n6969 , n6970 );
and ( n7355 , n6970 , n6972 );
and ( n7356 , n6969 , n6972 );
or ( n7357 , n7354 , n7355 , n7356 );
xor ( n7358 , n7353 , n7357 );
and ( n7359 , n4241 , n852 );
and ( n7360 , n4640 , n714 );
xor ( n7361 , n7359 , n7360 );
and ( n7362 , n5038 , n651 );
xor ( n7363 , n7361 , n7362 );
xor ( n7364 , n7358 , n7363 );
xor ( n7365 , n7349 , n7364 );
and ( n7366 , n6975 , n6976 );
and ( n7367 , n6976 , n7019 );
and ( n7368 , n6975 , n7019 );
or ( n7369 , n7366 , n7367 , n7368 );
and ( n7370 , n5434 , n488 );
and ( n7371 , n5832 , n411 );
xor ( n7372 , n7370 , n7371 );
and ( n7373 , n6230 , n375 );
xor ( n7374 , n7372 , n7373 );
xor ( n7375 , n7369 , n7374 );
and ( n7376 , n6623 , n312 );
and ( n7377 , n7018 , n288 );
xor ( n7378 , n7376 , n7377 );
and ( n7379 , n6987 , n6988 );
and ( n7380 , n6988 , n6992 );
and ( n7381 , n6987 , n6992 );
or ( n7382 , n7379 , n7380 , n7381 );
and ( n7383 , n6993 , n7005 );
xor ( n7384 , n7382 , n7383 );
and ( n7385 , n7000 , n7001 );
and ( n7386 , n7001 , n7003 );
and ( n7387 , n7000 , n7003 );
or ( n7388 , n7385 , n7386 , n7387 );
and ( n7389 , n6997 , n7004 );
xor ( n7390 , n7388 , n7389 );
and ( n7391 , n2206 , n1975 );
not ( n7392 , n1975 );
nor ( n7393 , n7391 , n7392 );
xor ( n7394 , n7390 , n7393 );
not ( n7395 , n1713 );
and ( n7396 , n2563 , n1713 );
nor ( n7397 , n7395 , n7396 );
and ( n7398 , n1935 , n2271 );
xor ( n7399 , n7397 , n7398 );
xor ( n7400 , n7394 , n7399 );
xor ( n7401 , n7384 , n7400 );
and ( n7402 , n6981 , n6982 );
and ( n7403 , n6982 , n7006 );
and ( n7404 , n6981 , n7006 );
or ( n7405 , n7402 , n7403 , n7404 );
xor ( n7406 , n7401 , n7405 );
and ( n7407 , n7007 , n7011 );
and ( n7408 , n7012 , n7015 );
or ( n7409 , n7407 , n7408 );
xor ( n7410 , n7406 , n7409 );
buf ( n7411 , n7410 );
buf ( n7412 , n7411 );
and ( n7413 , n7412 , n279 );
xor ( n7414 , n7378 , n7413 );
xor ( n7415 , n7375 , n7414 );
xor ( n7416 , n7365 , n7415 );
xor ( n7417 , n7345 , n7416 );
xor ( n7418 , n7314 , n7417 );
xor ( n7419 , n7296 , n7418 );
and ( n7420 , n6890 , n6894 );
and ( n7421 , n6894 , n7024 );
and ( n7422 , n6890 , n7024 );
or ( n7423 , n7420 , n7421 , n7422 );
xor ( n7424 , n7419 , n7423 );
and ( n7425 , n7025 , n7029 );
and ( n7426 , n7030 , n7033 );
or ( n7427 , n7425 , n7426 );
xor ( n7428 , n7424 , n7427 );
buf ( n7429 , n7428 );
buf ( n7430 , n7429 );
not ( n7431 , n7430 );
nor ( n7432 , n7431 , n2598 );
xor ( n7433 , n7287 , n7432 );
and ( n7434 , n6886 , n7038 );
and ( n7435 , n7039 , n7042 );
or ( n7436 , n7434 , n7435 );
xor ( n7437 , n7433 , n7436 );
buf ( n7438 , n7437 );
buf ( n7439 , n7438 );
not ( n7440 , n7439 );
buf ( n7441 , n269 );
not ( n7442 , n7441 );
nor ( n7443 , n7440 , n7442 );
xor ( n7444 , n7201 , n7443 );
xor ( n7445 , n7054 , n7198 );
nor ( n7446 , n7046 , n7442 );
and ( n7447 , n7445 , n7446 );
xor ( n7448 , n7445 , n7446 );
xor ( n7449 , n7058 , n7196 );
nor ( n7450 , n6651 , n7442 );
and ( n7451 , n7449 , n7450 );
xor ( n7452 , n7449 , n7450 );
xor ( n7453 , n7062 , n7194 );
nor ( n7454 , n6258 , n7442 );
and ( n7455 , n7453 , n7454 );
xor ( n7456 , n7453 , n7454 );
xor ( n7457 , n7066 , n7192 );
nor ( n7458 , n5860 , n7442 );
and ( n7459 , n7457 , n7458 );
xor ( n7460 , n7457 , n7458 );
xor ( n7461 , n7070 , n7190 );
nor ( n7462 , n5462 , n7442 );
and ( n7463 , n7461 , n7462 );
xor ( n7464 , n7461 , n7462 );
xor ( n7465 , n7074 , n7188 );
nor ( n7466 , n5066 , n7442 );
and ( n7467 , n7465 , n7466 );
xor ( n7468 , n7465 , n7466 );
xor ( n7469 , n7078 , n7186 );
nor ( n7470 , n4668 , n7442 );
and ( n7471 , n7469 , n7470 );
xor ( n7472 , n7469 , n7470 );
xor ( n7473 , n7082 , n7184 );
nor ( n7474 , n4269 , n7442 );
and ( n7475 , n7473 , n7474 );
xor ( n7476 , n7473 , n7474 );
xor ( n7477 , n7086 , n7182 );
nor ( n7478 , n3872 , n7442 );
and ( n7479 , n7477 , n7478 );
xor ( n7480 , n7477 , n7478 );
xor ( n7481 , n7090 , n7180 );
nor ( n7482 , n3473 , n7442 );
and ( n7483 , n7481 , n7482 );
xor ( n7484 , n7481 , n7482 );
xor ( n7485 , n7094 , n7178 );
nor ( n7486 , n3000 , n7442 );
and ( n7487 , n7485 , n7486 );
xor ( n7488 , n7485 , n7486 );
xor ( n7489 , n7098 , n7176 );
nor ( n7490 , n2688 , n7442 );
and ( n7491 , n7489 , n7490 );
xor ( n7492 , n7489 , n7490 );
xor ( n7493 , n7102 , n7174 );
nor ( n7494 , n3008 , n7442 );
and ( n7495 , n7493 , n7494 );
xor ( n7496 , n7493 , n7494 );
xor ( n7497 , n7106 , n7172 );
nor ( n7498 , n3017 , n7442 );
and ( n7499 , n7497 , n7498 );
xor ( n7500 , n7497 , n7498 );
xor ( n7501 , n7110 , n7170 );
nor ( n7502 , n3026 , n7442 );
and ( n7503 , n7501 , n7502 );
xor ( n7504 , n7501 , n7502 );
xor ( n7505 , n7114 , n7168 );
nor ( n7506 , n3035 , n7442 );
and ( n7507 , n7505 , n7506 );
xor ( n7508 , n7505 , n7506 );
xor ( n7509 , n7118 , n7166 );
nor ( n7510 , n3044 , n7442 );
and ( n7511 , n7509 , n7510 );
xor ( n7512 , n7509 , n7510 );
xor ( n7513 , n7122 , n7164 );
nor ( n7514 , n3053 , n7442 );
and ( n7515 , n7513 , n7514 );
xor ( n7516 , n7513 , n7514 );
xor ( n7517 , n7126 , n7162 );
nor ( n7518 , n3062 , n7442 );
and ( n7519 , n7517 , n7518 );
xor ( n7520 , n7517 , n7518 );
xor ( n7521 , n7130 , n7160 );
nor ( n7522 , n3071 , n7442 );
and ( n7523 , n7521 , n7522 );
xor ( n7524 , n7521 , n7522 );
xor ( n7525 , n7134 , n7158 );
nor ( n7526 , n3080 , n7442 );
and ( n7527 , n7525 , n7526 );
xor ( n7528 , n7525 , n7526 );
xor ( n7529 , n7138 , n7156 );
nor ( n7530 , n3089 , n7442 );
and ( n7531 , n7529 , n7530 );
xor ( n7532 , n7529 , n7530 );
xor ( n7533 , n7142 , n7154 );
nor ( n7534 , n3098 , n7442 );
and ( n7535 , n7533 , n7534 );
xor ( n7536 , n7533 , n7534 );
xor ( n7537 , n7147 , n7152 );
nor ( n7538 , n3107 , n7442 );
and ( n7539 , n7537 , n7538 );
xor ( n7540 , n7537 , n7538 );
xor ( n7541 , n7149 , n7150 );
buf ( n7542 , n7541 );
nor ( n7543 , n3116 , n7442 );
and ( n7544 , n7542 , n7543 );
xor ( n7545 , n7542 , n7543 );
nor ( n7546 , n3134 , n7048 );
buf ( n7547 , n7546 );
nor ( n7548 , n3125 , n7442 );
and ( n7549 , n7547 , n7548 );
buf ( n7550 , n7549 );
and ( n7551 , n7545 , n7550 );
or ( n7552 , n7544 , n7551 );
and ( n7553 , n7540 , n7552 );
or ( n7554 , n7539 , n7553 );
and ( n7555 , n7536 , n7554 );
or ( n7556 , n7535 , n7555 );
and ( n7557 , n7532 , n7556 );
or ( n7558 , n7531 , n7557 );
and ( n7559 , n7528 , n7558 );
or ( n7560 , n7527 , n7559 );
and ( n7561 , n7524 , n7560 );
or ( n7562 , n7523 , n7561 );
and ( n7563 , n7520 , n7562 );
or ( n7564 , n7519 , n7563 );
and ( n7565 , n7516 , n7564 );
or ( n7566 , n7515 , n7565 );
and ( n7567 , n7512 , n7566 );
or ( n7568 , n7511 , n7567 );
and ( n7569 , n7508 , n7568 );
or ( n7570 , n7507 , n7569 );
and ( n7571 , n7504 , n7570 );
or ( n7572 , n7503 , n7571 );
and ( n7573 , n7500 , n7572 );
or ( n7574 , n7499 , n7573 );
and ( n7575 , n7496 , n7574 );
or ( n7576 , n7495 , n7575 );
and ( n7577 , n7492 , n7576 );
or ( n7578 , n7491 , n7577 );
and ( n7579 , n7488 , n7578 );
or ( n7580 , n7487 , n7579 );
and ( n7581 , n7484 , n7580 );
or ( n7582 , n7483 , n7581 );
and ( n7583 , n7480 , n7582 );
or ( n7584 , n7479 , n7583 );
and ( n7585 , n7476 , n7584 );
or ( n7586 , n7475 , n7585 );
and ( n7587 , n7472 , n7586 );
or ( n7588 , n7471 , n7587 );
and ( n7589 , n7468 , n7588 );
or ( n7590 , n7467 , n7589 );
and ( n7591 , n7464 , n7590 );
or ( n7592 , n7463 , n7591 );
and ( n7593 , n7460 , n7592 );
or ( n7594 , n7459 , n7593 );
and ( n7595 , n7456 , n7594 );
or ( n7596 , n7455 , n7595 );
and ( n7597 , n7452 , n7596 );
or ( n7598 , n7451 , n7597 );
and ( n7599 , n7448 , n7598 );
or ( n7600 , n7447 , n7599 );
xor ( n7601 , n7444 , n7600 );
and ( n7602 , n285 , n2024 );
nor ( n7603 , n2025 , n7602 );
nor ( n7604 , n2300 , n305 );
xor ( n7605 , n7603 , n7604 );
and ( n7606 , n7203 , n7204 );
and ( n7607 , n7205 , n7208 );
or ( n7608 , n7606 , n7607 );
xor ( n7609 , n7605 , n7608 );
nor ( n7610 , n2596 , n336 );
xor ( n7611 , n7609 , n7610 );
and ( n7612 , n7209 , n7210 );
and ( n7613 , n7211 , n7214 );
or ( n7614 , n7612 , n7613 );
xor ( n7615 , n7611 , n7614 );
nor ( n7616 , n2991 , n386 );
xor ( n7617 , n7615 , n7616 );
and ( n7618 , n7215 , n7216 );
and ( n7619 , n7217 , n7220 );
or ( n7620 , n7618 , n7619 );
xor ( n7621 , n7617 , n7620 );
nor ( n7622 , n3464 , n458 );
xor ( n7623 , n7621 , n7622 );
and ( n7624 , n7221 , n7222 );
and ( n7625 , n7223 , n7226 );
or ( n7626 , n7624 , n7625 );
xor ( n7627 , n7623 , n7626 );
nor ( n7628 , n3863 , n551 );
xor ( n7629 , n7627 , n7628 );
and ( n7630 , n7227 , n7228 );
and ( n7631 , n7229 , n7232 );
or ( n7632 , n7630 , n7631 );
xor ( n7633 , n7629 , n7632 );
nor ( n7634 , n4260 , n665 );
xor ( n7635 , n7633 , n7634 );
and ( n7636 , n7233 , n7234 );
and ( n7637 , n7235 , n7238 );
or ( n7638 , n7636 , n7637 );
xor ( n7639 , n7635 , n7638 );
nor ( n7640 , n4659 , n797 );
xor ( n7641 , n7639 , n7640 );
and ( n7642 , n7239 , n7240 );
and ( n7643 , n7241 , n7244 );
or ( n7644 , n7642 , n7643 );
xor ( n7645 , n7641 , n7644 );
nor ( n7646 , n5057 , n954 );
xor ( n7647 , n7645 , n7646 );
and ( n7648 , n7245 , n7246 );
and ( n7649 , n7247 , n7250 );
or ( n7650 , n7648 , n7649 );
xor ( n7651 , n7647 , n7650 );
nor ( n7652 , n5453 , n1128 );
xor ( n7653 , n7651 , n7652 );
and ( n7654 , n7251 , n7252 );
and ( n7655 , n7253 , n7256 );
or ( n7656 , n7654 , n7655 );
xor ( n7657 , n7653 , n7656 );
nor ( n7658 , n5851 , n1320 );
xor ( n7659 , n7657 , n7658 );
and ( n7660 , n7257 , n7258 );
and ( n7661 , n7259 , n7262 );
or ( n7662 , n7660 , n7661 );
xor ( n7663 , n7659 , n7662 );
nor ( n7664 , n6249 , n1536 );
xor ( n7665 , n7663 , n7664 );
and ( n7666 , n7263 , n7264 );
and ( n7667 , n7265 , n7268 );
or ( n7668 , n7666 , n7667 );
xor ( n7669 , n7665 , n7668 );
nor ( n7670 , n6642 , n1773 );
xor ( n7671 , n7669 , n7670 );
and ( n7672 , n7269 , n7270 );
and ( n7673 , n7271 , n7274 );
or ( n7674 , n7672 , n7673 );
xor ( n7675 , n7671 , n7674 );
nor ( n7676 , n7037 , n2027 );
xor ( n7677 , n7675 , n7676 );
and ( n7678 , n7275 , n7276 );
and ( n7679 , n7277 , n7280 );
or ( n7680 , n7678 , n7679 );
xor ( n7681 , n7677 , n7680 );
nor ( n7682 , n7431 , n2302 );
xor ( n7683 , n7681 , n7682 );
and ( n7684 , n7281 , n7282 );
and ( n7685 , n7283 , n7286 );
or ( n7686 , n7684 , n7685 );
xor ( n7687 , n7683 , n7686 );
and ( n7688 , n7304 , n7308 );
and ( n7689 , n7308 , n7312 );
and ( n7690 , n7304 , n7312 );
or ( n7691 , n7688 , n7689 , n7690 );
and ( n7692 , n7300 , n7313 );
and ( n7693 , n7313 , n7417 );
and ( n7694 , n7300 , n7417 );
or ( n7695 , n7692 , n7693 , n7694 );
xor ( n7696 , n7691 , n7695 );
and ( n7697 , n7318 , n7344 );
and ( n7698 , n7344 , n7416 );
and ( n7699 , n7318 , n7416 );
or ( n7700 , n7697 , n7698 , n7699 );
and ( n7701 , n7332 , n7333 );
and ( n7702 , n7333 , n7335 );
and ( n7703 , n7332 , n7335 );
or ( n7704 , n7701 , n7702 , n7703 );
and ( n7705 , n7322 , n7326 );
and ( n7706 , n7326 , n7343 );
and ( n7707 , n7322 , n7343 );
or ( n7708 , n7705 , n7706 , n7707 );
xor ( n7709 , n7704 , n7708 );
not ( n7710 , n2001 );
and ( n7711 , n2406 , n2001 );
nor ( n7712 , n7710 , n7711 );
xor ( n7713 , n7709 , n7712 );
xor ( n7714 , n7700 , n7713 );
and ( n7715 , n7349 , n7364 );
and ( n7716 , n7364 , n7415 );
and ( n7717 , n7349 , n7415 );
or ( n7718 , n7715 , n7716 , n7717 );
and ( n7719 , n7331 , n7336 );
and ( n7720 , n7336 , n7342 );
and ( n7721 , n7331 , n7342 );
or ( n7722 , n7719 , n7720 , n7721 );
and ( n7723 , n7353 , n7357 );
and ( n7724 , n7357 , n7363 );
and ( n7725 , n7353 , n7363 );
or ( n7726 , n7723 , n7724 , n7725 );
xor ( n7727 , n7722 , n7726 );
and ( n7728 , n7338 , n7339 );
and ( n7729 , n7339 , n7341 );
and ( n7730 , n7338 , n7341 );
or ( n7731 , n7728 , n7729 , n7730 );
and ( n7732 , n2286 , n2138 );
and ( n7733 , n2581 , n1864 );
xor ( n7734 , n7732 , n7733 );
and ( n7735 , n2972 , n1753 );
xor ( n7736 , n7734 , n7735 );
xor ( n7737 , n7731 , n7736 );
and ( n7738 , n3445 , n1396 );
and ( n7739 , n3844 , n1302 );
xor ( n7740 , n7738 , n7739 );
and ( n7741 , n4241 , n1114 );
xor ( n7742 , n7740 , n7741 );
xor ( n7743 , n7737 , n7742 );
xor ( n7744 , n7727 , n7743 );
xor ( n7745 , n7718 , n7744 );
and ( n7746 , n7369 , n7374 );
and ( n7747 , n7374 , n7414 );
and ( n7748 , n7369 , n7414 );
or ( n7749 , n7746 , n7747 , n7748 );
and ( n7750 , n7359 , n7360 );
and ( n7751 , n7360 , n7362 );
and ( n7752 , n7359 , n7362 );
or ( n7753 , n7750 , n7751 , n7752 );
and ( n7754 , n7370 , n7371 );
and ( n7755 , n7371 , n7373 );
and ( n7756 , n7370 , n7373 );
or ( n7757 , n7754 , n7755 , n7756 );
xor ( n7758 , n7753 , n7757 );
and ( n7759 , n4640 , n852 );
and ( n7760 , n5038 , n714 );
xor ( n7761 , n7759 , n7760 );
and ( n7762 , n5434 , n651 );
xor ( n7763 , n7761 , n7762 );
xor ( n7764 , n7758 , n7763 );
xor ( n7765 , n7749 , n7764 );
and ( n7766 , n7376 , n7377 );
and ( n7767 , n7377 , n7413 );
and ( n7768 , n7376 , n7413 );
or ( n7769 , n7766 , n7767 , n7768 );
and ( n7770 , n5832 , n488 );
and ( n7771 , n6230 , n411 );
xor ( n7772 , n7770 , n7771 );
and ( n7773 , n6623 , n375 );
xor ( n7774 , n7772 , n7773 );
xor ( n7775 , n7769 , n7774 );
and ( n7776 , n7018 , n312 );
and ( n7777 , n7412 , n288 );
xor ( n7778 , n7776 , n7777 );
and ( n7779 , n7388 , n7389 );
and ( n7780 , n7389 , n7393 );
and ( n7781 , n7388 , n7393 );
or ( n7782 , n7779 , n7780 , n7781 );
and ( n7783 , n7394 , n7399 );
xor ( n7784 , n7782 , n7783 );
not ( n7785 , n1935 );
and ( n7786 , n2563 , n1935 );
nor ( n7787 , n7785 , n7786 );
and ( n7788 , n7397 , n7398 );
and ( n7789 , n2206 , n2271 );
not ( n7790 , n2271 );
nor ( n7791 , n7789 , n7790 );
xor ( n7792 , n7788 , n7791 );
xor ( n7793 , n7787 , n7792 );
xor ( n7794 , n7784 , n7793 );
and ( n7795 , n7382 , n7383 );
and ( n7796 , n7383 , n7400 );
and ( n7797 , n7382 , n7400 );
or ( n7798 , n7795 , n7796 , n7797 );
xor ( n7799 , n7794 , n7798 );
and ( n7800 , n7401 , n7405 );
and ( n7801 , n7406 , n7409 );
or ( n7802 , n7800 , n7801 );
xor ( n7803 , n7799 , n7802 );
buf ( n7804 , n7803 );
buf ( n7805 , n7804 );
and ( n7806 , n7805 , n279 );
xor ( n7807 , n7778 , n7806 );
xor ( n7808 , n7775 , n7807 );
xor ( n7809 , n7765 , n7808 );
xor ( n7810 , n7745 , n7809 );
xor ( n7811 , n7714 , n7810 );
xor ( n7812 , n7696 , n7811 );
and ( n7813 , n7291 , n7295 );
and ( n7814 , n7295 , n7418 );
and ( n7815 , n7291 , n7418 );
or ( n7816 , n7813 , n7814 , n7815 );
xor ( n7817 , n7812 , n7816 );
and ( n7818 , n7419 , n7423 );
and ( n7819 , n7424 , n7427 );
or ( n7820 , n7818 , n7819 );
xor ( n7821 , n7817 , n7820 );
buf ( n7822 , n7821 );
buf ( n7823 , n7822 );
not ( n7824 , n7823 );
nor ( n7825 , n7824 , n2598 );
xor ( n7826 , n7687 , n7825 );
and ( n7827 , n7287 , n7432 );
and ( n7828 , n7433 , n7436 );
or ( n7829 , n7827 , n7828 );
xor ( n7830 , n7826 , n7829 );
buf ( n7831 , n7830 );
buf ( n7832 , n7831 );
not ( n7833 , n7832 );
buf ( n7834 , n270 );
not ( n7835 , n7834 );
nor ( n7836 , n7833 , n7835 );
xor ( n7837 , n7601 , n7836 );
xor ( n7838 , n7448 , n7598 );
nor ( n7839 , n7440 , n7835 );
and ( n7840 , n7838 , n7839 );
xor ( n7841 , n7838 , n7839 );
xor ( n7842 , n7452 , n7596 );
nor ( n7843 , n7046 , n7835 );
and ( n7844 , n7842 , n7843 );
xor ( n7845 , n7842 , n7843 );
xor ( n7846 , n7456 , n7594 );
nor ( n7847 , n6651 , n7835 );
and ( n7848 , n7846 , n7847 );
xor ( n7849 , n7846 , n7847 );
xor ( n7850 , n7460 , n7592 );
nor ( n7851 , n6258 , n7835 );
and ( n7852 , n7850 , n7851 );
xor ( n7853 , n7850 , n7851 );
xor ( n7854 , n7464 , n7590 );
nor ( n7855 , n5860 , n7835 );
and ( n7856 , n7854 , n7855 );
xor ( n7857 , n7854 , n7855 );
xor ( n7858 , n7468 , n7588 );
nor ( n7859 , n5462 , n7835 );
and ( n7860 , n7858 , n7859 );
xor ( n7861 , n7858 , n7859 );
xor ( n7862 , n7472 , n7586 );
nor ( n7863 , n5066 , n7835 );
and ( n7864 , n7862 , n7863 );
xor ( n7865 , n7862 , n7863 );
xor ( n7866 , n7476 , n7584 );
nor ( n7867 , n4668 , n7835 );
and ( n7868 , n7866 , n7867 );
xor ( n7869 , n7866 , n7867 );
xor ( n7870 , n7480 , n7582 );
nor ( n7871 , n4269 , n7835 );
and ( n7872 , n7870 , n7871 );
xor ( n7873 , n7870 , n7871 );
xor ( n7874 , n7484 , n7580 );
nor ( n7875 , n3872 , n7835 );
and ( n7876 , n7874 , n7875 );
xor ( n7877 , n7874 , n7875 );
xor ( n7878 , n7488 , n7578 );
nor ( n7879 , n3473 , n7835 );
and ( n7880 , n7878 , n7879 );
xor ( n7881 , n7878 , n7879 );
xor ( n7882 , n7492 , n7576 );
nor ( n7883 , n3000 , n7835 );
and ( n7884 , n7882 , n7883 );
xor ( n7885 , n7882 , n7883 );
xor ( n7886 , n7496 , n7574 );
nor ( n7887 , n2688 , n7835 );
and ( n7888 , n7886 , n7887 );
xor ( n7889 , n7886 , n7887 );
xor ( n7890 , n7500 , n7572 );
nor ( n7891 , n3008 , n7835 );
and ( n7892 , n7890 , n7891 );
xor ( n7893 , n7890 , n7891 );
xor ( n7894 , n7504 , n7570 );
nor ( n7895 , n3017 , n7835 );
and ( n7896 , n7894 , n7895 );
xor ( n7897 , n7894 , n7895 );
xor ( n7898 , n7508 , n7568 );
nor ( n7899 , n3026 , n7835 );
and ( n7900 , n7898 , n7899 );
xor ( n7901 , n7898 , n7899 );
xor ( n7902 , n7512 , n7566 );
nor ( n7903 , n3035 , n7835 );
and ( n7904 , n7902 , n7903 );
xor ( n7905 , n7902 , n7903 );
xor ( n7906 , n7516 , n7564 );
nor ( n7907 , n3044 , n7835 );
and ( n7908 , n7906 , n7907 );
xor ( n7909 , n7906 , n7907 );
xor ( n7910 , n7520 , n7562 );
nor ( n7911 , n3053 , n7835 );
and ( n7912 , n7910 , n7911 );
xor ( n7913 , n7910 , n7911 );
xor ( n7914 , n7524 , n7560 );
nor ( n7915 , n3062 , n7835 );
and ( n7916 , n7914 , n7915 );
xor ( n7917 , n7914 , n7915 );
xor ( n7918 , n7528 , n7558 );
nor ( n7919 , n3071 , n7835 );
and ( n7920 , n7918 , n7919 );
xor ( n7921 , n7918 , n7919 );
xor ( n7922 , n7532 , n7556 );
nor ( n7923 , n3080 , n7835 );
and ( n7924 , n7922 , n7923 );
xor ( n7925 , n7922 , n7923 );
xor ( n7926 , n7536 , n7554 );
nor ( n7927 , n3089 , n7835 );
and ( n7928 , n7926 , n7927 );
xor ( n7929 , n7926 , n7927 );
xor ( n7930 , n7540 , n7552 );
nor ( n7931 , n3098 , n7835 );
and ( n7932 , n7930 , n7931 );
xor ( n7933 , n7930 , n7931 );
xor ( n7934 , n7545 , n7550 );
nor ( n7935 , n3107 , n7835 );
and ( n7936 , n7934 , n7935 );
xor ( n7937 , n7934 , n7935 );
xor ( n7938 , n7547 , n7548 );
buf ( n7939 , n7938 );
nor ( n7940 , n3116 , n7835 );
and ( n7941 , n7939 , n7940 );
xor ( n7942 , n7939 , n7940 );
nor ( n7943 , n3134 , n7442 );
buf ( n7944 , n7943 );
nor ( n7945 , n3125 , n7835 );
and ( n7946 , n7944 , n7945 );
buf ( n7947 , n7946 );
and ( n7948 , n7942 , n7947 );
or ( n7949 , n7941 , n7948 );
and ( n7950 , n7937 , n7949 );
or ( n7951 , n7936 , n7950 );
and ( n7952 , n7933 , n7951 );
or ( n7953 , n7932 , n7952 );
and ( n7954 , n7929 , n7953 );
or ( n7955 , n7928 , n7954 );
and ( n7956 , n7925 , n7955 );
or ( n7957 , n7924 , n7956 );
and ( n7958 , n7921 , n7957 );
or ( n7959 , n7920 , n7958 );
and ( n7960 , n7917 , n7959 );
or ( n7961 , n7916 , n7960 );
and ( n7962 , n7913 , n7961 );
or ( n7963 , n7912 , n7962 );
and ( n7964 , n7909 , n7963 );
or ( n7965 , n7908 , n7964 );
and ( n7966 , n7905 , n7965 );
or ( n7967 , n7904 , n7966 );
and ( n7968 , n7901 , n7967 );
or ( n7969 , n7900 , n7968 );
and ( n7970 , n7897 , n7969 );
or ( n7971 , n7896 , n7970 );
and ( n7972 , n7893 , n7971 );
or ( n7973 , n7892 , n7972 );
and ( n7974 , n7889 , n7973 );
or ( n7975 , n7888 , n7974 );
and ( n7976 , n7885 , n7975 );
or ( n7977 , n7884 , n7976 );
and ( n7978 , n7881 , n7977 );
or ( n7979 , n7880 , n7978 );
and ( n7980 , n7877 , n7979 );
or ( n7981 , n7876 , n7980 );
and ( n7982 , n7873 , n7981 );
or ( n7983 , n7872 , n7982 );
and ( n7984 , n7869 , n7983 );
or ( n7985 , n7868 , n7984 );
and ( n7986 , n7865 , n7985 );
or ( n7987 , n7864 , n7986 );
and ( n7988 , n7861 , n7987 );
or ( n7989 , n7860 , n7988 );
and ( n7990 , n7857 , n7989 );
or ( n7991 , n7856 , n7990 );
and ( n7992 , n7853 , n7991 );
or ( n7993 , n7852 , n7992 );
and ( n7994 , n7849 , n7993 );
or ( n7995 , n7848 , n7994 );
and ( n7996 , n7845 , n7995 );
or ( n7997 , n7844 , n7996 );
and ( n7998 , n7841 , n7997 );
or ( n7999 , n7840 , n7998 );
xor ( n8000 , n7837 , n7999 );
and ( n8001 , n285 , n2299 );
nor ( n8002 , n2300 , n8001 );
nor ( n8003 , n2596 , n305 );
xor ( n8004 , n8002 , n8003 );
and ( n8005 , n7603 , n7604 );
and ( n8006 , n7605 , n7608 );
or ( n8007 , n8005 , n8006 );
xor ( n8008 , n8004 , n8007 );
nor ( n8009 , n2991 , n336 );
xor ( n8010 , n8008 , n8009 );
and ( n8011 , n7609 , n7610 );
and ( n8012 , n7611 , n7614 );
or ( n8013 , n8011 , n8012 );
xor ( n8014 , n8010 , n8013 );
nor ( n8015 , n3464 , n386 );
xor ( n8016 , n8014 , n8015 );
and ( n8017 , n7615 , n7616 );
and ( n8018 , n7617 , n7620 );
or ( n8019 , n8017 , n8018 );
xor ( n8020 , n8016 , n8019 );
nor ( n8021 , n3863 , n458 );
xor ( n8022 , n8020 , n8021 );
and ( n8023 , n7621 , n7622 );
and ( n8024 , n7623 , n7626 );
or ( n8025 , n8023 , n8024 );
xor ( n8026 , n8022 , n8025 );
nor ( n8027 , n4260 , n551 );
xor ( n8028 , n8026 , n8027 );
and ( n8029 , n7627 , n7628 );
and ( n8030 , n7629 , n7632 );
or ( n8031 , n8029 , n8030 );
xor ( n8032 , n8028 , n8031 );
nor ( n8033 , n4659 , n665 );
xor ( n8034 , n8032 , n8033 );
and ( n8035 , n7633 , n7634 );
and ( n8036 , n7635 , n7638 );
or ( n8037 , n8035 , n8036 );
xor ( n8038 , n8034 , n8037 );
nor ( n8039 , n5057 , n797 );
xor ( n8040 , n8038 , n8039 );
and ( n8041 , n7639 , n7640 );
and ( n8042 , n7641 , n7644 );
or ( n8043 , n8041 , n8042 );
xor ( n8044 , n8040 , n8043 );
nor ( n8045 , n5453 , n954 );
xor ( n8046 , n8044 , n8045 );
and ( n8047 , n7645 , n7646 );
and ( n8048 , n7647 , n7650 );
or ( n8049 , n8047 , n8048 );
xor ( n8050 , n8046 , n8049 );
nor ( n8051 , n5851 , n1128 );
xor ( n8052 , n8050 , n8051 );
and ( n8053 , n7651 , n7652 );
and ( n8054 , n7653 , n7656 );
or ( n8055 , n8053 , n8054 );
xor ( n8056 , n8052 , n8055 );
nor ( n8057 , n6249 , n1320 );
xor ( n8058 , n8056 , n8057 );
and ( n8059 , n7657 , n7658 );
and ( n8060 , n7659 , n7662 );
or ( n8061 , n8059 , n8060 );
xor ( n8062 , n8058 , n8061 );
nor ( n8063 , n6642 , n1536 );
xor ( n8064 , n8062 , n8063 );
and ( n8065 , n7663 , n7664 );
and ( n8066 , n7665 , n7668 );
or ( n8067 , n8065 , n8066 );
xor ( n8068 , n8064 , n8067 );
nor ( n8069 , n7037 , n1773 );
xor ( n8070 , n8068 , n8069 );
and ( n8071 , n7669 , n7670 );
and ( n8072 , n7671 , n7674 );
or ( n8073 , n8071 , n8072 );
xor ( n8074 , n8070 , n8073 );
nor ( n8075 , n7431 , n2027 );
xor ( n8076 , n8074 , n8075 );
and ( n8077 , n7675 , n7676 );
and ( n8078 , n7677 , n7680 );
or ( n8079 , n8077 , n8078 );
xor ( n8080 , n8076 , n8079 );
nor ( n8081 , n7824 , n2302 );
xor ( n8082 , n8080 , n8081 );
and ( n8083 , n7681 , n7682 );
and ( n8084 , n7683 , n7686 );
or ( n8085 , n8083 , n8084 );
xor ( n8086 , n8082 , n8085 );
and ( n8087 , n7704 , n7708 );
and ( n8088 , n7708 , n7712 );
and ( n8089 , n7704 , n7712 );
or ( n8090 , n8087 , n8088 , n8089 );
and ( n8091 , n7700 , n7713 );
and ( n8092 , n7713 , n7810 );
and ( n8093 , n7700 , n7810 );
or ( n8094 , n8091 , n8092 , n8093 );
xor ( n8095 , n8090 , n8094 );
and ( n8096 , n7718 , n7744 );
and ( n8097 , n7744 , n7809 );
and ( n8098 , n7718 , n7809 );
or ( n8099 , n8096 , n8097 , n8098 );
and ( n8100 , n7732 , n7733 );
and ( n8101 , n7733 , n7735 );
and ( n8102 , n7732 , n7735 );
or ( n8103 , n8100 , n8101 , n8102 );
and ( n8104 , n7722 , n7726 );
and ( n8105 , n7726 , n7743 );
and ( n8106 , n7722 , n7743 );
or ( n8107 , n8104 , n8105 , n8106 );
xor ( n8108 , n8103 , n8107 );
not ( n8109 , n2286 );
and ( n8110 , n2406 , n2286 );
nor ( n8111 , n8109 , n8110 );
xor ( n8112 , n8108 , n8111 );
xor ( n8113 , n8099 , n8112 );
and ( n8114 , n7749 , n7764 );
and ( n8115 , n7764 , n7808 );
and ( n8116 , n7749 , n7808 );
or ( n8117 , n8114 , n8115 , n8116 );
and ( n8118 , n7731 , n7736 );
and ( n8119 , n7736 , n7742 );
and ( n8120 , n7731 , n7742 );
or ( n8121 , n8118 , n8119 , n8120 );
and ( n8122 , n7753 , n7757 );
and ( n8123 , n7757 , n7763 );
and ( n8124 , n7753 , n7763 );
or ( n8125 , n8122 , n8123 , n8124 );
xor ( n8126 , n8121 , n8125 );
and ( n8127 , n7738 , n7739 );
and ( n8128 , n7739 , n7741 );
and ( n8129 , n7738 , n7741 );
or ( n8130 , n8127 , n8128 , n8129 );
and ( n8131 , n2581 , n2138 );
and ( n8132 , n2972 , n1864 );
xor ( n8133 , n8131 , n8132 );
and ( n8134 , n3445 , n1753 );
xor ( n8135 , n8133 , n8134 );
xor ( n8136 , n8130 , n8135 );
and ( n8137 , n3844 , n1396 );
and ( n8138 , n4241 , n1302 );
xor ( n8139 , n8137 , n8138 );
and ( n8140 , n4640 , n1114 );
xor ( n8141 , n8139 , n8140 );
xor ( n8142 , n8136 , n8141 );
xor ( n8143 , n8126 , n8142 );
xor ( n8144 , n8117 , n8143 );
and ( n8145 , n7769 , n7774 );
and ( n8146 , n7774 , n7807 );
and ( n8147 , n7769 , n7807 );
or ( n8148 , n8145 , n8146 , n8147 );
and ( n8149 , n7759 , n7760 );
and ( n8150 , n7760 , n7762 );
and ( n8151 , n7759 , n7762 );
or ( n8152 , n8149 , n8150 , n8151 );
and ( n8153 , n7770 , n7771 );
and ( n8154 , n7771 , n7773 );
and ( n8155 , n7770 , n7773 );
or ( n8156 , n8153 , n8154 , n8155 );
xor ( n8157 , n8152 , n8156 );
and ( n8158 , n5038 , n852 );
and ( n8159 , n5434 , n714 );
xor ( n8160 , n8158 , n8159 );
and ( n8161 , n5832 , n651 );
xor ( n8162 , n8160 , n8161 );
xor ( n8163 , n8157 , n8162 );
xor ( n8164 , n8148 , n8163 );
and ( n8165 , n7776 , n7777 );
and ( n8166 , n7777 , n7806 );
and ( n8167 , n7776 , n7806 );
or ( n8168 , n8165 , n8166 , n8167 );
and ( n8169 , n6230 , n488 );
and ( n8170 , n6623 , n411 );
xor ( n8171 , n8169 , n8170 );
and ( n8172 , n7018 , n375 );
xor ( n8173 , n8171 , n8172 );
xor ( n8174 , n8168 , n8173 );
and ( n8175 , n7412 , n312 );
and ( n8176 , n7805 , n288 );
xor ( n8177 , n8175 , n8176 );
and ( n8178 , n7788 , n7791 );
and ( n8179 , n7787 , n7792 );
xor ( n8180 , n8178 , n8179 );
and ( n8181 , n2205 , n2562 );
xor ( n8182 , n8180 , n8181 );
and ( n8183 , n7782 , n7783 );
and ( n8184 , n7783 , n7793 );
and ( n8185 , n7782 , n7793 );
or ( n8186 , n8183 , n8184 , n8185 );
xor ( n8187 , n8182 , n8186 );
and ( n8188 , n7794 , n7798 );
and ( n8189 , n7799 , n7802 );
or ( n8190 , n8188 , n8189 );
xor ( n8191 , n8187 , n8190 );
buf ( n8192 , n8191 );
buf ( n8193 , n8192 );
and ( n8194 , n8193 , n279 );
xor ( n8195 , n8177 , n8194 );
xor ( n8196 , n8174 , n8195 );
xor ( n8197 , n8164 , n8196 );
xor ( n8198 , n8144 , n8197 );
xor ( n8199 , n8113 , n8198 );
xor ( n8200 , n8095 , n8199 );
and ( n8201 , n7691 , n7695 );
and ( n8202 , n7695 , n7811 );
and ( n8203 , n7691 , n7811 );
or ( n8204 , n8201 , n8202 , n8203 );
xor ( n8205 , n8200 , n8204 );
and ( n8206 , n7812 , n7816 );
and ( n8207 , n7817 , n7820 );
or ( n8208 , n8206 , n8207 );
xor ( n8209 , n8205 , n8208 );
buf ( n8210 , n8209 );
buf ( n8211 , n8210 );
not ( n8212 , n8211 );
nor ( n8213 , n8212 , n2598 );
xor ( n8214 , n8086 , n8213 );
and ( n8215 , n7687 , n7825 );
and ( n8216 , n7826 , n7829 );
or ( n8217 , n8215 , n8216 );
xor ( n8218 , n8214 , n8217 );
buf ( n8219 , n8218 );
buf ( n8220 , n8219 );
not ( n8221 , n8220 );
buf ( n8222 , n271 );
not ( n8223 , n8222 );
nor ( n8224 , n8221 , n8223 );
xor ( n8225 , n8000 , n8224 );
xor ( n8226 , n7841 , n7997 );
nor ( n8227 , n7833 , n8223 );
and ( n8228 , n8226 , n8227 );
xor ( n8229 , n8226 , n8227 );
xor ( n8230 , n7845 , n7995 );
nor ( n8231 , n7440 , n8223 );
and ( n8232 , n8230 , n8231 );
xor ( n8233 , n8230 , n8231 );
xor ( n8234 , n7849 , n7993 );
nor ( n8235 , n7046 , n8223 );
and ( n8236 , n8234 , n8235 );
xor ( n8237 , n8234 , n8235 );
xor ( n8238 , n7853 , n7991 );
nor ( n8239 , n6651 , n8223 );
and ( n8240 , n8238 , n8239 );
xor ( n8241 , n8238 , n8239 );
xor ( n8242 , n7857 , n7989 );
nor ( n8243 , n6258 , n8223 );
and ( n8244 , n8242 , n8243 );
xor ( n8245 , n8242 , n8243 );
xor ( n8246 , n7861 , n7987 );
nor ( n8247 , n5860 , n8223 );
and ( n8248 , n8246 , n8247 );
xor ( n8249 , n8246 , n8247 );
xor ( n8250 , n7865 , n7985 );
nor ( n8251 , n5462 , n8223 );
and ( n8252 , n8250 , n8251 );
xor ( n8253 , n8250 , n8251 );
xor ( n8254 , n7869 , n7983 );
nor ( n8255 , n5066 , n8223 );
and ( n8256 , n8254 , n8255 );
xor ( n8257 , n8254 , n8255 );
xor ( n8258 , n7873 , n7981 );
nor ( n8259 , n4668 , n8223 );
and ( n8260 , n8258 , n8259 );
xor ( n8261 , n8258 , n8259 );
xor ( n8262 , n7877 , n7979 );
nor ( n8263 , n4269 , n8223 );
and ( n8264 , n8262 , n8263 );
xor ( n8265 , n8262 , n8263 );
xor ( n8266 , n7881 , n7977 );
nor ( n8267 , n3872 , n8223 );
and ( n8268 , n8266 , n8267 );
xor ( n8269 , n8266 , n8267 );
xor ( n8270 , n7885 , n7975 );
nor ( n8271 , n3473 , n8223 );
and ( n8272 , n8270 , n8271 );
xor ( n8273 , n8270 , n8271 );
xor ( n8274 , n7889 , n7973 );
nor ( n8275 , n3000 , n8223 );
and ( n8276 , n8274 , n8275 );
xor ( n8277 , n8274 , n8275 );
xor ( n8278 , n7893 , n7971 );
nor ( n8279 , n2688 , n8223 );
and ( n8280 , n8278 , n8279 );
xor ( n8281 , n8278 , n8279 );
xor ( n8282 , n7897 , n7969 );
nor ( n8283 , n3008 , n8223 );
and ( n8284 , n8282 , n8283 );
xor ( n8285 , n8282 , n8283 );
xor ( n8286 , n7901 , n7967 );
nor ( n8287 , n3017 , n8223 );
and ( n8288 , n8286 , n8287 );
xor ( n8289 , n8286 , n8287 );
xor ( n8290 , n7905 , n7965 );
nor ( n8291 , n3026 , n8223 );
and ( n8292 , n8290 , n8291 );
xor ( n8293 , n8290 , n8291 );
xor ( n8294 , n7909 , n7963 );
nor ( n8295 , n3035 , n8223 );
and ( n8296 , n8294 , n8295 );
xor ( n8297 , n8294 , n8295 );
xor ( n8298 , n7913 , n7961 );
nor ( n8299 , n3044 , n8223 );
and ( n8300 , n8298 , n8299 );
xor ( n8301 , n8298 , n8299 );
xor ( n8302 , n7917 , n7959 );
nor ( n8303 , n3053 , n8223 );
and ( n8304 , n8302 , n8303 );
xor ( n8305 , n8302 , n8303 );
xor ( n8306 , n7921 , n7957 );
nor ( n8307 , n3062 , n8223 );
and ( n8308 , n8306 , n8307 );
xor ( n8309 , n8306 , n8307 );
xor ( n8310 , n7925 , n7955 );
nor ( n8311 , n3071 , n8223 );
and ( n8312 , n8310 , n8311 );
xor ( n8313 , n8310 , n8311 );
xor ( n8314 , n7929 , n7953 );
nor ( n8315 , n3080 , n8223 );
and ( n8316 , n8314 , n8315 );
xor ( n8317 , n8314 , n8315 );
xor ( n8318 , n7933 , n7951 );
nor ( n8319 , n3089 , n8223 );
and ( n8320 , n8318 , n8319 );
xor ( n8321 , n8318 , n8319 );
xor ( n8322 , n7937 , n7949 );
nor ( n8323 , n3098 , n8223 );
and ( n8324 , n8322 , n8323 );
xor ( n8325 , n8322 , n8323 );
xor ( n8326 , n7942 , n7947 );
nor ( n8327 , n3107 , n8223 );
and ( n8328 , n8326 , n8327 );
xor ( n8329 , n8326 , n8327 );
xor ( n8330 , n7944 , n7945 );
buf ( n8331 , n8330 );
nor ( n8332 , n3116 , n8223 );
and ( n8333 , n8331 , n8332 );
xor ( n8334 , n8331 , n8332 );
nor ( n8335 , n3134 , n7835 );
buf ( n8336 , n8335 );
nor ( n8337 , n3125 , n8223 );
and ( n8338 , n8336 , n8337 );
buf ( n8339 , n8338 );
and ( n8340 , n8334 , n8339 );
or ( n8341 , n8333 , n8340 );
and ( n8342 , n8329 , n8341 );
or ( n8343 , n8328 , n8342 );
and ( n8344 , n8325 , n8343 );
or ( n8345 , n8324 , n8344 );
and ( n8346 , n8321 , n8345 );
or ( n8347 , n8320 , n8346 );
and ( n8348 , n8317 , n8347 );
or ( n8349 , n8316 , n8348 );
and ( n8350 , n8313 , n8349 );
or ( n8351 , n8312 , n8350 );
and ( n8352 , n8309 , n8351 );
or ( n8353 , n8308 , n8352 );
and ( n8354 , n8305 , n8353 );
or ( n8355 , n8304 , n8354 );
and ( n8356 , n8301 , n8355 );
or ( n8357 , n8300 , n8356 );
and ( n8358 , n8297 , n8357 );
or ( n8359 , n8296 , n8358 );
and ( n8360 , n8293 , n8359 );
or ( n8361 , n8292 , n8360 );
and ( n8362 , n8289 , n8361 );
or ( n8363 , n8288 , n8362 );
and ( n8364 , n8285 , n8363 );
or ( n8365 , n8284 , n8364 );
and ( n8366 , n8281 , n8365 );
or ( n8367 , n8280 , n8366 );
and ( n8368 , n8277 , n8367 );
or ( n8369 , n8276 , n8368 );
and ( n8370 , n8273 , n8369 );
or ( n8371 , n8272 , n8370 );
and ( n8372 , n8269 , n8371 );
or ( n8373 , n8268 , n8372 );
and ( n8374 , n8265 , n8373 );
or ( n8375 , n8264 , n8374 );
and ( n8376 , n8261 , n8375 );
or ( n8377 , n8260 , n8376 );
and ( n8378 , n8257 , n8377 );
or ( n8379 , n8256 , n8378 );
and ( n8380 , n8253 , n8379 );
or ( n8381 , n8252 , n8380 );
and ( n8382 , n8249 , n8381 );
or ( n8383 , n8248 , n8382 );
and ( n8384 , n8245 , n8383 );
or ( n8385 , n8244 , n8384 );
and ( n8386 , n8241 , n8385 );
or ( n8387 , n8240 , n8386 );
and ( n8388 , n8237 , n8387 );
or ( n8389 , n8236 , n8388 );
and ( n8390 , n8233 , n8389 );
or ( n8391 , n8232 , n8390 );
and ( n8392 , n8229 , n8391 );
or ( n8393 , n8228 , n8392 );
xor ( n8394 , n8225 , n8393 );
and ( n8395 , n285 , n2595 );
nor ( n8396 , n2596 , n8395 );
nor ( n8397 , n2991 , n305 );
xor ( n8398 , n8396 , n8397 );
and ( n8399 , n8002 , n8003 );
and ( n8400 , n8004 , n8007 );
or ( n8401 , n8399 , n8400 );
xor ( n8402 , n8398 , n8401 );
nor ( n8403 , n3464 , n336 );
xor ( n8404 , n8402 , n8403 );
and ( n8405 , n8008 , n8009 );
and ( n8406 , n8010 , n8013 );
or ( n8407 , n8405 , n8406 );
xor ( n8408 , n8404 , n8407 );
nor ( n8409 , n3863 , n386 );
xor ( n8410 , n8408 , n8409 );
and ( n8411 , n8014 , n8015 );
and ( n8412 , n8016 , n8019 );
or ( n8413 , n8411 , n8412 );
xor ( n8414 , n8410 , n8413 );
nor ( n8415 , n4260 , n458 );
xor ( n8416 , n8414 , n8415 );
and ( n8417 , n8020 , n8021 );
and ( n8418 , n8022 , n8025 );
or ( n8419 , n8417 , n8418 );
xor ( n8420 , n8416 , n8419 );
nor ( n8421 , n4659 , n551 );
xor ( n8422 , n8420 , n8421 );
and ( n8423 , n8026 , n8027 );
and ( n8424 , n8028 , n8031 );
or ( n8425 , n8423 , n8424 );
xor ( n8426 , n8422 , n8425 );
nor ( n8427 , n5057 , n665 );
xor ( n8428 , n8426 , n8427 );
and ( n8429 , n8032 , n8033 );
and ( n8430 , n8034 , n8037 );
or ( n8431 , n8429 , n8430 );
xor ( n8432 , n8428 , n8431 );
nor ( n8433 , n5453 , n797 );
xor ( n8434 , n8432 , n8433 );
and ( n8435 , n8038 , n8039 );
and ( n8436 , n8040 , n8043 );
or ( n8437 , n8435 , n8436 );
xor ( n8438 , n8434 , n8437 );
nor ( n8439 , n5851 , n954 );
xor ( n8440 , n8438 , n8439 );
and ( n8441 , n8044 , n8045 );
and ( n8442 , n8046 , n8049 );
or ( n8443 , n8441 , n8442 );
xor ( n8444 , n8440 , n8443 );
nor ( n8445 , n6249 , n1128 );
xor ( n8446 , n8444 , n8445 );
and ( n8447 , n8050 , n8051 );
and ( n8448 , n8052 , n8055 );
or ( n8449 , n8447 , n8448 );
xor ( n8450 , n8446 , n8449 );
nor ( n8451 , n6642 , n1320 );
xor ( n8452 , n8450 , n8451 );
and ( n8453 , n8056 , n8057 );
and ( n8454 , n8058 , n8061 );
or ( n8455 , n8453 , n8454 );
xor ( n8456 , n8452 , n8455 );
nor ( n8457 , n7037 , n1536 );
xor ( n8458 , n8456 , n8457 );
and ( n8459 , n8062 , n8063 );
and ( n8460 , n8064 , n8067 );
or ( n8461 , n8459 , n8460 );
xor ( n8462 , n8458 , n8461 );
nor ( n8463 , n7431 , n1773 );
xor ( n8464 , n8462 , n8463 );
and ( n8465 , n8068 , n8069 );
and ( n8466 , n8070 , n8073 );
or ( n8467 , n8465 , n8466 );
xor ( n8468 , n8464 , n8467 );
nor ( n8469 , n7824 , n2027 );
xor ( n8470 , n8468 , n8469 );
and ( n8471 , n8074 , n8075 );
and ( n8472 , n8076 , n8079 );
or ( n8473 , n8471 , n8472 );
xor ( n8474 , n8470 , n8473 );
nor ( n8475 , n8212 , n2302 );
xor ( n8476 , n8474 , n8475 );
and ( n8477 , n8080 , n8081 );
and ( n8478 , n8082 , n8085 );
or ( n8479 , n8477 , n8478 );
xor ( n8480 , n8476 , n8479 );
and ( n8481 , n8103 , n8107 );
and ( n8482 , n8107 , n8111 );
and ( n8483 , n8103 , n8111 );
or ( n8484 , n8481 , n8482 , n8483 );
and ( n8485 , n8099 , n8112 );
and ( n8486 , n8112 , n8198 );
and ( n8487 , n8099 , n8198 );
or ( n8488 , n8485 , n8486 , n8487 );
xor ( n8489 , n8484 , n8488 );
and ( n8490 , n8117 , n8143 );
and ( n8491 , n8143 , n8197 );
and ( n8492 , n8117 , n8197 );
or ( n8493 , n8490 , n8491 , n8492 );
and ( n8494 , n8131 , n8132 );
and ( n8495 , n8132 , n8134 );
and ( n8496 , n8131 , n8134 );
or ( n8497 , n8494 , n8495 , n8496 );
and ( n8498 , n8121 , n8125 );
and ( n8499 , n8125 , n8142 );
and ( n8500 , n8121 , n8142 );
or ( n8501 , n8498 , n8499 , n8500 );
xor ( n8502 , n8497 , n8501 );
not ( n8503 , n2581 );
and ( n8504 , n2406 , n2581 );
nor ( n8505 , n8503 , n8504 );
xor ( n8506 , n8502 , n8505 );
xor ( n8507 , n8493 , n8506 );
and ( n8508 , n8148 , n8163 );
and ( n8509 , n8163 , n8196 );
and ( n8510 , n8148 , n8196 );
or ( n8511 , n8508 , n8509 , n8510 );
and ( n8512 , n8130 , n8135 );
and ( n8513 , n8135 , n8141 );
and ( n8514 , n8130 , n8141 );
or ( n8515 , n8512 , n8513 , n8514 );
and ( n8516 , n8152 , n8156 );
and ( n8517 , n8156 , n8162 );
and ( n8518 , n8152 , n8162 );
or ( n8519 , n8516 , n8517 , n8518 );
xor ( n8520 , n8515 , n8519 );
and ( n8521 , n8137 , n8138 );
and ( n8522 , n8138 , n8140 );
and ( n8523 , n8137 , n8140 );
or ( n8524 , n8521 , n8522 , n8523 );
and ( n8525 , n2972 , n2138 );
and ( n8526 , n3445 , n1864 );
xor ( n8527 , n8525 , n8526 );
and ( n8528 , n3844 , n1753 );
xor ( n8529 , n8527 , n8528 );
xor ( n8530 , n8524 , n8529 );
and ( n8531 , n4241 , n1396 );
and ( n8532 , n4640 , n1302 );
xor ( n8533 , n8531 , n8532 );
and ( n8534 , n5038 , n1114 );
xor ( n8535 , n8533 , n8534 );
xor ( n8536 , n8530 , n8535 );
xor ( n8537 , n8520 , n8536 );
xor ( n8538 , n8511 , n8537 );
and ( n8539 , n8168 , n8173 );
and ( n8540 , n8173 , n8195 );
and ( n8541 , n8168 , n8195 );
or ( n8542 , n8539 , n8540 , n8541 );
and ( n8543 , n8158 , n8159 );
and ( n8544 , n8159 , n8161 );
and ( n8545 , n8158 , n8161 );
or ( n8546 , n8543 , n8544 , n8545 );
and ( n8547 , n8169 , n8170 );
and ( n8548 , n8170 , n8172 );
and ( n8549 , n8169 , n8172 );
or ( n8550 , n8547 , n8548 , n8549 );
xor ( n8551 , n8546 , n8550 );
and ( n8552 , n5434 , n852 );
and ( n8553 , n5832 , n714 );
xor ( n8554 , n8552 , n8553 );
and ( n8555 , n6230 , n651 );
xor ( n8556 , n8554 , n8555 );
xor ( n8557 , n8551 , n8556 );
xor ( n8558 , n8542 , n8557 );
and ( n8559 , n8175 , n8176 );
and ( n8560 , n8176 , n8194 );
and ( n8561 , n8175 , n8194 );
or ( n8562 , n8559 , n8560 , n8561 );
and ( n8563 , n6623 , n488 );
and ( n8564 , n7018 , n411 );
xor ( n8565 , n8563 , n8564 );
and ( n8566 , n7412 , n375 );
xor ( n8567 , n8565 , n8566 );
xor ( n8568 , n8562 , n8567 );
and ( n8569 , n7805 , n312 );
and ( n8570 , n8193 , n288 );
xor ( n8571 , n8569 , n8570 );
and ( n8572 , n8179 , n8181 );
and ( n8573 , n8178 , n8181 );
or ( n8574 , 1'b0 , n8572 , n8573 );
and ( n8575 , n8182 , n8186 );
and ( n8576 , n8187 , n8190 );
or ( n8577 , n8575 , n8576 );
xor ( n8578 , n8574 , n8577 );
buf ( n8579 , n8578 );
buf ( n8580 , n8579 );
not ( n8581 , n8580 );
and ( n8582 , n8581 , n279 );
not ( n8583 , n279 );
nor ( n8584 , n8582 , n8583 );
xor ( n8585 , n8571 , n8584 );
xor ( n8586 , n8568 , n8585 );
xor ( n8587 , n8558 , n8586 );
xor ( n8588 , n8538 , n8587 );
xor ( n8589 , n8507 , n8588 );
xor ( n8590 , n8489 , n8589 );
and ( n8591 , n8090 , n8094 );
and ( n8592 , n8094 , n8199 );
and ( n8593 , n8090 , n8199 );
or ( n8594 , n8591 , n8592 , n8593 );
xor ( n8595 , n8590 , n8594 );
and ( n8596 , n8200 , n8204 );
and ( n8597 , n8205 , n8208 );
or ( n8598 , n8596 , n8597 );
xor ( n8599 , n8595 , n8598 );
buf ( n8600 , n8599 );
buf ( n8601 , n8600 );
not ( n8602 , n8601 );
nor ( n8603 , n8602 , n2598 );
xor ( n8604 , n8480 , n8603 );
and ( n8605 , n8086 , n8213 );
and ( n8606 , n8214 , n8217 );
or ( n8607 , n8605 , n8606 );
xor ( n8608 , n8604 , n8607 );
buf ( n8609 , n8608 );
buf ( n8610 , n8609 );
not ( n8611 , n8610 );
buf ( n8612 , n272 );
not ( n8613 , n8612 );
nor ( n8614 , n8611 , n8613 );
xor ( n8615 , n8394 , n8614 );
xor ( n8616 , n8229 , n8391 );
nor ( n8617 , n8221 , n8613 );
and ( n8618 , n8616 , n8617 );
xor ( n8619 , n8616 , n8617 );
xor ( n8620 , n8233 , n8389 );
nor ( n8621 , n7833 , n8613 );
and ( n8622 , n8620 , n8621 );
xor ( n8623 , n8620 , n8621 );
xor ( n8624 , n8237 , n8387 );
nor ( n8625 , n7440 , n8613 );
and ( n8626 , n8624 , n8625 );
xor ( n8627 , n8624 , n8625 );
xor ( n8628 , n8241 , n8385 );
nor ( n8629 , n7046 , n8613 );
and ( n8630 , n8628 , n8629 );
xor ( n8631 , n8628 , n8629 );
xor ( n8632 , n8245 , n8383 );
nor ( n8633 , n6651 , n8613 );
and ( n8634 , n8632 , n8633 );
xor ( n8635 , n8632 , n8633 );
xor ( n8636 , n8249 , n8381 );
nor ( n8637 , n6258 , n8613 );
and ( n8638 , n8636 , n8637 );
xor ( n8639 , n8636 , n8637 );
xor ( n8640 , n8253 , n8379 );
nor ( n8641 , n5860 , n8613 );
and ( n8642 , n8640 , n8641 );
xor ( n8643 , n8640 , n8641 );
xor ( n8644 , n8257 , n8377 );
nor ( n8645 , n5462 , n8613 );
and ( n8646 , n8644 , n8645 );
xor ( n8647 , n8644 , n8645 );
xor ( n8648 , n8261 , n8375 );
nor ( n8649 , n5066 , n8613 );
and ( n8650 , n8648 , n8649 );
xor ( n8651 , n8648 , n8649 );
xor ( n8652 , n8265 , n8373 );
nor ( n8653 , n4668 , n8613 );
and ( n8654 , n8652 , n8653 );
xor ( n8655 , n8652 , n8653 );
xor ( n8656 , n8269 , n8371 );
nor ( n8657 , n4269 , n8613 );
and ( n8658 , n8656 , n8657 );
xor ( n8659 , n8656 , n8657 );
xor ( n8660 , n8273 , n8369 );
nor ( n8661 , n3872 , n8613 );
and ( n8662 , n8660 , n8661 );
xor ( n8663 , n8660 , n8661 );
xor ( n8664 , n8277 , n8367 );
nor ( n8665 , n3473 , n8613 );
and ( n8666 , n8664 , n8665 );
xor ( n8667 , n8664 , n8665 );
xor ( n8668 , n8281 , n8365 );
nor ( n8669 , n3000 , n8613 );
and ( n8670 , n8668 , n8669 );
xor ( n8671 , n8668 , n8669 );
xor ( n8672 , n8285 , n8363 );
nor ( n8673 , n2688 , n8613 );
and ( n8674 , n8672 , n8673 );
xor ( n8675 , n8672 , n8673 );
xor ( n8676 , n8289 , n8361 );
nor ( n8677 , n3008 , n8613 );
and ( n8678 , n8676 , n8677 );
xor ( n8679 , n8676 , n8677 );
xor ( n8680 , n8293 , n8359 );
nor ( n8681 , n3017 , n8613 );
and ( n8682 , n8680 , n8681 );
xor ( n8683 , n8680 , n8681 );
xor ( n8684 , n8297 , n8357 );
nor ( n8685 , n3026 , n8613 );
and ( n8686 , n8684 , n8685 );
xor ( n8687 , n8684 , n8685 );
xor ( n8688 , n8301 , n8355 );
nor ( n8689 , n3035 , n8613 );
and ( n8690 , n8688 , n8689 );
xor ( n8691 , n8688 , n8689 );
xor ( n8692 , n8305 , n8353 );
nor ( n8693 , n3044 , n8613 );
and ( n8694 , n8692 , n8693 );
xor ( n8695 , n8692 , n8693 );
xor ( n8696 , n8309 , n8351 );
nor ( n8697 , n3053 , n8613 );
and ( n8698 , n8696 , n8697 );
xor ( n8699 , n8696 , n8697 );
xor ( n8700 , n8313 , n8349 );
nor ( n8701 , n3062 , n8613 );
and ( n8702 , n8700 , n8701 );
xor ( n8703 , n8700 , n8701 );
xor ( n8704 , n8317 , n8347 );
nor ( n8705 , n3071 , n8613 );
and ( n8706 , n8704 , n8705 );
xor ( n8707 , n8704 , n8705 );
xor ( n8708 , n8321 , n8345 );
nor ( n8709 , n3080 , n8613 );
and ( n8710 , n8708 , n8709 );
xor ( n8711 , n8708 , n8709 );
xor ( n8712 , n8325 , n8343 );
nor ( n8713 , n3089 , n8613 );
and ( n8714 , n8712 , n8713 );
xor ( n8715 , n8712 , n8713 );
xor ( n8716 , n8329 , n8341 );
nor ( n8717 , n3098 , n8613 );
and ( n8718 , n8716 , n8717 );
xor ( n8719 , n8716 , n8717 );
xor ( n8720 , n8334 , n8339 );
nor ( n8721 , n3107 , n8613 );
and ( n8722 , n8720 , n8721 );
xor ( n8723 , n8720 , n8721 );
xor ( n8724 , n8336 , n8337 );
buf ( n8725 , n8724 );
nor ( n8726 , n3116 , n8613 );
and ( n8727 , n8725 , n8726 );
xor ( n8728 , n8725 , n8726 );
nor ( n8729 , n3134 , n8223 );
buf ( n8730 , n8729 );
nor ( n8731 , n3125 , n8613 );
and ( n8732 , n8730 , n8731 );
buf ( n8733 , n8732 );
and ( n8734 , n8728 , n8733 );
or ( n8735 , n8727 , n8734 );
and ( n8736 , n8723 , n8735 );
or ( n8737 , n8722 , n8736 );
and ( n8738 , n8719 , n8737 );
or ( n8739 , n8718 , n8738 );
and ( n8740 , n8715 , n8739 );
or ( n8741 , n8714 , n8740 );
and ( n8742 , n8711 , n8741 );
or ( n8743 , n8710 , n8742 );
and ( n8744 , n8707 , n8743 );
or ( n8745 , n8706 , n8744 );
and ( n8746 , n8703 , n8745 );
or ( n8747 , n8702 , n8746 );
and ( n8748 , n8699 , n8747 );
or ( n8749 , n8698 , n8748 );
and ( n8750 , n8695 , n8749 );
or ( n8751 , n8694 , n8750 );
and ( n8752 , n8691 , n8751 );
or ( n8753 , n8690 , n8752 );
and ( n8754 , n8687 , n8753 );
or ( n8755 , n8686 , n8754 );
and ( n8756 , n8683 , n8755 );
or ( n8757 , n8682 , n8756 );
and ( n8758 , n8679 , n8757 );
or ( n8759 , n8678 , n8758 );
and ( n8760 , n8675 , n8759 );
or ( n8761 , n8674 , n8760 );
and ( n8762 , n8671 , n8761 );
or ( n8763 , n8670 , n8762 );
and ( n8764 , n8667 , n8763 );
or ( n8765 , n8666 , n8764 );
and ( n8766 , n8663 , n8765 );
or ( n8767 , n8662 , n8766 );
and ( n8768 , n8659 , n8767 );
or ( n8769 , n8658 , n8768 );
and ( n8770 , n8655 , n8769 );
or ( n8771 , n8654 , n8770 );
and ( n8772 , n8651 , n8771 );
or ( n8773 , n8650 , n8772 );
and ( n8774 , n8647 , n8773 );
or ( n8775 , n8646 , n8774 );
and ( n8776 , n8643 , n8775 );
or ( n8777 , n8642 , n8776 );
and ( n8778 , n8639 , n8777 );
or ( n8779 , n8638 , n8778 );
and ( n8780 , n8635 , n8779 );
or ( n8781 , n8634 , n8780 );
and ( n8782 , n8631 , n8781 );
or ( n8783 , n8630 , n8782 );
and ( n8784 , n8627 , n8783 );
or ( n8785 , n8626 , n8784 );
and ( n8786 , n8623 , n8785 );
or ( n8787 , n8622 , n8786 );
and ( n8788 , n8619 , n8787 );
or ( n8789 , n8618 , n8788 );
xor ( n8790 , n8615 , n8789 );
buf ( n8791 , n8790 );
buf ( n8792 , n8791 );
xor ( n8793 , n8619 , n8787 );
buf ( n8794 , n8793 );
buf ( n8795 , n8794 );
xor ( n8796 , n8623 , n8785 );
buf ( n8797 , n8796 );
buf ( n8798 , n8797 );
xor ( n8799 , n8627 , n8783 );
buf ( n8800 , n8799 );
buf ( n8801 , n8800 );
xor ( n8802 , n8631 , n8781 );
buf ( n8803 , n8802 );
buf ( n8804 , n8803 );
xor ( n8805 , n8635 , n8779 );
buf ( n8806 , n8805 );
buf ( n8807 , n8806 );
xor ( n8808 , n8639 , n8777 );
buf ( n8809 , n8808 );
buf ( n8810 , n8809 );
xor ( n8811 , n8643 , n8775 );
buf ( n8812 , n8811 );
buf ( n8813 , n8812 );
xor ( n8814 , n8647 , n8773 );
buf ( n8815 , n8814 );
buf ( n8816 , n8815 );
xor ( n8817 , n8651 , n8771 );
buf ( n8818 , n8817 );
buf ( n8819 , n8818 );
xor ( n8820 , n8655 , n8769 );
buf ( n8821 , n8820 );
buf ( n8822 , n8821 );
xor ( n8823 , n8659 , n8767 );
buf ( n8824 , n8823 );
buf ( n8825 , n8824 );
xor ( n8826 , n8663 , n8765 );
buf ( n8827 , n8826 );
buf ( n8828 , n8827 );
xor ( n8829 , n8667 , n8763 );
buf ( n8830 , n8829 );
buf ( n8831 , n8830 );
xor ( n8832 , n8671 , n8761 );
buf ( n8833 , n8832 );
buf ( n8834 , n8833 );
xor ( n8835 , n8675 , n8759 );
buf ( n8836 , n8835 );
buf ( n8837 , n8836 );
endmodule

