//
// Conformal-LEC Version 16.10-d005 ( 21-Apr-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 ;
output n2048 , n2049 ;

wire n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , 
     n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , 
     n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , 
     n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , 
     n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , 
     n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , 
     n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , 
     n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , 
     n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , 
     n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , 
     n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , 
     n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , 
     n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , 
     n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , 
     n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , 
     n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , 
     n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , 
     n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , 
     n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , 
     n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , 
     n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , 
     n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , 
     n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , 
     n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , 
     n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , 
     n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , 
     n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , 
     n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , 
     n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , 
     n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , 
     n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , 
     n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , 
     n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , 
     n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , 
     n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , 
     n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , 
     n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , 
     n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , 
     n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , 
     n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , 
     n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , 
     n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , 
     n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , 
     n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , 
     n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , 
     n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , 
     n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , 
     n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , 
     n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , 
     n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , 
     n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , 
     n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , 
     n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , 
     n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , 
     n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , 
     n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , 
     n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , 
     n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , 
     n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , 
     n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , 
     n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , 
     n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , 
     n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , 
     n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , 
     n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , 
     n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , 
     n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , 
     n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , 
     n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , 
     n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , 
     n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , 
     n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , 
     n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , 
     n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , 
     n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , 
     n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , 
     n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , 
     n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , 
     n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , 
     n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , 
     n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , 
     n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , 
     n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , 
     n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , 
     n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , 
     n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , 
     n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , 
     n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , 
     n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , 
     n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , 
     n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , 
     n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , 
     n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , 
     n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , 
     n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , 
     n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , 
     n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , 
     n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , 
     n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , 
     n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , 
     n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , 
     n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , 
     n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , 
     n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , 
     n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , 
     n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , 
     n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , 
     n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , 
     n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , 
     n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , 
     n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , 
     n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , 
     n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , 
     n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , 
     n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , 
     n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , 
     n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , 
     n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , 
     n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , 
     n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , 
     n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , 
     n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , 
     n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , 
     n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , 
     n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , 
     n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , 
     n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , 
     n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , 
     n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , 
     n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , 
     n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , 
     n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , 
     n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , 
     n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , 
     n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , 
     n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , 
     n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , 
     n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , 
     n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , 
     n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , 
     n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , 
     n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , 
     n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , 
     n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , 
     n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , 
     n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , 
     n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , 
     n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , 
     n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , 
     n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , 
     n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , 
     n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , 
     n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , 
     n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , 
     n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , 
     n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , 
     n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , 
     n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , 
     n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , 
     n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , 
     n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , 
     n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , 
     n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , 
     n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , 
     n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , 
     n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , 
     n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , 
     n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , 
     n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , 
     n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , 
     n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , 
     n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , 
     n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , 
     n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , 
     n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , 
     n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , 
     n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , 
     n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , 
     n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , 
     n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , 
     n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , 
     n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , 
     n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , 
     n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , 
     n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , 
     n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , 
     n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , 
     n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , 
     n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , 
     n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , 
     n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , 
     n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , 
     n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , 
     n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , 
     n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , 
     n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , 
     n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , 
     n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , 
     n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , 
     n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , 
     n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , 
     n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , 
     n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , 
     n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , 
     n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , 
     n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , 
     n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , 
     n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , 
     n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , 
     n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , 
     n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , 
     n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , 
     n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , 
     n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , 
     n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , 
     n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , 
     n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , 
     n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , 
     n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , 
     n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , 
     n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , 
     n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , 
     n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , 
     n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , 
     n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , 
     n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , 
     n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , 
     n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , 
     n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , 
     n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , 
     n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , 
     n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , 
     n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , 
     n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , 
     n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , 
     n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , 
     n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , 
     n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , 
     n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , 
     n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , 
     n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , 
     n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , 
     n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , 
     n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , 
     n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , 
     n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , 
     n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , 
     n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , 
     n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , 
     n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , 
     n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , 
     n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , 
     n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , 
     n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , 
     n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , 
     n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , 
     n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , 
     n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , 
     n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , 
     n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , 
     n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , 
     n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , 
     n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , 
     n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , 
     n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , 
     n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , 
     n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , 
     n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , 
     n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , 
     n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , 
     n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , 
     n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , 
     n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , 
     n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , 
     n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , 
     n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , 
     n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , 
     n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , 
     n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , 
     n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , 
     n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , 
     n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , 
     n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , 
     n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , 
     n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , 
     n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , 
     n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , 
     n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , 
     n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , 
     n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , 
     n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , 
     n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , 
     n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , 
     n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , 
     n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , 
     n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , 
     n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , 
     n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , 
     n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , 
     n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , 
     n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , 
     n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , 
     n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , 
     n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , 
     n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , 
     n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , 
     n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , 
     n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , 
     n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , 
     n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , 
     n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , 
     n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , 
     n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , 
     n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , 
     n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , 
     n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , 
     n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , 
     n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , 
     n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , 
     n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , 
     n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , 
     n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , 
     n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , 
     n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , 
     n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , 
     n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , 
     n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , 
     n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , 
     n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , 
     n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , 
     n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , 
     n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , 
     n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , 
     n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , 
     n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , 
     n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , 
     n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , 
     n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , 
     n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , 
     n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , 
     n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , 
     n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , 
     n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , 
     n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , 
     n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , 
     n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , 
     n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , 
     n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , 
     n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , 
     n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , 
     n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , 
     n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , 
     n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , 
     n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , 
     n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , 
     n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , 
     n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , 
     n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , 
     n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , 
     n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , 
     n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , 
     n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , 
     n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , 
     n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , 
     n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , 
     n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , 
     n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , 
     n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , 
     n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , 
     n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , 
     n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , 
     n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , 
     n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , 
     n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , 
     n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , 
     n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , 
     n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , 
     n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , 
     n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , 
     n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , 
     n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , 
     n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , 
     n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , 
     n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , 
     n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , 
     n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , 
     n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , 
     n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , 
     n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , 
     n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , 
     n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , 
     n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , 
     n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , 
     n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , 
     n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , 
     n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , 
     n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , 
     n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , 
     n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , 
     n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , 
     n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , 
     n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , 
     n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , 
     n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , 
     n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , 
     n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , 
     n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , 
     n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , 
     n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , 
     n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , 
     n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , 
     n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , 
     n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , 
     n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , 
     n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , 
     n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , 
     n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , 
     n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , 
     n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , 
     n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , 
     n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , 
     n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , 
     n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , 
     n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , 
     n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , 
     n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , 
     n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , 
     n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , 
     n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , 
     n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , 
     n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , 
     n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , 
     n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , 
     n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , 
     n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , 
     n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , 
     n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , 
     n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , 
     n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , 
     n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , 
     n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , 
     n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , 
     n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , 
     n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , 
     n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , 
     n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , 
     n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , 
     n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , 
     n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , 
     n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , 
     n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , 
     n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , 
     n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , 
     n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , 
     n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , 
     n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , 
     n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , 
     n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , 
     n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , 
     n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , 
     n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , 
     n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , 
     n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , 
     n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , 
     n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , 
     n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , 
     n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , 
     n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , 
     n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , 
     n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , 
     n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , 
     n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , 
     n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , 
     n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , 
     n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , 
     n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , 
     n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , 
     n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , 
     n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , 
     n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , 
     n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , 
     n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , 
     n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , 
     n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , 
     n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , 
     n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , 
     n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , 
     n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , 
     n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , 
     n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , 
     n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , 
     n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , 
     n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , 
     n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , 
     n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , 
     n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , 
     n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , 
     n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , 
     n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , 
     n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , 
     n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , 
     n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , 
     n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , 
     n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , 
     n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , 
     n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , 
     n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , 
     n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , 
     n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , 
     n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , 
     n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , 
     n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , 
     n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , 
     n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , 
     n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , 
     n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , 
     n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , 
     n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , 
     n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , 
     n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , 
     n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , 
     n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , 
     n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , 
     n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , 
     n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , 
     n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , 
     n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , 
     n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , 
     n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , 
     n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , 
     n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , 
     n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , 
     n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , 
     n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , 
     n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , 
     n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , 
     n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , 
     n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , 
     n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , 
     n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , 
     n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , 
     n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , 
     n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , 
     n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , 
     n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , 
     n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , 
     n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , 
     n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , 
     n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , 
     n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , 
     n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , 
     n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , 
     n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , 
     n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , 
     n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , 
     n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , 
     n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , 
     n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , 
     n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , 
     n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , 
     n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , 
     n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , 
     n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , 
     n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , 
     n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , 
     n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , 
     n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , 
     n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , 
     n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , 
     n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , 
     n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , 
     n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , 
     n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , 
     n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , 
     n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , 
     n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , 
     n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , 
     n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , 
     n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , 
     n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , 
     n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , 
     n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , 
     n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , 
     n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , 
     n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , 
     n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , 
     n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , 
     n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , 
     n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , 
     n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , 
     n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , 
     n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , 
     n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , 
     n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , 
     n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , 
     n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , 
     n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , 
     n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , 
     n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , 
     n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , 
     n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , 
     n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , 
     n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , 
     n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , 
     n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , 
     n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , 
     n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , 
     n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , 
     n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , 
     n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , 
     n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , 
     n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , 
     n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , 
     n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , 
     n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , 
     n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , 
     n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , 
     n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , 
     n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , 
     n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , 
     n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , 
     n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , 
     n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , 
     n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , 
     n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , 
     n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , 
     n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , 
     n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , 
     n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , 
     n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , 
     n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , 
     n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , 
     n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , 
     n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , 
     n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , 
     n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , 
     n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , 
     n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , 
     n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , 
     n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , 
     n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , 
     n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , 
     n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , 
     n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , 
     n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , 
     n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , 
     n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , 
     n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , 
     n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , 
     n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , 
     n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , 
     n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , 
     n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , 
     n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , 
     n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , 
     n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , 
     n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , 
     n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , 
     n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , 
     n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , 
     n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , 
     n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , 
     n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , 
     n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , 
     n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , 
     n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , 
     n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , 
     n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , 
     n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , 
     n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , 
     n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , 
     n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , 
     n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , 
     n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , 
     n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , 
     n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , 
     n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , 
     n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , 
     n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , 
     n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , 
     n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , 
     n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , 
     n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , 
     n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , 
     n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , 
     n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , 
     n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , 
     n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , 
     n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , 
     n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , 
     n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , 
     n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , 
     n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , 
     n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , 
     n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , 
     n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , 
     n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , 
     n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , 
     n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , 
     n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , 
     n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , 
     n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , 
     n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , 
     n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , 
     n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , 
     n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , 
     n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , 
     n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , 
     n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , 
     n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , 
     n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , 
     n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , 
     n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , 
     n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , 
     n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , 
     n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , 
     n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , 
     n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , 
     n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , 
     n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , 
     n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , 
     n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , 
     n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , 
     n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , 
     n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , 
     n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , 
     n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , 
     n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , 
     n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , 
     n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , 
     n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , 
     n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , 
     n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , 
     n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , 
     n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , 
     n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , 
     n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , 
     n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , 
     n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , 
     n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , 
     n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , 
     n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , 
     n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , 
     n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , 
     n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , 
     n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , 
     n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , 
     n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , 
     n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , 
     n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , 
     n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , 
     n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , 
     n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , 
     n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , 
     n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , 
     n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , 
     n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , 
     n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , 
     n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , 
     n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , 
     n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , 
     n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , 
     n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , 
     n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , 
     n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , 
     n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , 
     n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , 
     n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , 
     n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , 
     n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , 
     n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , 
     n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , 
     n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , 
     n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , 
     n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , 
     n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , 
     n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , 
     n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , 
     n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , 
     n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , 
     n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , 
     n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , 
     n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , 
     n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , 
     n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , 
     n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , 
     n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , 
     n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , 
     n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , 
     n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , 
     n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , 
     n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , 
     n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , 
     n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , 
     n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , 
     n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , 
     n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , 
     n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , 
     n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , 
     n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , 
     n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , 
     n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , 
     n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , 
     n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , 
     n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , 
     n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , 
     n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , 
     n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , 
     n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , 
     n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , 
     n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , 
     n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , 
     n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , 
     n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , 
     n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , 
     n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , 
     n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , 
     n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , 
     n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , 
     n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , 
     n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , 
     n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , 
     n12319 ;
buf ( n2049 , n8230 );
buf ( n2048 , n12319 );
buf ( n4102 , n1034 );
buf ( n4103 , n1592 );
buf ( n4104 , n603 );
buf ( n4105 , n200 );
buf ( n4106 , n1580 );
buf ( n4107 , n605 );
buf ( n4108 , n1607 );
buf ( n4109 , n1303 );
buf ( n4110 , n1812 );
buf ( n4111 , n1722 );
buf ( n4112 , n331 );
buf ( n4113 , n519 );
buf ( n4114 , n1521 );
buf ( n4115 , n2043 );
buf ( n4116 , n968 );
buf ( n4117 , n239 );
buf ( n4118 , n1450 );
buf ( n4119 , n711 );
buf ( n4120 , n139 );
buf ( n4121 , n640 );
buf ( n4122 , n1570 );
buf ( n4123 , n1898 );
buf ( n4124 , n1140 );
buf ( n4125 , n1586 );
buf ( n4126 , n1479 );
buf ( n4127 , n197 );
buf ( n4128 , n1579 );
buf ( n4129 , n1588 );
buf ( n4130 , n1384 );
buf ( n4131 , n1772 );
buf ( n4132 , n42 );
buf ( n4133 , n196 );
buf ( n4134 , n1274 );
buf ( n4135 , n1259 );
buf ( n4136 , n1223 );
buf ( n4137 , n1466 );
buf ( n4138 , n932 );
buf ( n4139 , n849 );
buf ( n4140 , n166 );
buf ( n4141 , n269 );
buf ( n4142 , n1454 );
buf ( n4143 , n513 );
buf ( n4144 , n1201 );
buf ( n4145 , n428 );
buf ( n4146 , n1745 );
buf ( n4147 , n1290 );
buf ( n4148 , n1950 );
buf ( n4149 , n1769 );
buf ( n4150 , n1126 );
buf ( n4151 , n1119 );
buf ( n4152 , n62 );
buf ( n4153 , n67 );
buf ( n4154 , n1306 );
buf ( n4155 , n50 );
buf ( n4156 , n412 );
buf ( n4157 , n477 );
buf ( n4158 , n1678 );
buf ( n4159 , n1826 );
buf ( n4160 , n108 );
buf ( n4161 , n504 );
buf ( n4162 , n116 );
buf ( n4163 , n1979 );
buf ( n4164 , n1214 );
buf ( n4165 , n1092 );
buf ( n4166 , n620 );
buf ( n4167 , n1339 );
buf ( n4168 , n533 );
buf ( n4169 , n1374 );
buf ( n4170 , n153 );
buf ( n4171 , n1787 );
buf ( n4172 , n332 );
buf ( n4173 , n317 );
buf ( n4174 , n273 );
buf ( n4175 , n1221 );
buf ( n4176 , n921 );
buf ( n4177 , n1493 );
buf ( n4178 , n1297 );
buf ( n4179 , n452 );
buf ( n4180 , n319 );
buf ( n4181 , n2012 );
buf ( n4182 , n365 );
buf ( n4183 , n442 );
buf ( n4184 , n824 );
buf ( n4185 , n1855 );
buf ( n4186 , n105 );
buf ( n4187 , n421 );
buf ( n4188 , n1704 );
buf ( n4189 , n1863 );
buf ( n4190 , n1512 );
buf ( n4191 , n1325 );
buf ( n4192 , n1867 );
buf ( n4193 , n1362 );
buf ( n4194 , n143 );
buf ( n4195 , n486 );
buf ( n4196 , n1546 );
buf ( n4197 , n1947 );
buf ( n4198 , n543 );
buf ( n4199 , n1050 );
buf ( n4200 , n604 );
buf ( n4201 , n725 );
buf ( n4202 , n1878 );
buf ( n4203 , n1616 );
buf ( n4204 , n1228 );
buf ( n4205 , n422 );
buf ( n4206 , n1539 );
buf ( n4207 , n1727 );
buf ( n4208 , n910 );
buf ( n4209 , n1079 );
buf ( n4210 , n1977 );
buf ( n4211 , n393 );
buf ( n4212 , n1107 );
buf ( n4213 , n10 );
buf ( n4214 , n696 );
buf ( n4215 , n606 );
buf ( n4216 , n1625 );
buf ( n4217 , n1915 );
buf ( n4218 , n133 );
buf ( n4219 , n23 );
buf ( n4220 , n2035 );
buf ( n4221 , n1970 );
buf ( n4222 , n1462 );
buf ( n4223 , n549 );
buf ( n4224 , n236 );
buf ( n4225 , n1052 );
buf ( n4226 , n903 );
buf ( n4227 , n520 );
buf ( n4228 , n447 );
buf ( n4229 , n17 );
buf ( n4230 , n76 );
buf ( n4231 , n1061 );
buf ( n4232 , n354 );
buf ( n4233 , n1830 );
buf ( n4234 , n1721 );
buf ( n4235 , n212 );
buf ( n4236 , n1912 );
buf ( n4237 , n61 );
buf ( n4238 , n288 );
buf ( n4239 , n1525 );
buf ( n4240 , n850 );
buf ( n4241 , n1729 );
buf ( n4242 , n1265 );
buf ( n4243 , n1491 );
buf ( n4244 , n453 );
buf ( n4245 , n780 );
buf ( n4246 , n1463 );
buf ( n4247 , n267 );
buf ( n4248 , n1480 );
buf ( n4249 , n841 );
buf ( n4250 , n250 );
buf ( n4251 , n1299 );
buf ( n4252 , n1406 );
buf ( n4253 , n207 );
buf ( n4254 , n807 );
buf ( n4255 , n814 );
buf ( n4256 , n713 );
buf ( n4257 , n1846 );
buf ( n4258 , n72 );
buf ( n4259 , n485 );
buf ( n4260 , n1414 );
buf ( n4261 , n6 );
buf ( n4262 , n1139 );
buf ( n4263 , n1674 );
buf ( n4264 , n931 );
buf ( n4265 , n1386 );
buf ( n4266 , n1023 );
buf ( n4267 , n1888 );
buf ( n4268 , n114 );
buf ( n4269 , n2013 );
buf ( n4270 , n854 );
buf ( n4271 , n141 );
buf ( n4272 , n709 );
buf ( n4273 , n1753 );
buf ( n4274 , n1695 );
buf ( n4275 , n381 );
buf ( n4276 , n1518 );
buf ( n4277 , n348 );
buf ( n4278 , n1789 );
buf ( n4279 , n1123 );
buf ( n4280 , n85 );
buf ( n4281 , n1442 );
buf ( n4282 , n2047 );
buf ( n4283 , n411 );
buf ( n4284 , n661 );
buf ( n4285 , n118 );
buf ( n4286 , n1815 );
buf ( n4287 , n482 );
buf ( n4288 , n457 );
buf ( n4289 , n460 );
buf ( n4290 , n906 );
buf ( n4291 , n1756 );
buf ( n4292 , n917 );
buf ( n4293 , n612 );
buf ( n4294 , n1711 );
buf ( n4295 , n2019 );
buf ( n4296 , n1051 );
buf ( n4297 , n1664 );
buf ( n4298 , n619 );
buf ( n4299 , n1540 );
buf ( n4300 , n1234 );
buf ( n4301 , n461 );
buf ( n4302 , n1193 );
buf ( n4303 , n1305 );
buf ( n4304 , n1268 );
buf ( n4305 , n1792 );
buf ( n4306 , n78 );
buf ( n4307 , n1513 );
buf ( n4308 , n1937 );
buf ( n4309 , n1387 );
buf ( n4310 , n1459 );
buf ( n4311 , n803 );
buf ( n4312 , n530 );
buf ( n4313 , n1300 );
buf ( n4314 , n602 );
buf ( n4315 , n1901 );
buf ( n4316 , n1866 );
buf ( n4317 , n1658 );
buf ( n4318 , n318 );
buf ( n4319 , n1966 );
buf ( n4320 , n1243 );
buf ( n4321 , n601 );
buf ( n4322 , n515 );
buf ( n4323 , n21 );
buf ( n4324 , n1741 );
buf ( n4325 , n753 );
buf ( n4326 , n1334 );
buf ( n4327 , n1522 );
buf ( n4328 , n480 );
buf ( n4329 , n792 );
buf ( n4330 , n1983 );
buf ( n4331 , n1085 );
buf ( n4332 , n426 );
buf ( n4333 , n728 );
buf ( n4334 , n1785 );
buf ( n4335 , n364 );
buf ( n4336 , n275 );
buf ( n4337 , n1993 );
buf ( n4338 , n1652 );
buf ( n4339 , n1408 );
buf ( n4340 , n1590 );
buf ( n4341 , n801 );
buf ( n4342 , n403 );
buf ( n4343 , n87 );
buf ( n4344 , n900 );
buf ( n4345 , n208 );
buf ( n4346 , n636 );
buf ( n4347 , n205 );
buf ( n4348 , n534 );
buf ( n4349 , n1739 );
buf ( n4350 , n1360 );
buf ( n4351 , n1895 );
buf ( n4352 , n1113 );
buf ( n4353 , n2041 );
buf ( n4354 , n419 );
buf ( n4355 , n1015 );
buf ( n4356 , n1449 );
buf ( n4357 , n1240 );
buf ( n4358 , n537 );
buf ( n4359 , n1719 );
buf ( n4360 , n1885 );
buf ( n4361 , n1301 );
buf ( n4362 , n876 );
buf ( n4363 , n1563 );
buf ( n4364 , n104 );
buf ( n4365 , n1813 );
buf ( n4366 , n993 );
buf ( n4367 , n1533 );
buf ( n4368 , n1634 );
buf ( n4369 , n1713 );
buf ( n4370 , n1246 );
buf ( n4371 , n1037 );
buf ( n4372 , n1069 );
buf ( n4373 , n981 );
buf ( n4374 , n1531 );
buf ( n4375 , n1500 );
buf ( n4376 , n242 );
buf ( n4377 , n132 );
buf ( n4378 , n215 );
buf ( n4379 , n1419 );
buf ( n4380 , n443 );
buf ( n4381 , n1110 );
buf ( n4382 , n135 );
buf ( n4383 , n333 );
buf ( n4384 , n416 );
buf ( n4385 , n1078 );
buf ( n4386 , n1671 );
buf ( n4387 , n994 );
buf ( n4388 , n1155 );
buf ( n4389 , n24 );
buf ( n4390 , n873 );
buf ( n4391 , n1173 );
buf ( n4392 , n666 );
buf ( n4393 , n608 );
buf ( n4394 , n37 );
buf ( n4395 , n1180 );
buf ( n4396 , n1168 );
buf ( n4397 , n48 );
buf ( n4398 , n256 );
buf ( n4399 , n1838 );
buf ( n4400 , n1861 );
buf ( n4401 , n1556 );
buf ( n4402 , n1284 );
buf ( n4403 , n472 );
buf ( n4404 , n1868 );
buf ( n4405 , n1715 );
buf ( n4406 , n1817 );
buf ( n4407 , n1743 );
buf ( n4408 , n1629 );
buf ( n4409 , n220 );
buf ( n4410 , n1716 );
buf ( n4411 , n586 );
buf ( n4412 , n1129 );
buf ( n4413 , n405 );
buf ( n4414 , n1683 );
buf ( n4415 , n833 );
buf ( n4416 , n1095 );
buf ( n4417 , n301 );
buf ( n4418 , n597 );
buf ( n4419 , n395 );
buf ( n4420 , n440 );
buf ( n4421 , n82 );
buf ( n4422 , n1314 );
buf ( n4423 , n1611 );
buf ( n4424 , n309 );
buf ( n4425 , n1899 );
buf ( n4426 , n81 );
buf ( n4427 , n1006 );
buf ( n4428 , n925 );
buf ( n4429 , n1814 );
buf ( n4430 , n739 );
buf ( n4431 , n1413 );
buf ( n4432 , n307 );
buf ( n4433 , n956 );
buf ( n4434 , n1004 );
buf ( n4435 , n529 );
buf ( n4436 , n1251 );
buf ( n4437 , n176 );
buf ( n4438 , n1364 );
buf ( n4439 , n1465 );
buf ( n4440 , n1728 );
buf ( n4441 , n362 );
buf ( n4442 , n1130 );
buf ( n4443 , n140 );
buf ( n4444 , n89 );
buf ( n4445 , n1025 );
buf ( n4446 , n632 );
buf ( n4447 , n1014 );
buf ( n4448 , n662 );
buf ( n4449 , n1096 );
buf ( n4450 , n641 );
buf ( n4451 , n1288 );
buf ( n4452 , n1975 );
buf ( n4453 , n60 );
buf ( n4454 , n1519 );
buf ( n4455 , n1998 );
buf ( n4456 , n1390 );
buf ( n4457 , n1506 );
buf ( n4458 , n1780 );
buf ( n4459 , n1412 );
buf ( n4460 , n154 );
buf ( n4461 , n1477 );
buf ( n4462 , n1072 );
buf ( n4463 , n1401 );
buf ( n4464 , n249 );
buf ( n4465 , n1091 );
buf ( n4466 , n1138 );
buf ( n4467 , n229 );
buf ( n4468 , n262 );
buf ( n4469 , n1543 );
buf ( n4470 , n984 );
buf ( n4471 , n415 );
buf ( n4472 , n1794 );
buf ( n4473 , n1175 );
buf ( n4474 , n1074 );
buf ( n4475 , n2015 );
buf ( n4476 , n1624 );
buf ( n4477 , n1242 );
buf ( n4478 , n1797 );
buf ( n4479 , n804 );
buf ( n4480 , n1508 );
buf ( n4481 , n145 );
buf ( n4482 , n1116 );
buf ( n4483 , n957 );
buf ( n4484 , n1375 );
buf ( n4485 , n1802 );
buf ( n4486 , n1420 );
buf ( n4487 , n1710 );
buf ( n4488 , n1942 );
buf ( n4489 , n178 );
buf ( n4490 , n1100 );
buf ( n4491 , n893 );
buf ( n4492 , n432 );
buf ( n4493 , n1448 );
buf ( n4494 , n1646 );
buf ( n4495 , n1694 );
buf ( n4496 , n375 );
buf ( n4497 , n1017 );
buf ( n4498 , n714 );
buf ( n4499 , n858 );
buf ( n4500 , n1117 );
buf ( n4501 , n785 );
buf ( n4502 , n450 );
buf ( n4503 , n328 );
buf ( n4504 , n659 );
buf ( n4505 , n1263 );
buf ( n4506 , n870 );
buf ( n4507 , n649 );
buf ( n4508 , n1285 );
buf ( n4509 , n1574 );
buf ( n4510 , n391 );
buf ( n4511 , n1232 );
buf ( n4512 , n1090 );
buf ( n4513 , n535 );
buf ( n4514 , n15 );
buf ( n4515 , n563 );
buf ( n4516 , n1149 );
buf ( n4517 , n1595 );
buf ( n4518 , n744 );
buf ( n4519 , n798 );
buf ( n4520 , n949 );
buf ( n4521 , n888 );
buf ( n4522 , n437 );
buf ( n4523 , n20 );
buf ( n4524 , n823 );
buf ( n4525 , n1900 );
buf ( n4526 , n195 );
buf ( n4527 , n772 );
buf ( n4528 , n304 );
buf ( n4529 , n1407 );
buf ( n4530 , n1395 );
buf ( n4531 , n2023 );
buf ( n4532 , n871 );
buf ( n4533 , n77 );
buf ( n4534 , n315 );
buf ( n4535 , n905 );
buf ( n4536 , n918 );
buf ( n4537 , n1593 );
buf ( n4538 , n406 );
buf ( n4539 , n506 );
buf ( n4540 , n4 );
buf ( n4541 , n1114 );
buf ( n4542 , n650 );
buf ( n4543 , n1967 );
buf ( n4544 , n424 );
buf ( n4545 , n1350 );
buf ( n4546 , n127 );
buf ( n4547 , n173 );
buf ( n4548 , n291 );
buf ( n4549 , n478 );
buf ( n4550 , n400 );
buf ( n4551 , n891 );
buf ( n4552 , n223 );
buf ( n4553 , n1793 );
buf ( n4554 , n1904 );
buf ( n4555 , n682 );
buf ( n4556 , n404 );
buf ( n4557 , n1619 );
buf ( n4558 , n1478 );
buf ( n4559 , n1709 );
buf ( n4560 , n466 );
buf ( n4561 , n1112 );
buf ( n4562 , n169 );
buf ( n4563 , n413 );
buf ( n4564 , n1514 );
buf ( n4565 , n99 );
buf ( n4566 , n560 );
buf ( n4567 , n1765 );
buf ( n4568 , n368 );
buf ( n4569 , n719 );
buf ( n4570 , n103 );
buf ( n4571 , n298 );
buf ( n4572 , n1596 );
buf ( n4573 , n617 );
buf ( n4574 , n710 );
buf ( n4575 , n686 );
buf ( n4576 , n1162 );
buf ( n4577 , n1876 );
buf ( n4578 , n435 );
buf ( n4579 , n98 );
buf ( n4580 , n1106 );
buf ( n4581 , n1222 );
buf ( n4582 , n55 );
buf ( n4583 , n1920 );
buf ( n4584 , n1191 );
buf ( n4585 , n265 );
buf ( n4586 , n507 );
buf ( n4587 , n1145 );
buf ( n4588 , n731 );
buf ( n4589 , n1172 );
buf ( n4590 , n584 );
buf ( n4591 , n1089 );
buf ( n4592 , n2026 );
buf ( n4593 , n57 );
buf ( n4594 , n587 );
buf ( n4595 , n1803 );
buf ( n4596 , n1071 );
buf ( n4597 , n1544 );
buf ( n4598 , n759 );
buf ( n4599 , n321 );
buf ( n4600 , n1795 );
buf ( n4601 , n732 );
buf ( n4602 , n908 );
buf ( n4603 , n627 );
buf ( n4604 , n1639 );
buf ( n4605 , n138 );
buf ( n4606 , n613 );
buf ( n4607 , n1688 );
buf ( n4608 , n342 );
buf ( n4609 , n1734 );
buf ( n4610 , n1919 );
buf ( n4611 , n2 );
buf ( n4612 , n377 );
buf ( n4613 , n1086 );
buf ( n4614 , n0 );
buf ( n4615 , n271 );
buf ( n4616 , n863 );
buf ( n4617 , n624 );
buf ( n4618 , n1905 );
buf ( n4619 , n648 );
buf ( n4620 , n829 );
buf ( n4621 , n1693 );
buf ( n4622 , n963 );
buf ( n4623 , n1818 );
buf ( n4624 , n944 );
buf ( n4625 , n1954 );
buf ( n4626 , n90 );
buf ( n4627 , n693 );
buf ( n4628 , n285 );
buf ( n4629 , n164 );
buf ( n4630 , n745 );
buf ( n4631 , n717 );
buf ( n4632 , n1827 );
buf ( n4633 , n456 );
buf ( n4634 , n923 );
buf ( n4635 , n654 );
buf ( n4636 , n1237 );
buf ( n4637 , n80 );
buf ( n4638 , n95 );
buf ( n4639 , n1557 );
buf ( n4640 , n2002 );
buf ( n4641 , n1087 );
buf ( n4642 , n474 );
buf ( n4643 , n626 );
buf ( n4644 , n247 );
buf ( n4645 , n545 );
buf ( n4646 , n112 );
buf ( n4647 , n1668 );
buf ( n4648 , n973 );
buf ( n4649 , n361 );
buf ( n4650 , n600 );
buf ( n4651 , n959 );
buf ( n4652 , n1859 );
buf ( n4653 , n1952 );
buf ( n4654 , n1307 );
buf ( n4655 , n227 );
buf ( n4656 , n1589 );
buf ( n4657 , n524 );
buf ( n4658 , n694 );
buf ( n4659 , n1971 );
buf ( n4660 , n1151 );
buf ( n4661 , n1978 );
buf ( n4662 , n1615 );
buf ( n4663 , n1893 );
buf ( n4664 , n1985 );
buf ( n4665 , n1053 );
buf ( n4666 , n157 );
buf ( n4667 , n997 );
buf ( n4668 , n1313 );
buf ( n4669 , n1842 );
buf ( n4670 , n1333 );
buf ( n4671 , n1181 );
buf ( n4672 , n230 );
buf ( n4673 , n928 );
buf ( n4674 , n1501 );
buf ( n4675 , n805 );
buf ( n4676 , n922 );
buf ( n4677 , n344 );
buf ( n4678 , n683 );
buf ( n4679 , n1620 );
buf ( n4680 , n786 );
buf ( n4681 , n889 );
buf ( n4682 , n299 );
buf ( n4683 , n747 );
buf ( n4684 , n282 );
buf ( n4685 , n768 );
buf ( n4686 , n467 );
buf ( n4687 , n1216 );
buf ( n4688 , n779 );
buf ( n4689 , n1272 );
buf ( n4690 , n1594 );
buf ( n4691 , n1064 );
buf ( n4692 , n1577 );
buf ( n4693 , n540 );
buf ( n4694 , n618 );
buf ( n4695 , n1599 );
buf ( n4696 , n565 );
buf ( n4697 , n360 );
buf ( n4698 , n645 );
buf ( n4699 , n1718 );
buf ( n4700 , n552 );
buf ( n4701 , n1653 );
buf ( n4702 , n1804 );
buf ( n4703 , n1505 );
buf ( n4704 , n1336 );
buf ( n4705 , n414 );
buf ( n4706 , n1335 );
buf ( n4707 , n1393 );
buf ( n4708 , n1680 );
buf ( n4709 , n1516 );
buf ( n4710 , n972 );
buf ( n4711 , n16 );
buf ( n4712 , n448 );
buf ( n4713 , n1354 );
buf ( n4714 , n1663 );
buf ( n4715 , n2020 );
buf ( n4716 , n1410 );
buf ( n4717 , n946 );
buf ( n4718 , n1641 );
buf ( n4719 , n1943 );
buf ( n4720 , n444 );
buf ( n4721 , n1186 );
buf ( n4722 , n26 );
buf ( n4723 , n384 );
buf ( n4724 , n36 );
buf ( n4725 , n856 );
buf ( n4726 , n548 );
buf ( n4727 , n1345 );
buf ( n4728 , n667 );
buf ( n4729 , n1136 );
buf ( n4730 , n302 );
buf ( n4731 , n567 );
buf ( n4732 , n1109 );
buf ( n4733 , n869 );
buf ( n4734 , n1060 );
buf ( n4735 , n1949 );
buf ( n4736 , n1982 );
buf ( n4737 , n836 );
buf ( n4738 , n1628 );
buf ( n4739 , n1849 );
buf ( n4740 , n673 );
buf ( n4741 , n1132 );
buf ( n4742 , n1264 );
buf ( n4743 , n1542 );
buf ( n4744 , n1127 );
buf ( n4745 , n1897 );
buf ( n4746 , n999 );
buf ( n4747 , n611 );
buf ( n4748 , n652 );
buf ( n4749 , n1559 );
buf ( n4750 , n1147 );
buf ( n4751 , n795 );
buf ( n4752 , n264 );
buf ( n4753 , n1343 );
buf ( n4754 , n163 );
buf ( n4755 , n799 );
buf ( n4756 , n1731 );
buf ( n4757 , n1361 );
buf ( n4758 , n892 );
buf ( n4759 , n27 );
buf ( n4760 , n570 );
buf ( n4761 , n1561 );
buf ( n4762 , n1926 );
buf ( n4763 , n834 );
buf ( n4764 , n238 );
buf ( n4765 , n1312 );
buf ( n4766 , n1647 );
buf ( n4767 , n203 );
buf ( n4768 , n532 );
buf ( n4769 , n1294 );
buf ( n4770 , n1602 );
buf ( n4771 , n1160 );
buf ( n4772 , n1576 );
buf ( n4773 , n787 );
buf ( n4774 , n46 );
buf ( n4775 , n1638 );
buf ( n4776 , n29 );
buf ( n4777 , n1070 );
buf ( n4778 , n1411 );
buf ( n4779 , n1115 );
buf ( n4780 , n1875 );
buf ( n4781 , n681 );
buf ( n4782 , n1040 );
buf ( n4783 , n1778 );
buf ( n4784 , n769 );
buf ( n4785 , n1640 );
buf ( n4786 , n1524 );
buf ( n4787 , n1029 );
buf ( n4788 , n609 );
buf ( n4789 , n1308 );
buf ( n4790 , n399 );
buf ( n4791 , n1931 );
buf ( n4792 , n475 );
buf ( n4793 , n1185 );
buf ( n4794 , n137 );
buf ( n4795 , n578 );
buf ( n4796 , n754 );
buf ( n4797 , n66 );
buf ( n4798 , n688 );
buf ( n4799 , n2034 );
buf ( n4800 , n1621 );
buf ( n4801 , n64 );
buf ( n4802 , n1084 );
buf ( n4803 , n30 );
buf ( n4804 , n1761 );
buf ( n4805 , n868 );
buf ( n4806 , n329 );
buf ( n4807 , n1691 );
buf ( n4808 , n907 );
buf ( n4809 , n1908 );
buf ( n4810 , n953 );
buf ( n4811 , n1582 );
buf ( n4812 , n1992 );
buf ( n4813 , n1337 );
buf ( n4814 , n1323 );
buf ( n4815 , n1224 );
buf ( n4816 , n1400 );
buf ( n4817 , n820 );
buf ( n4818 , n1244 );
buf ( n4819 , n1169 );
buf ( n4820 , n1083 );
buf ( n4821 , n909 );
buf ( n4822 , n837 );
buf ( n4823 , n912 );
buf ( n4824 , n185 );
buf ( n4825 , n1356 );
buf ( n4826 , n950 );
buf ( n4827 , n989 );
buf ( n4828 , n933 );
buf ( n4829 , n281 );
buf ( n4830 , n1651 );
buf ( n4831 , n1437 );
buf ( n4832 , n1417 );
buf ( n4833 , n568 );
buf ( n4834 , n1573 );
buf ( n4835 , n505 );
buf ( n4836 , n1566 );
buf ( n4837 , n885 );
buf ( n4838 , n1751 );
buf ( n4839 , n637 );
buf ( n4840 , n767 );
buf ( n4841 , n674 );
buf ( n4842 , n1484 );
buf ( n4843 , n54 );
buf ( n4844 , n748 );
buf ( n4845 , n1791 );
buf ( n4846 , n2000 );
buf ( n4847 , n358 );
buf ( n4848 , n251 );
buf ( n4849 , n1012 );
buf ( n4850 , n1275 );
buf ( n4851 , n1784 );
buf ( n4852 , n1930 );
buf ( n4853 , n41 );
buf ( n4854 , n1617 );
buf ( n4855 , n240 );
buf ( n4856 , n224 );
buf ( n4857 , n712 );
buf ( n4858 , n974 );
buf ( n4859 , n211 );
buf ( n4860 , n1669 );
buf ( n4861 , n896 );
buf ( n4862 , n373 );
buf ( n4863 , n1230 );
buf ( n4864 , n1179 );
buf ( n4865 , n1035 );
buf ( n4866 , n1445 );
buf ( n4867 , n431 );
buf ( n4868 , n557 );
buf ( n4869 , n287 );
buf ( n4870 , n1174 );
buf ( n4871 , n1892 );
buf ( n4872 , n487 );
buf ( n4873 , n2005 );
buf ( n4874 , n177 );
buf ( n4875 , n884 );
buf ( n4876 , n1874 );
buf ( n4877 , n1324 );
buf ( n4878 , n1605 );
buf ( n4879 , n1380 );
buf ( n4880 , n1247 );
buf ( n4881 , n1257 );
buf ( n4882 , n1613 );
buf ( n4883 , n1645 );
buf ( n4884 , n156 );
buf ( n4885 , n920 );
buf ( n4886 , n663 );
buf ( n4887 , n468 );
buf ( n4888 , n599 );
buf ( n4889 , n621 );
buf ( n4890 , n2006 );
buf ( n4891 , n1883 );
buf ( n4892 , n1065 );
buf ( n4893 , n802 );
buf ( n4894 , n1256 );
buf ( n4895 , n1196 );
buf ( n4896 , n1927 );
buf ( n4897 , n919 );
buf ( n4898 , n1889 );
buf ( n4899 , n1575 );
buf ( n4900 , n97 );
buf ( n4901 , n1122 );
buf ( n4902 , n148 );
buf ( n4903 , n1972 );
buf ( n4904 , n1409 );
buf ( n4905 , n958 );
buf ( n4906 , n336 );
buf ( n4907 , n261 );
buf ( n4908 , n1124 );
buf ( n4909 , n1002 );
buf ( n4910 , n326 );
buf ( n4911 , n1963 );
buf ( n4912 , n826 );
buf ( n4913 , n1187 );
buf ( n4914 , n1824 );
buf ( n4915 , n228 );
buf ( n4916 , n1032 );
buf ( n4917 , n1144 );
buf ( n4918 , n665 );
buf ( n4919 , n1276 );
buf ( n4920 , n1248 );
buf ( n4921 , n125 );
buf ( n4922 , n1279 );
buf ( n4923 , n1523 );
buf ( n4924 , n1742 );
buf ( n4925 , n1021 );
buf ( n4926 , n425 );
buf ( n4927 , n726 );
buf ( n4928 , n1073 );
buf ( n4929 , n1503 );
buf ( n4930 , n1098 );
buf ( n4931 , n350 );
buf ( n4932 , n1598 );
buf ( n4933 , n703 );
buf ( n4934 , n1882 );
buf ( n4935 , n865 );
buf ( n4936 , n1990 );
buf ( n4937 , n1567 );
buf ( n4938 , n1850 );
buf ( n4939 , n985 );
buf ( n4940 , n1923 );
buf ( n4941 , n2044 );
buf ( n4942 , n253 );
buf ( n4943 , n1746 );
buf ( n4944 , n45 );
buf ( n4945 , n766 );
buf ( n4946 , n180 );
buf ( n4947 , n1702 );
buf ( n4948 , n1808 );
buf ( n4949 , n1271 );
buf ( n4950 , n2025 );
buf ( n4951 , n1764 );
buf ( n4952 , n1282 );
buf ( n4953 , n1028 );
buf ( n4954 , n990 );
buf ( n4955 , n793 );
buf ( n4956 , n1103 );
buf ( n4957 , n1158 );
buf ( n4958 , n1555 );
buf ( n4959 , n1632 );
buf ( n4960 , n1042 );
buf ( n4961 , n252 );
buf ( n4962 , n1515 );
buf ( n4963 , n1648 );
buf ( n4964 , n455 );
buf ( n4965 , n794 );
buf ( n4966 , n490 );
buf ( n4967 , n1610 );
buf ( n4968 , n1270 );
buf ( n4969 , n353 );
buf ( n4970 , n462 );
buf ( n4971 , n1690 );
buf ( n4972 , n1022 );
buf ( n4973 , n341 );
buf ( n4974 , n1453 );
buf ( n4975 , n1907 );
buf ( n4976 , n704 );
buf ( n4977 , n550 );
buf ( n4978 , n107 );
buf ( n4979 , n1428 );
buf ( n4980 , n1399 );
buf ( n4981 , n1862 );
buf ( n4982 , n459 );
buf ( n4983 , n1212 );
buf ( n4984 , n1805 );
buf ( n4985 , n809 );
buf ( n4986 , n1890 );
buf ( n4987 , n186 );
buf ( n4988 , n1969 );
buf ( n4989 , n2039 );
buf ( n4990 , n1148 );
buf ( n4991 , n687 );
buf ( n4992 , n1939 );
buf ( n4993 , n1752 );
buf ( n4994 , n303 );
buf ( n4995 , n1363 );
buf ( n4996 , n1726 );
buf ( n4997 , n635 );
buf ( n4998 , n740 );
buf ( n4999 , n1649 );
buf ( n5000 , n758 );
buf ( n5001 , n1161 );
buf ( n5002 , n872 );
buf ( n5003 , n575 );
buf ( n5004 , n1054 );
buf ( n5005 , n1154 );
buf ( n5006 , n322 );
buf ( n5007 , n987 );
buf ( n5008 , n1534 );
buf ( n5009 , n49 );
buf ( n5010 , n1679 );
buf ( n5011 , n1750 );
buf ( n5012 , n308 );
buf ( n5013 , n862 );
buf ( n5014 , n124 );
buf ( n5015 , n1822 );
buf ( n5016 , n1261 );
buf ( n5017 , n825 );
buf ( n5018 , n1137 );
buf ( n5019 , n1475 );
buf ( n5020 , n1344 );
buf ( n5021 , n1366 );
buf ( n5022 , n1504 );
buf ( n5023 , n1913 );
buf ( n5024 , n878 );
buf ( n5025 , n516 );
buf ( n5026 , n470 );
buf ( n5027 , n843 );
buf ( n5028 , n1315 );
buf ( n5029 , n1706 );
buf ( n5030 , n616 );
buf ( n5031 , n698 );
buf ( n5032 , n554 );
buf ( n5033 , n842 );
buf ( n5034 , n723 );
buf ( n5035 , n1564 );
buf ( n5036 , n623 );
buf ( n5037 , n538 );
buf ( n5038 , n630 );
buf ( n5039 , n816 );
buf ( n5040 , n1790 );
buf ( n5041 , n1435 );
buf ( n5042 , n83 );
buf ( n5043 , n1675 );
buf ( n5044 , n1707 );
buf ( n5045 , n1848 );
buf ( n5046 , n2029 );
buf ( n5047 , n1066 );
buf ( n5048 , n280 );
buf ( n5049 , n1733 );
buf ( n5050 , n720 );
buf ( n5051 , n1281 );
buf ( n5052 , n857 );
buf ( n5053 , n995 );
buf ( n5054 , n1490 );
buf ( n5055 , n237 );
buf ( n5056 , n1183 );
buf ( n5057 , n1856 );
buf ( n5058 , n1806 );
buf ( n5059 , n234 );
buf ( n5060 , n316 );
buf ( n5061 , n756 );
buf ( n5062 , n1163 );
buf ( n5063 , n1461 );
buf ( n5064 , n160 );
buf ( n5065 , n564 );
buf ( n5066 , n469 );
buf ( n5067 , n942 );
buf ( n5068 , n2017 );
buf ( n5069 , n1552 );
buf ( n5070 , n1886 );
buf ( n5071 , n454 );
buf ( n5072 , n1832 );
buf ( n5073 , n1517 );
buf ( n5074 , n1820 );
buf ( n5075 , n607 );
buf ( n5076 , n1860 );
buf ( n5077 , n937 );
buf ( n5078 , n1879 );
buf ( n5079 , n774 );
buf ( n5080 , n386 );
buf ( n5081 , n1167 );
buf ( n5082 , n679 );
buf ( n5083 , n1799 );
buf ( n5084 , n518 );
buf ( n5085 , n1436 );
buf ( n5086 , n1870 );
buf ( n5087 , n479 );
buf ( n5088 , n651 );
buf ( n5089 , n1302 );
buf ( n5090 , n1771 );
buf ( n5091 , n1839 );
buf ( n5092 , n189 );
buf ( n5093 , n1269 );
buf ( n5094 , n1385 );
buf ( n5095 , n31 );
buf ( n5096 , n63 );
buf ( n5097 , n655 );
buf ( n5098 , n784 );
buf ( n5099 , n297 );
buf ( n5100 , n311 );
buf ( n5101 , n131 );
buf ( n5102 , n775 );
buf ( n5103 , n954 );
buf ( n5104 , n853 );
buf ( n5105 , n1146 );
buf ( n5106 , n977 );
buf ( n5107 , n1195 );
buf ( n5108 , n1553 );
buf ( n5109 , n491 );
buf ( n5110 , n201 );
buf ( n5111 , n434 );
buf ( n5112 , n1622 );
buf ( n5113 , n499 );
buf ( n5114 , n325 );
buf ( n5115 , n898 );
buf ( n5116 , n914 );
buf ( n5117 , n1165 );
buf ( n5118 , n992 );
buf ( n5119 , n1955 );
buf ( n5120 , n752 );
buf ( n5121 , n511 );
buf ( n5122 , n1929 );
buf ( n5123 , n1831 );
buf ( n5124 , n423 );
buf ( n5125 , n684 );
buf ( n5126 , n1705 );
buf ( n5127 , n2016 );
buf ( n5128 , n1944 );
buf ( n5129 , n1397 );
buf ( n5130 , n79 );
buf ( n5131 , n770 );
buf ( n5132 , n1038 );
buf ( n5133 , n1046 );
buf ( n5134 , n144 );
buf ( n5135 , n1736 );
buf ( n5136 , n270 );
buf ( n5137 , n1206 );
buf ( n5138 , n685 );
buf ( n5139 , n497 );
buf ( n5140 , n1441 );
buf ( n5141 , n939 );
buf ( n5142 , n536 );
buf ( n5143 , n1869 );
buf ( n5144 , n245 );
buf ( n5145 , n1968 );
buf ( n5146 , n840 );
buf ( n5147 , n815 );
buf ( n5148 , n1171 );
buf ( n5149 , n1398 );
buf ( n5150 , n970 );
buf ( n5151 , n827 );
buf ( n5152 , n1538 );
buf ( n5153 , n1775 );
buf ( n5154 , n1473 );
buf ( n5155 , n1215 );
buf ( n5156 , n1220 );
buf ( n5157 , n1976 );
buf ( n5158 , n1768 );
buf ( n5159 , n1614 );
buf ( n5160 , n1847 );
buf ( n5161 , n1601 );
buf ( n5162 , n1834 );
buf ( n5163 , n349 );
buf ( n5164 , n527 );
buf ( n5165 , n1684 );
buf ( n5166 , n278 );
buf ( n5167 , n1447 );
buf ( n5168 , n19 );
buf ( n5169 , n1654 );
buf ( n5170 , n689 );
buf ( n5171 , n1133 );
buf ( n5172 , n1851 );
buf ( n5173 , n737 );
buf ( n5174 , n1700 );
buf ( n5175 , n323 );
buf ( n5176 , n2037 );
buf ( n5177 , n846 );
buf ( n5178 , n1328 );
buf ( n5179 , n751 );
buf ( n5180 , n1346 );
buf ( n5181 , n1935 );
buf ( n5182 , n1604 );
buf ( n5183 , n1005 );
buf ( n5184 , n777 );
buf ( n5185 , n1933 );
buf ( n5186 , n1612 );
buf ( n5187 , n279 );
buf ( n5188 , n913 );
buf ( n5189 , n555 );
buf ( n5190 , n1906 );
buf ( n5191 , n1104 );
buf ( n5192 , n1320 );
buf ( n5193 , n644 );
buf ( n5194 , n1458 );
buf ( n5195 , n1854 );
buf ( n5196 , n1101 );
buf ( n5197 , n1884 );
buf ( n5198 , n596 );
buf ( n5199 , n473 );
buf ( n5200 , n13 );
buf ( n5201 , n1696 );
buf ( n5202 , n1527 );
buf ( n5203 , n1495 );
buf ( n5204 , n187 );
buf ( n5205 , n1075 );
buf ( n5206 , n1211 );
buf ( n5207 , n3 );
buf ( n5208 , n292 );
buf ( n5209 , n1426 );
buf ( n5210 , n938 );
buf ( n5211 , n2036 );
buf ( n5212 , n1030 );
buf ( n5213 , n1438 );
buf ( n5214 , n1379 );
buf ( n5215 , n874 );
buf ( n5216 , n1082 );
buf ( n5217 , n1063 );
buf ( n5218 , n646 );
buf ( n5219 , n883 );
buf ( n5220 , n796 );
buf ( n5221 , n142 );
buf ( n5222 , n168 );
buf ( n5223 , n1205 );
buf ( n5224 , n1973 );
buf ( n5225 , n706 );
buf ( n5226 , n975 );
buf ( n5227 , n1916 );
buf ( n5228 , n221 );
buf ( n5229 , n561 );
buf ( n5230 , n1581 );
buf ( n5231 , n1455 );
buf ( n5232 , n254 );
buf ( n5233 , n967 );
buf ( n5234 , n1033 );
buf ( n5235 , n243 );
buf ( n5236 , n396 );
buf ( n5237 , n1909 );
buf ( n5238 , n222 );
buf ( n5239 , n115 );
buf ( n5240 , n1056 );
buf ( n5241 , n1198 );
buf ( n5242 , n1801 );
buf ( n5243 , n813 );
buf ( n5244 , n1108 );
buf ( n5245 , n1487 );
buf ( n5246 , n1287 );
buf ( n5247 , n1499 );
buf ( n5248 , n409 );
buf ( n5249 , n1392 );
buf ( n5250 , n1828 );
buf ( n5251 , n1476 );
buf ( n5252 , n1088 );
buf ( n5253 , n1673 );
buf ( n5254 , n324 );
buf ( n5255 , n730 );
buf ( n5256 , n1770 );
buf ( n5257 , n1877 );
buf ( n5258 , n28 );
buf ( n5259 , n1485 );
buf ( n5260 , n113 );
buf ( n5261 , n1941 );
buf ( n5262 , n971 );
buf ( n5263 , n1946 );
buf ( n5264 , n494 );
buf ( n5265 , n512 );
buf ( n5266 , n2009 );
buf ( n5267 , n193 );
buf ( n5268 , n1011 );
buf ( n5269 , n2031 );
buf ( n5270 , n351 );
buf ( n5271 , n622 );
buf ( n5272 , n1097 );
buf ( n5273 , n1697 );
buf ( n5274 , n439 );
buf ( n5275 , n1368 );
buf ( n5276 , n1327 );
buf ( n5277 , n1483 );
buf ( n5278 , n911 );
buf ( n5279 , n210 );
buf ( n5280 , n383 );
buf ( n5281 , n1618 );
buf ( n5282 , n1027 );
buf ( n5283 , n1623 );
buf ( n5284 , n1304 );
buf ( n5285 , n2038 );
buf ( n5286 , n1661 );
buf ( n5287 , n129 );
buf ( n5288 , n445 );
buf ( n5289 , n130 );
buf ( n5290 , n1988 );
buf ( n5291 , n615 );
buf ( n5292 , n1178 );
buf ( n5293 , n5 );
buf ( n5294 , n1404 );
buf ( n5295 , n765 );
buf ( n5296 , n691 );
buf ( n5297 , n25 );
buf ( n5298 , n559 );
buf ( n5299 , n2014 );
buf ( n5300 , n1910 );
buf ( n5301 , n1965 );
buf ( n5302 , n1235 );
buf ( n5303 , n217 );
buf ( n5304 , n1451 );
buf ( n5305 , n38 );
buf ( n5306 , n1405 );
buf ( n5307 , n498 );
buf ( n5308 , n558 );
buf ( n5309 , n930 );
buf ( n5310 , n1472 );
buf ( n5311 , n1583 );
buf ( n5312 , n742 );
buf ( n5313 , n2021 );
buf ( n5314 , n1218 );
buf ( n5315 , n1260 );
buf ( n5316 , n1587 );
buf ( n5317 , n158 );
buf ( n5318 , n1763 );
buf ( n5319 , n1980 );
buf ( n5320 , n172 );
buf ( n5321 , n1600 );
buf ( n5322 , n1311 );
buf ( n5323 , n268 );
buf ( n5324 , n191 );
buf ( n5325 , n969 );
buf ( n5326 , n755 );
buf ( n5327 , n1188 );
buf ( n5328 , n22 );
buf ( n5329 , n1203 );
buf ( n5330 , n52 );
buf ( n5331 , n1134 );
buf ( n5332 , n1541 );
buf ( n5333 , n680 );
buf ( n5334 , n1317 );
buf ( n5335 , n1960 );
buf ( n5336 , n757 );
buf ( n5337 , n522 );
buf ( n5338 , n75 );
buf ( n5339 , n366 );
buf ( n5340 , n514 );
buf ( n5341 , n1330 );
buf ( n5342 , n1606 );
buf ( n5343 , n634 );
buf ( n5344 , n1219 );
buf ( n5345 , n1309 );
buf ( n5346 , n695 );
buf ( n5347 , n1321 );
buf ( n5348 , n690 );
buf ( n5349 , n492 );
buf ( n5350 , n1568 );
buf ( n5351 , n420 );
buf ( n5352 , n1585 );
buf ( n5353 , n1571 );
buf ( n5354 , n1938 );
buf ( n5355 , n904 );
buf ( n5356 , n1460 );
buf ( n5357 , n1249 );
buf ( n5358 , n830 );
buf ( n5359 , n763 );
buf ( n5360 , n2010 );
buf ( n5361 , n1894 );
buf ( n5362 , n998 );
buf ( n5363 , n225 );
buf ( n5364 , n1532 );
buf ( n5365 , n1800 );
buf ( n5366 , n1857 );
buf ( n5367 , n1956 );
buf ( n5368 , n70 );
buf ( n5369 , n1773 );
buf ( n5370 , n1781 );
buf ( n5371 , n387 );
buf ( n5372 , n1865 );
buf ( n5373 , n1911 );
buf ( n5374 , n800 );
buf ( n5375 , n159 );
buf ( n5376 , n1626 );
buf ( n5377 , n2030 );
buf ( n5378 , n831 );
buf ( n5379 , n1530 );
buf ( n5380 , n209 );
buf ( n5381 , n746 );
buf ( n5382 , n149 );
buf ( n5383 , n1105 );
buf ( n5384 , n465 );
buf ( n5385 , n40 );
buf ( n5386 , n1009 );
buf ( n5387 , n656 );
buf ( n5388 , n1373 );
buf ( n5389 , n1170 );
buf ( n5390 , n1914 );
buf ( n5391 , n1332 );
buf ( n5392 , n1951 );
buf ( n5393 , n1767 );
buf ( n5394 , n181 );
buf ( n5395 , n1974 );
buf ( n5396 , n146 );
buf ( n5397 , n7 );
buf ( n5398 , n1928 );
buf ( n5399 , n1762 );
buf ( n5400 , n1241 );
buf ( n5401 , n1227 );
buf ( n5402 , n1444 );
buf ( n5403 , n314 );
buf ( n5404 , n1043 );
buf ( n5405 , n629 );
buf ( n5406 , n901 );
buf ( n5407 , n1266 );
buf ( n5408 , n1226 );
buf ( n5409 , n633 );
buf ( n5410 , n595 );
buf ( n5411 , n231 );
buf ( n5412 , n1996 );
buf ( n5413 , n1048 );
buf ( n5414 , n783 );
buf ( n5415 , n284 );
buf ( n5416 , n1369 );
buf ( n5417 , n1550 );
buf ( n5418 , n789 );
buf ( n5419 , n1469 );
buf ( n5420 , n1948 );
buf ( n5421 , n283 );
buf ( n5422 , n1210 );
buf ( n5423 , n1560 );
buf ( n5424 , n708 );
buf ( n5425 , n390 );
buf ( n5426 , n1659 );
buf ( n5427 , n668 );
buf ( n5428 , n276 );
buf ( n5429 , n313 );
buf ( n5430 , n369 );
buf ( n5431 , n1255 );
buf ( n5432 , n675 );
buf ( n5433 , n610 );
buf ( n5434 , n1357 );
buf ( n5435 , n481 );
buf ( n5436 , n1819 );
buf ( n5437 , n1184 );
buf ( n5438 , n1486 );
buf ( n5439 , n219 );
buf ( n5440 , n1962 );
buf ( n5441 , n206 );
buf ( n5442 , n449 );
buf ( n5443 , n91 );
buf ( n5444 , n1807 );
buf ( n5445 , n1423 );
buf ( n5446 , n1482 );
buf ( n5447 , n1758 );
buf ( n5448 , n589 );
buf ( n5449 , n488 );
buf ( n5450 , n1010 );
buf ( n5451 , n86 );
buf ( n5452 , n643 );
buf ( n5453 , n1997 );
buf ( n5454 , n1725 );
buf ( n5455 , n402 );
buf ( n5456 , n152 );
buf ( n5457 , n1662 );
buf ( n5458 , n1331 );
buf ( n5459 , n1045 );
buf ( n5460 , n1026 );
buf ( n5461 , n1959 );
buf ( n5462 , n881 );
buf ( n5463 , n266 );
buf ( n5464 , n1633 );
buf ( n5465 , n1267 );
buf ( n5466 , n1316 );
buf ( n5467 , n371 );
buf ( n5468 , n312 );
buf ( n5469 , n32 );
buf ( n5470 , n1896 );
buf ( n5471 , n320 );
buf ( n5472 , n1007 );
buf ( n5473 , n1016 );
buf ( n5474 , n1391 );
buf ( n5475 , n806 );
buf ( n5476 , n1443 );
buf ( n5477 , n1657 );
buf ( n5478 , n1591 );
buf ( n5479 , n272 );
buf ( n5480 , n1347 );
buf ( n5481 , n1231 );
buf ( n5482 , n727 );
buf ( n5483 , n1748 );
buf ( n5484 , n1740 );
buf ( n5485 , n9 );
buf ( n5486 , n372 );
buf ( n5487 , n356 );
buf ( n5488 , n750 );
buf ( n5489 , n1755 );
buf ( n5490 , n1703 );
buf ( n5491 , n718 );
buf ( n5492 , n128 );
buf ( n5493 , n782 );
buf ( n5494 , n760 );
buf ( n5495 , n852 );
buf ( n5496 , n1578 );
buf ( n5497 , n1456 );
buf ( n5498 , n924 );
buf ( n5499 , n1425 );
buf ( n5500 , n1744 );
buf ( n5501 , n34 );
buf ( n5502 , n771 );
buf ( n5503 , n867 );
buf ( n5504 , n1421 );
buf ( n5505 , n246 );
buf ( n5506 , n1777 );
buf ( n5507 , n838 );
buf ( n5508 , n670 );
buf ( n5509 , n1511 );
buf ( n5510 , n1627 );
buf ( n5511 , n451 );
buf ( n5512 , n65 );
buf ( n5513 , n1239 );
buf ( n5514 , n1388 );
buf ( n5515 , n2027 );
buf ( n5516 , n51 );
buf ( n5517 , n2045 );
buf ( n5518 , n2028 );
buf ( n5519 , n71 );
buf ( n5520 , n1496 );
buf ( n5521 , n1650 );
buf ( n5522 , n1816 );
buf ( n5523 , n948 );
buf ( n5524 , n179 );
buf ( n5525 , n1670 );
buf ( n5526 , n1685 );
buf ( n5527 , n1554 );
buf ( n5528 , n170 );
buf ( n5529 , n1143 );
buf ( n5530 , n1403 );
buf ( n5531 , n471 );
buf ( n5532 , n510 );
buf ( n5533 , n1989 );
buf ( n5534 , n509 );
buf ( n5535 , n1166 );
buf ( n5536 , n875 );
buf ( n5537 , n1432 );
buf ( n5538 , n374 );
buf ( n5539 , n202 );
buf ( n5540 , n12 );
buf ( n5541 , n389 );
buf ( n5542 , n161 );
buf ( n5543 , n531 );
buf ( n5544 , n263 );
buf ( n5545 , n1994 );
buf ( n5546 , n1253 );
buf ( n5547 , n260 );
buf ( n5548 , n2003 );
buf ( n5549 , n1776 );
buf ( n5550 , n1194 );
buf ( n5551 , n150 );
buf ( n5552 , n1551 );
buf ( n5553 , n539 );
buf ( n5554 , n503 );
buf ( n5555 , n743 );
buf ( n5556 , n1000 );
buf ( n5557 , n1835 );
buf ( n5558 , n1666 );
buf ( n5559 , n1296 );
buf ( n5560 , n736 );
buf ( n5561 , n734 );
buf ( n5562 , n346 );
buf ( n5563 , n847 );
buf ( n5564 , n1470 );
buf ( n5565 , n1440 );
buf ( n5566 , n716 );
buf ( n5567 , n1200 );
buf ( n5568 , n1643 );
buf ( n5569 , n1433 );
buf ( n5570 , n715 );
buf ( n5571 , n1031 );
buf ( n5572 , n1262 );
buf ( n5573 , n1430 );
buf ( n5574 , n408 );
buf ( n5575 , n1457 );
buf ( n5576 , n625 );
buf ( n5577 , n583 );
buf ( n5578 , n947 );
buf ( n5579 , n1494 );
buf ( n5580 , n1424 );
buf ( n5581 , n1068 );
buf ( n5582 , n2042 );
buf ( n5583 , n338 );
buf ( n5584 , n73 );
buf ( n5585 , n1286 );
buf ( n5586 , n190 );
buf ( n5587 , n53 );
buf ( n5588 , n701 );
buf ( n5589 , n1358 );
buf ( n5590 , n1565 );
buf ( n5591 , n812 );
buf ( n5592 , n821 );
buf ( n5593 , n1152 );
buf ( n5594 , n677 );
buf ( n5595 , n1001 );
buf ( n5596 , n588 );
buf ( n5597 , n1342 );
buf ( n5598 , n1754 );
buf ( n5599 , n631 );
buf ( n5600 , n484 );
buf ( n5601 , n1759 );
buf ( n5602 , n1153 );
buf ( n5603 , n628 );
buf ( n5604 , n35 );
buf ( n5605 , n556 );
buf ( n5606 , n1872 );
buf ( n5607 , n647 );
buf ( n5608 , n1672 );
buf ( n5609 , n1841 );
buf ( n5610 , n579 );
buf ( n5611 , n155 );
buf ( n5612 , n817 );
buf ( n5613 , n69 );
buf ( n5614 , n382 );
buf ( n5615 , n1984 );
buf ( n5616 , n241 );
buf ( n5617 , n1699 );
buf ( n5618 , n1783 );
buf ( n5619 , n355 );
buf ( n5620 , n1291 );
buf ( n5621 , n255 );
buf ( n5622 , n1603 );
buf ( n5623 , n1289 );
buf ( n5624 , n1635 );
buf ( n5625 , n1003 );
buf ( n5626 , n1389 );
buf ( n5627 , n464 );
buf ( n5628 , n544 );
buf ( n5629 , n11 );
buf ( n5630 , n707 );
buf ( n5631 , n855 );
buf ( n5632 , n171 );
buf ( n5633 , n676 );
buf ( n5634 , n2008 );
buf ( n5635 , n1844 );
buf ( n5636 , n257 );
buf ( n5637 , n359 );
buf ( n5638 , n397 );
buf ( n5639 , n1076 );
buf ( n5640 , n1348 );
buf ( n5641 , n489 );
buf ( n5642 , n101 );
buf ( n5643 , n1686 );
buf ( n5644 , n1724 );
buf ( n5645 , n121 );
buf ( n5646 , n370 );
buf ( n5647 , n1416 );
buf ( n5648 , n1549 );
buf ( n5649 , n962 );
buf ( n5650 , n398 );
buf ( n5651 , n1940 );
buf ( n5652 , n1676 );
buf ( n5653 , n702 );
buf ( n5654 , n378 );
buf ( n5655 , n213 );
buf ( n5656 , n1526 );
buf ( n5657 , n401 );
buf ( n5658 , n1131 );
buf ( n5659 , n286 );
buf ( n5660 , n657 );
buf ( n5661 , n1536 );
buf ( n5662 , n1120 );
buf ( n5663 , n678 );
buf ( n5664 , n376 );
buf ( n5665 , n1836 );
buf ( n5666 , n1548 );
buf ( n5667 , n1991 );
buf ( n5668 , n1427 );
buf ( n5669 , n1189 );
buf ( n5670 , n1925 );
buf ( n5671 , n175 );
buf ( n5672 , n1921 );
buf ( n5673 , n339 );
buf ( n5674 , n1535 );
buf ( n5675 , n811 );
buf ( n5676 , n493 );
buf ( n5677 , n343 );
buf ( n5678 , n58 );
buf ( n5679 , n1020 );
buf ( n5680 , n1584 );
buf ( n5681 , n880 );
buf ( n5682 , n1298 );
buf ( n5683 , n1637 );
buf ( n5684 , n1902 );
buf ( n5685 , n1418 );
buf ( n5686 , n1008 );
buf ( n5687 , n2018 );
buf ( n5688 , n886 );
buf ( n5689 , n394 );
buf ( n5690 , n672 );
buf ( n5691 , n964 );
buf ( n5692 , n986 );
buf ( n5693 , n1058 );
buf ( n5694 , n248 );
buf ( n5695 , n864 );
buf ( n5696 , n100 );
buf ( n5697 , n1782 );
buf ( n5698 , n1636 );
buf ( n5699 , n1371 );
buf ( n5700 , n1749 );
buf ( n5701 , n1864 );
buf ( n5702 , n790 );
buf ( n5703 , n310 );
buf ( n5704 , n978 );
buf ( n5705 , n738 );
buf ( n5706 , n1537 );
buf ( n5707 , n94 );
buf ( n5708 , n1190 );
buf ( n5709 , n1277 );
buf ( n5710 , n1319 );
buf ( n5711 , n43 );
buf ( n5712 , n845 );
buf ( n5713 , n1280 );
buf ( n5714 , n501 );
buf ( n5715 , n1431 );
buf ( n5716 , n1840 );
buf ( n5717 , n860 );
buf ( n5718 , n340 );
buf ( n5719 , n1936 );
buf ( n5720 , n1677 );
buf ( n5721 , n1209 );
buf ( n5722 , n126 );
buf ( n5723 , n1310 );
buf ( n5724 , n569 );
buf ( n5725 , n388 );
buf ( n5726 , n1121 );
buf ( n5727 , n109 );
buf ( n5728 , n1446 );
buf ( n5729 , n1047 );
buf ( n5730 , n1439 );
buf ( n5731 , n1737 );
buf ( n5732 , n1608 );
buf ( n5733 , n577 );
buf ( n5734 , n277 );
buf ( n5735 , n585 );
buf ( n5736 , n357 );
buf ( n5737 , n1871 );
buf ( n5738 , n562 );
buf ( n5739 , n1717 );
buf ( n5740 , n983 );
buf ( n5741 , n1059 );
buf ( n5742 , n940 );
buf ( n5743 , n194 );
buf ( n5744 , n929 );
buf ( n5745 , n1995 );
buf ( n5746 , n1359 );
buf ( n5747 , n1182 );
buf ( n5748 , n899 );
buf ( n5749 , n441 );
buf ( n5750 , n705 );
buf ( n5751 , n1987 );
buf ( n5752 , n1837 );
buf ( n5753 , n788 );
buf ( n5754 , n1245 );
buf ( n5755 , n1233 );
buf ( n5756 , n819 );
buf ( n5757 , n887 );
buf ( n5758 , n1341 );
buf ( n5759 , n1292 );
buf ( n5760 , n1062 );
buf ( n5761 , n1099 );
buf ( n5762 , n1081 );
buf ( n5763 , n1917 );
buf ( n5764 , n1502 );
buf ( n5765 , n1102 );
buf ( n5766 , n1177 );
buf ( n5767 , n430 );
buf ( n5768 , n1957 );
buf ( n5769 , n2022 );
buf ( n5770 , n902 );
buf ( n5771 , n1452 );
buf ( n5772 , n352 );
buf ( n5773 , n1204 );
buf ( n5774 , n1786 );
buf ( n5775 , n1492 );
buf ( n5776 , n327 );
buf ( n5777 , n1708 );
buf ( n5778 , n182 );
buf ( n5779 , n1377 );
buf ( n5780 , n1509 );
buf ( n5781 , n1562 );
buf ( n5782 , n848 );
buf ( n5783 , n1125 );
buf ( n5784 , n367 );
buf ( n5785 , n204 );
buf ( n5786 , n1164 );
buf ( n5787 , n218 );
buf ( n5788 , n991 );
buf ( n5789 , n1986 );
buf ( n5790 , n1774 );
buf ( n5791 , n594 );
buf ( n5792 , n446 );
buf ( n5793 , n1981 );
buf ( n5794 , n1258 );
buf ( n5795 , n122 );
buf ( n5796 , n84 );
buf ( n5797 , n700 );
buf ( n5798 , n188 );
buf ( n5799 , n476 );
buf ( n5800 , n935 );
buf ( n5801 , n1903 );
buf ( n5802 , n952 );
buf ( n5803 , n290 );
buf ( n5804 , n120 );
buf ( n5805 , n571 );
buf ( n5806 , n580 );
buf ( n5807 , n1507 );
buf ( n5808 , n433 );
buf ( n5809 , n1353 );
buf ( n5810 , n890 );
buf ( n5811 , n300 );
buf ( n5812 , n111 );
buf ( n5813 , n1642 );
buf ( n5814 , n335 );
buf ( n5815 , n92 );
buf ( n5816 , n232 );
buf ( n5817 , n1351 );
buf ( n5818 , n1067 );
buf ( n5819 , n1880 );
buf ( n5820 , n1192 );
buf ( n5821 , n18 );
buf ( n5822 , n136 );
buf ( n5823 , n123 );
buf ( n5824 , n1422 );
buf ( n5825 , n1217 );
buf ( n5826 , n44 );
buf ( n5827 , n866 );
buf ( n5828 , n1964 );
buf ( n5829 , n296 );
buf ( n5830 , n1922 );
buf ( n5831 , n1510 );
buf ( n5832 , n379 );
buf ( n5833 , n106 );
buf ( n5834 , n295 );
buf ( n5835 , n638 );
buf ( n5836 , n1881 );
buf ( n5837 , n818 );
buf ( n5838 , n1468 );
buf ( n5839 , n363 );
buf ( n5840 , n1118 );
buf ( n5841 , n1660 );
buf ( n5842 , n722 );
buf ( n5843 , n521 );
buf ( n5844 , n1340 );
buf ( n5845 , n1093 );
buf ( n5846 , n2011 );
buf ( n5847 , n1 );
buf ( n5848 , n1825 );
buf ( n5849 , n1891 );
buf ( n5850 , n192 );
buf ( n5851 , n1999 );
buf ( n5852 , n791 );
buf ( n5853 , n764 );
buf ( n5854 , n1701 );
buf ( n5855 , n761 );
buf ( n5856 , n1572 );
buf ( n5857 , n293 );
buf ( n5858 , n1498 );
buf ( n5859 , n119 );
buf ( n5860 , n151 );
buf ( n5861 , n1077 );
buf ( n5862 , n1934 );
buf ( n5863 , n380 );
buf ( n5864 , n581 );
buf ( n5865 , n733 );
buf ( n5866 , n496 );
buf ( n5867 , n966 );
buf ( n5868 , n418 );
buf ( n5869 , n1547 );
buf ( n5870 , n525 );
buf ( n5871 , n258 );
buf ( n5872 , n927 );
buf ( n5873 , n1208 );
buf ( n5874 , n508 );
buf ( n5875 , n1429 );
buf ( n5876 , n1199 );
buf ( n5877 , n797 );
buf ( n5878 , n951 );
buf ( n5879 , n102 );
buf ( n5880 , n134 );
buf ( n5881 , n1958 );
buf ( n5882 , n1057 );
buf ( n5883 , n955 );
buf ( n5884 , n1156 );
buf ( n5885 , n56 );
buf ( n5886 , n1692 );
buf ( n5887 , n822 );
buf ( n5888 , n1352 );
buf ( n5889 , n1464 );
buf ( n5890 , n735 );
buf ( n5891 , n410 );
buf ( n5892 , n1811 );
buf ( n5893 , n980 );
buf ( n5894 , n1714 );
buf ( n5895 , n523 );
buf ( n5896 , n1349 );
buf ( n5897 , n915 );
buf ( n5898 , n692 );
buf ( n5899 , n941 );
buf ( n5900 , n1809 );
buf ( n5901 , n1631 );
buf ( n5902 , n614 );
buf ( n5903 , n1887 );
buf ( n5904 , n1735 );
buf ( n5905 , n1520 );
buf ( n5906 , n483 );
buf ( n5907 , n33 );
buf ( n5908 , n877 );
buf ( n5909 , n1853 );
buf ( n5910 , n882 );
buf ( n5911 , n39 );
buf ( n5912 , n1024 );
buf ( n5913 , n658 );
buf ( n5914 , n244 );
buf ( n5915 , n1326 );
buf ( n5916 , n574 );
buf ( n5917 , n162 );
buf ( n5918 , n417 );
buf ( n5919 , n1682 );
buf ( n5920 , n1760 );
buf ( n5921 , n1961 );
buf ( n5922 , n1609 );
buf ( n5923 , n214 );
buf ( n5924 , n781 );
buf ( n5925 , n542 );
buf ( n5926 , n553 );
buf ( n5927 , n1630 );
buf ( n5928 , n590 );
buf ( n5929 , n1322 );
buf ( n5930 , n835 );
buf ( n5931 , n226 );
buf ( n5932 , n861 );
buf ( n5933 , n495 );
buf ( n5934 , n1013 );
buf ( n5935 , n669 );
buf ( n5936 , n289 );
buf ( n5937 , n1681 );
buf ( n5938 , n216 );
buf ( n5939 , n1415 );
buf ( n5940 , n895 );
buf ( n5941 , n500 );
buf ( n5942 , n1732 );
buf ( n5943 , n839 );
buf ( n5944 , n438 );
buf ( n5945 , n330 );
buf ( n5946 , n1250 );
buf ( n5947 , n1381 );
buf ( n5948 , n1018 );
buf ( n5949 , n233 );
buf ( n5950 , n88 );
buf ( n5951 , n551 );
buf ( n5952 , n832 );
buf ( n5953 , n916 );
buf ( n5954 , n1141 );
buf ( n5955 , n879 );
buf ( n5956 , n1597 );
buf ( n5957 , n1474 );
buf ( n5958 , n117 );
buf ( n5959 , n1396 );
buf ( n5960 , n598 );
buf ( n5961 , n1779 );
buf ( n5962 , n1197 );
buf ( n5963 , n392 );
buf ( n5964 , n844 );
buf ( n5965 , n165 );
buf ( n5966 , n988 );
buf ( n5967 , n1689 );
buf ( n5968 , n1159 );
buf ( n5969 , n1273 );
buf ( n5970 , n945 );
buf ( n5971 , n546 );
buf ( n5972 , n2040 );
buf ( n5973 , n1528 );
buf ( n5974 , n1766 );
buf ( n5975 , n1529 );
buf ( n5976 , n96 );
buf ( n5977 , n1953 );
buf ( n5978 , n1918 );
buf ( n5979 , n572 );
buf ( n5980 , n1295 );
buf ( n5981 , n2004 );
buf ( n5982 , n965 );
buf ( n5983 , n566 );
buf ( n5984 , n1376 );
buf ( n5985 , n1225 );
buf ( n5986 , n1207 );
buf ( n5987 , n664 );
buf ( n5988 , n147 );
buf ( n5989 , n1665 );
buf ( n5990 , n345 );
buf ( n5991 , n943 );
buf ( n5992 , n1757 );
buf ( n5993 , n2032 );
buf ( n5994 , n721 );
buf ( n5995 , n294 );
buf ( n5996 , n183 );
buf ( n5997 , n1932 );
buf ( n5998 , n773 );
buf ( n5999 , n1055 );
buf ( n6000 , n1213 );
buf ( n6001 , n1829 );
buf ( n6002 , n1655 );
buf ( n6003 , n894 );
buf ( n6004 , n1810 );
buf ( n6005 , n1355 );
buf ( n6006 , n337 );
buf ( n6007 , n1945 );
buf ( n6008 , n1924 );
buf ( n6009 , n926 );
buf ( n6010 , n639 );
buf ( n6011 , n1569 );
buf ( n6012 , n653 );
buf ( n6013 , n1656 );
buf ( n6014 , n1382 );
buf ( n6015 , n74 );
buf ( n6016 , n1329 );
buf ( n6017 , n463 );
buf ( n6018 , n2033 );
buf ( n6019 , n582 );
buf ( n6020 , n68 );
buf ( n6021 , n776 );
buf ( n6022 , n1019 );
buf ( n6023 , n2024 );
buf ( n6024 , n1434 );
buf ( n6025 , n259 );
buf ( n6026 , n1738 );
buf ( n6027 , n1318 );
buf ( n6028 , n198 );
buf ( n6029 , n808 );
buf ( n6030 , n699 );
buf ( n6031 , n1497 );
buf ( n6032 , n167 );
buf ( n6033 , n517 );
buf ( n6034 , n982 );
buf ( n6035 , n110 );
buf ( n6036 , n2007 );
buf ( n6037 , n1044 );
buf ( n6038 , n429 );
buf ( n6039 , n576 );
buf ( n6040 , n528 );
buf ( n6041 , n47 );
buf ( n6042 , n1378 );
buf ( n6043 , n235 );
buf ( n6044 , n427 );
buf ( n6045 , n436 );
buf ( n6046 , n828 );
buf ( n6047 , n1798 );
buf ( n6048 , n1747 );
buf ( n6049 , n859 );
buf ( n6050 , n1202 );
buf ( n6051 , n1833 );
buf ( n6052 , n1365 );
buf ( n6053 , n1788 );
buf ( n6054 , n1796 );
buf ( n6055 , n976 );
buf ( n6056 , n1150 );
buf ( n6057 , n306 );
buf ( n6058 , n741 );
buf ( n6059 , n778 );
buf ( n6060 , n1252 );
buf ( n6061 , n1852 );
buf ( n6062 , n93 );
buf ( n6063 , n1229 );
buf ( n6064 , n1080 );
buf ( n6065 , n1142 );
buf ( n6066 , n810 );
buf ( n6067 , n407 );
buf ( n6068 , n593 );
buf ( n6069 , n934 );
buf ( n6070 , n1372 );
buf ( n6071 , n1545 );
buf ( n6072 , n1687 );
buf ( n6073 , n526 );
buf ( n6074 , n1489 );
buf ( n6075 , n1283 );
buf ( n6076 , n1049 );
buf ( n6077 , n14 );
buf ( n6078 , n1036 );
buf ( n6079 , n697 );
buf ( n6080 , n1481 );
buf ( n6081 , n174 );
buf ( n6082 , n591 );
buf ( n6083 , n334 );
buf ( n6084 , n458 );
buf ( n6085 , n1471 );
buf ( n6086 , n184 );
buf ( n6087 , n724 );
buf ( n6088 , n1254 );
buf ( n6089 , n979 );
buf ( n6090 , n1821 );
buf ( n6091 , n936 );
buf ( n6092 , n199 );
buf ( n6093 , n1094 );
buf ( n6094 , n573 );
buf ( n6095 , n1858 );
buf ( n6096 , n1383 );
buf ( n6097 , n305 );
buf ( n6098 , n385 );
buf ( n6099 , n592 );
buf ( n6100 , n749 );
buf ( n6101 , n1845 );
buf ( n6102 , n1823 );
buf ( n6103 , n2001 );
buf ( n6104 , n541 );
buf ( n6105 , n1236 );
buf ( n6106 , n1723 );
buf ( n6107 , n1367 );
buf ( n6108 , n1558 );
buf ( n6109 , n897 );
buf ( n6110 , n1402 );
buf ( n6111 , n1176 );
buf ( n6112 , n996 );
buf ( n6113 , n1712 );
buf ( n6114 , n1278 );
buf ( n6115 , n1488 );
buf ( n6116 , n762 );
buf ( n6117 , n347 );
buf ( n6118 , n1667 );
buf ( n6119 , n1644 );
buf ( n6120 , n1467 );
buf ( n6121 , n1843 );
buf ( n6122 , n1238 );
buf ( n6123 , n502 );
buf ( n6124 , n1873 );
buf ( n6125 , n1157 );
buf ( n6126 , n671 );
buf ( n6127 , n1135 );
buf ( n6128 , n2046 );
buf ( n6129 , n729 );
buf ( n6130 , n1293 );
buf ( n6131 , n1128 );
buf ( n6132 , n1338 );
buf ( n6133 , n961 );
buf ( n6134 , n274 );
buf ( n6135 , n1720 );
buf ( n6136 , n1730 );
buf ( n6137 , n851 );
buf ( n6138 , n8 );
buf ( n6139 , n1039 );
buf ( n6140 , n1041 );
buf ( n6141 , n960 );
buf ( n6142 , n1394 );
buf ( n6143 , n1370 );
buf ( n6144 , n660 );
buf ( n6145 , n642 );
buf ( n6146 , n1698 );
buf ( n6147 , n1111 );
buf ( n6148 , n59 );
buf ( n6149 , n547 );
buf ( n6150 , n5126 );
buf ( n6151 , n5127 );
or ( n6152 , n6150 , n6151 );
buf ( n6153 , n5128 );
or ( n6154 , n6152 , n6153 );
buf ( n6155 , n5129 );
or ( n6156 , n6154 , n6155 );
buf ( n6157 , n5130 );
or ( n6158 , n6156 , n6157 );
buf ( n6159 , n5131 );
or ( n6160 , n6158 , n6159 );
buf ( n6161 , n5132 );
or ( n6162 , n6160 , n6161 );
buf ( n6163 , n5133 );
or ( n6164 , n6162 , n6163 );
buf ( n6165 , n5134 );
or ( n6166 , n6164 , n6165 );
buf ( n6167 , n5135 );
or ( n6168 , n6166 , n6167 );
buf ( n6169 , n5136 );
or ( n6170 , n6168 , n6169 );
buf ( n6171 , n5137 );
or ( n6172 , n6170 , n6171 );
buf ( n6173 , n5138 );
or ( n6174 , n6172 , n6173 );
buf ( n6175 , n5139 );
or ( n6176 , n6174 , n6175 );
buf ( n6177 , n5140 );
or ( n6178 , n6176 , n6177 );
buf ( n6179 , n5141 );
or ( n6180 , n6178 , n6179 );
buf ( n6181 , n5142 );
or ( n6182 , n6180 , n6181 );
buf ( n6183 , n5143 );
or ( n6184 , n6182 , n6183 );
buf ( n6185 , n5144 );
or ( n6186 , n6184 , n6185 );
buf ( n6187 , n5145 );
or ( n6188 , n6186 , n6187 );
buf ( n6189 , n5146 );
or ( n6190 , n6188 , n6189 );
buf ( n6191 , n5147 );
or ( n6192 , n6190 , n6191 );
buf ( n6193 , n5148 );
or ( n6194 , n6192 , n6193 );
buf ( n6195 , n5149 );
or ( n6196 , n6194 , n6195 );
buf ( n6197 , n5150 );
or ( n6198 , n6196 , n6197 );
buf ( n6199 , n5151 );
or ( n6200 , n6198 , n6199 );
buf ( n6201 , n5152 );
or ( n6202 , n6200 , n6201 );
buf ( n6203 , n5153 );
or ( n6204 , n6202 , n6203 );
buf ( n6205 , n5154 );
or ( n6206 , n6204 , n6205 );
buf ( n6207 , n5155 );
or ( n6208 , n6206 , n6207 );
buf ( n6209 , n5156 );
or ( n6210 , n6208 , n6209 );
buf ( n6211 , n5157 );
or ( n6212 , n6210 , n6211 );
buf ( n6213 , n5158 );
or ( n6214 , n6212 , n6213 );
buf ( n6215 , n5159 );
or ( n6216 , n6214 , n6215 );
buf ( n6217 , n5160 );
or ( n6218 , n6216 , n6217 );
buf ( n6219 , n5161 );
or ( n6220 , n6218 , n6219 );
buf ( n6221 , n5162 );
or ( n6222 , n6220 , n6221 );
buf ( n6223 , n5163 );
or ( n6224 , n6222 , n6223 );
buf ( n6225 , n5164 );
or ( n6226 , n6224 , n6225 );
buf ( n6227 , n5165 );
or ( n6228 , n6226 , n6227 );
buf ( n6229 , n5166 );
or ( n6230 , n6228 , n6229 );
buf ( n6231 , n5167 );
or ( n6232 , n6230 , n6231 );
buf ( n6233 , n5168 );
or ( n6234 , n6232 , n6233 );
buf ( n6235 , n5169 );
or ( n6236 , n6234 , n6235 );
buf ( n6237 , n5170 );
or ( n6238 , n6236 , n6237 );
buf ( n6239 , n5171 );
or ( n6240 , n6238 , n6239 );
buf ( n6241 , n5172 );
or ( n6242 , n6240 , n6241 );
buf ( n6243 , n5173 );
or ( n6244 , n6242 , n6243 );
buf ( n6245 , n5174 );
or ( n6246 , n6244 , n6245 );
buf ( n6247 , n5175 );
or ( n6248 , n6246 , n6247 );
buf ( n6249 , n5176 );
or ( n6250 , n6248 , n6249 );
buf ( n6251 , n5177 );
or ( n6252 , n6250 , n6251 );
buf ( n6253 , n5178 );
or ( n6254 , n6252 , n6253 );
buf ( n6255 , n5179 );
or ( n6256 , n6254 , n6255 );
buf ( n6257 , n5180 );
or ( n6258 , n6256 , n6257 );
buf ( n6259 , n5181 );
or ( n6260 , n6258 , n6259 );
buf ( n6261 , n5182 );
or ( n6262 , n6260 , n6261 );
buf ( n6263 , n5183 );
or ( n6264 , n6262 , n6263 );
buf ( n6265 , n5184 );
or ( n6266 , n6264 , n6265 );
buf ( n6267 , n5185 );
or ( n6268 , n6266 , n6267 );
buf ( n6269 , n5186 );
or ( n6270 , n6268 , n6269 );
buf ( n6271 , n5187 );
or ( n6272 , n6270 , n6271 );
buf ( n6273 , n5188 );
or ( n6274 , n6272 , n6273 );
buf ( n6275 , n5189 );
or ( n6276 , n6274 , n6275 );
buf ( n6277 , n5190 );
or ( n6278 , n6276 , n6277 );
buf ( n6279 , n5191 );
or ( n6280 , n6278 , n6279 );
buf ( n6281 , n5192 );
or ( n6282 , n6280 , n6281 );
buf ( n6283 , n5193 );
or ( n6284 , n6282 , n6283 );
buf ( n6285 , n5194 );
or ( n6286 , n6284 , n6285 );
buf ( n6287 , n5195 );
or ( n6288 , n6286 , n6287 );
buf ( n6289 , n5196 );
or ( n6290 , n6288 , n6289 );
buf ( n6291 , n5197 );
or ( n6292 , n6290 , n6291 );
buf ( n6293 , n5198 );
or ( n6294 , n6292 , n6293 );
buf ( n6295 , n5199 );
or ( n6296 , n6294 , n6295 );
buf ( n6297 , n5200 );
or ( n6298 , n6296 , n6297 );
buf ( n6299 , n5201 );
or ( n6300 , n6298 , n6299 );
buf ( n6301 , n5202 );
or ( n6302 , n6300 , n6301 );
buf ( n6303 , n5203 );
or ( n6304 , n6302 , n6303 );
buf ( n6305 , n5204 );
or ( n6306 , n6304 , n6305 );
buf ( n6307 , n5205 );
or ( n6308 , n6306 , n6307 );
buf ( n6309 , n5206 );
or ( n6310 , n6308 , n6309 );
buf ( n6311 , n5207 );
or ( n6312 , n6310 , n6311 );
buf ( n6313 , n5208 );
or ( n6314 , n6312 , n6313 );
buf ( n6315 , n5209 );
or ( n6316 , n6314 , n6315 );
buf ( n6317 , n5210 );
or ( n6318 , n6316 , n6317 );
buf ( n6319 , n5211 );
or ( n6320 , n6318 , n6319 );
buf ( n6321 , n5212 );
or ( n6322 , n6320 , n6321 );
buf ( n6323 , n5213 );
or ( n6324 , n6322 , n6323 );
buf ( n6325 , n5214 );
or ( n6326 , n6324 , n6325 );
buf ( n6327 , n5215 );
or ( n6328 , n6326 , n6327 );
buf ( n6329 , n5216 );
or ( n6330 , n6328 , n6329 );
buf ( n6331 , n5217 );
or ( n6332 , n6330 , n6331 );
buf ( n6333 , n5218 );
or ( n6334 , n6332 , n6333 );
buf ( n6335 , n5219 );
or ( n6336 , n6334 , n6335 );
buf ( n6337 , n5220 );
or ( n6338 , n6336 , n6337 );
buf ( n6339 , n5221 );
or ( n6340 , n6338 , n6339 );
buf ( n6341 , n5222 );
or ( n6342 , n6340 , n6341 );
buf ( n6343 , n5223 );
or ( n6344 , n6342 , n6343 );
buf ( n6345 , n5224 );
or ( n6346 , n6344 , n6345 );
buf ( n6347 , n5225 );
or ( n6348 , n6346 , n6347 );
buf ( n6349 , n5226 );
or ( n6350 , n6348 , n6349 );
buf ( n6351 , n5227 );
or ( n6352 , n6350 , n6351 );
buf ( n6353 , n5228 );
or ( n6354 , n6352 , n6353 );
buf ( n6355 , n5229 );
or ( n6356 , n6354 , n6355 );
buf ( n6357 , n5230 );
or ( n6358 , n6356 , n6357 );
buf ( n6359 , n5231 );
or ( n6360 , n6358 , n6359 );
buf ( n6361 , n5232 );
or ( n6362 , n6360 , n6361 );
buf ( n6363 , n5233 );
or ( n6364 , n6362 , n6363 );
buf ( n6365 , n5234 );
or ( n6366 , n6364 , n6365 );
buf ( n6367 , n5235 );
or ( n6368 , n6366 , n6367 );
buf ( n6369 , n5236 );
or ( n6370 , n6368 , n6369 );
buf ( n6371 , n5237 );
or ( n6372 , n6370 , n6371 );
buf ( n6373 , n5238 );
or ( n6374 , n6372 , n6373 );
buf ( n6375 , n5239 );
or ( n6376 , n6374 , n6375 );
buf ( n6377 , n5240 );
or ( n6378 , n6376 , n6377 );
buf ( n6379 , n5241 );
or ( n6380 , n6378 , n6379 );
buf ( n6381 , n5242 );
or ( n6382 , n6380 , n6381 );
buf ( n6383 , n5243 );
or ( n6384 , n6382 , n6383 );
buf ( n6385 , n5244 );
or ( n6386 , n6384 , n6385 );
buf ( n6387 , n5245 );
or ( n6388 , n6386 , n6387 );
buf ( n6389 , n5246 );
or ( n6390 , n6388 , n6389 );
buf ( n6391 , n5247 );
or ( n6392 , n6390 , n6391 );
buf ( n6393 , n5248 );
or ( n6394 , n6392 , n6393 );
buf ( n6395 , n5249 );
or ( n6396 , n6394 , n6395 );
buf ( n6397 , n5250 );
or ( n6398 , n6396 , n6397 );
buf ( n6399 , n5251 );
or ( n6400 , n6398 , n6399 );
buf ( n6401 , n5252 );
or ( n6402 , n6400 , n6401 );
buf ( n6403 , n5253 );
or ( n6404 , n6402 , n6403 );
buf ( n6405 , n5254 );
or ( n6406 , n6404 , n6405 );
buf ( n6407 , n5255 );
or ( n6408 , n6406 , n6407 );
buf ( n6409 , n5256 );
or ( n6410 , n6408 , n6409 );
buf ( n6411 , n5257 );
or ( n6412 , n6410 , n6411 );
buf ( n6413 , n5258 );
or ( n6414 , n6412 , n6413 );
buf ( n6415 , n5259 );
or ( n6416 , n6414 , n6415 );
buf ( n6417 , n5260 );
or ( n6418 , n6416 , n6417 );
buf ( n6419 , n5261 );
or ( n6420 , n6418 , n6419 );
buf ( n6421 , n5262 );
or ( n6422 , n6420 , n6421 );
buf ( n6423 , n5263 );
or ( n6424 , n6422 , n6423 );
buf ( n6425 , n5264 );
or ( n6426 , n6424 , n6425 );
buf ( n6427 , n5265 );
or ( n6428 , n6426 , n6427 );
buf ( n6429 , n5266 );
or ( n6430 , n6428 , n6429 );
buf ( n6431 , n5267 );
or ( n6432 , n6430 , n6431 );
buf ( n6433 , n5268 );
or ( n6434 , n6432 , n6433 );
buf ( n6435 , n5269 );
or ( n6436 , n6434 , n6435 );
buf ( n6437 , n5270 );
or ( n6438 , n6436 , n6437 );
buf ( n6439 , n5271 );
or ( n6440 , n6438 , n6439 );
buf ( n6441 , n5272 );
or ( n6442 , n6440 , n6441 );
buf ( n6443 , n5273 );
or ( n6444 , n6442 , n6443 );
buf ( n6445 , n5274 );
or ( n6446 , n6444 , n6445 );
buf ( n6447 , n5275 );
or ( n6448 , n6446 , n6447 );
buf ( n6449 , n5276 );
or ( n6450 , n6448 , n6449 );
buf ( n6451 , n5277 );
or ( n6452 , n6450 , n6451 );
buf ( n6453 , n5278 );
or ( n6454 , n6452 , n6453 );
buf ( n6455 , n5279 );
or ( n6456 , n6454 , n6455 );
buf ( n6457 , n5280 );
or ( n6458 , n6456 , n6457 );
buf ( n6459 , n5281 );
or ( n6460 , n6458 , n6459 );
buf ( n6461 , n5282 );
or ( n6462 , n6460 , n6461 );
buf ( n6463 , n5283 );
or ( n6464 , n6462 , n6463 );
buf ( n6465 , n5284 );
or ( n6466 , n6464 , n6465 );
buf ( n6467 , n5285 );
or ( n6468 , n6466 , n6467 );
buf ( n6469 , n5286 );
or ( n6470 , n6468 , n6469 );
buf ( n6471 , n5287 );
or ( n6472 , n6470 , n6471 );
buf ( n6473 , n5288 );
or ( n6474 , n6472 , n6473 );
buf ( n6475 , n5289 );
or ( n6476 , n6474 , n6475 );
buf ( n6477 , n5290 );
or ( n6478 , n6476 , n6477 );
buf ( n6479 , n5291 );
or ( n6480 , n6478 , n6479 );
buf ( n6481 , n5292 );
or ( n6482 , n6480 , n6481 );
buf ( n6483 , n5293 );
or ( n6484 , n6482 , n6483 );
buf ( n6485 , n5294 );
or ( n6486 , n6484 , n6485 );
buf ( n6487 , n5295 );
or ( n6488 , n6486 , n6487 );
buf ( n6489 , n5296 );
or ( n6490 , n6488 , n6489 );
buf ( n6491 , n5297 );
or ( n6492 , n6490 , n6491 );
buf ( n6493 , n5298 );
or ( n6494 , n6492 , n6493 );
buf ( n6495 , n5299 );
or ( n6496 , n6494 , n6495 );
buf ( n6497 , n5300 );
or ( n6498 , n6496 , n6497 );
buf ( n6499 , n5301 );
or ( n6500 , n6498 , n6499 );
buf ( n6501 , n5302 );
or ( n6502 , n6500 , n6501 );
buf ( n6503 , n5303 );
or ( n6504 , n6502 , n6503 );
buf ( n6505 , n5304 );
or ( n6506 , n6504 , n6505 );
buf ( n6507 , n5305 );
or ( n6508 , n6506 , n6507 );
buf ( n6509 , n5306 );
or ( n6510 , n6508 , n6509 );
buf ( n6511 , n5307 );
or ( n6512 , n6510 , n6511 );
buf ( n6513 , n5308 );
or ( n6514 , n6512 , n6513 );
buf ( n6515 , n5309 );
or ( n6516 , n6514 , n6515 );
buf ( n6517 , n5310 );
or ( n6518 , n6516 , n6517 );
buf ( n6519 , n5311 );
or ( n6520 , n6518 , n6519 );
buf ( n6521 , n5312 );
or ( n6522 , n6520 , n6521 );
buf ( n6523 , n5313 );
or ( n6524 , n6522 , n6523 );
buf ( n6525 , n5314 );
or ( n6526 , n6524 , n6525 );
buf ( n6527 , n5315 );
or ( n6528 , n6526 , n6527 );
buf ( n6529 , n5316 );
or ( n6530 , n6528 , n6529 );
buf ( n6531 , n5317 );
or ( n6532 , n6530 , n6531 );
buf ( n6533 , n5318 );
or ( n6534 , n6532 , n6533 );
buf ( n6535 , n5319 );
or ( n6536 , n6534 , n6535 );
buf ( n6537 , n5320 );
or ( n6538 , n6536 , n6537 );
buf ( n6539 , n5321 );
or ( n6540 , n6538 , n6539 );
buf ( n6541 , n5322 );
or ( n6542 , n6540 , n6541 );
buf ( n6543 , n5323 );
or ( n6544 , n6542 , n6543 );
buf ( n6545 , n5324 );
or ( n6546 , n6544 , n6545 );
buf ( n6547 , n5325 );
or ( n6548 , n6546 , n6547 );
buf ( n6549 , n5326 );
or ( n6550 , n6548 , n6549 );
buf ( n6551 , n5327 );
or ( n6552 , n6550 , n6551 );
buf ( n6553 , n5328 );
or ( n6554 , n6552 , n6553 );
buf ( n6555 , n5329 );
or ( n6556 , n6554 , n6555 );
buf ( n6557 , n5330 );
or ( n6558 , n6556 , n6557 );
buf ( n6559 , n5331 );
or ( n6560 , n6558 , n6559 );
buf ( n6561 , n5332 );
or ( n6562 , n6560 , n6561 );
buf ( n6563 , n5333 );
or ( n6564 , n6562 , n6563 );
buf ( n6565 , n5334 );
or ( n6566 , n6564 , n6565 );
buf ( n6567 , n5335 );
or ( n6568 , n6566 , n6567 );
buf ( n6569 , n5336 );
or ( n6570 , n6568 , n6569 );
buf ( n6571 , n5337 );
or ( n6572 , n6570 , n6571 );
buf ( n6573 , n5338 );
or ( n6574 , n6572 , n6573 );
buf ( n6575 , n5339 );
or ( n6576 , n6574 , n6575 );
buf ( n6577 , n5340 );
or ( n6578 , n6576 , n6577 );
buf ( n6579 , n5341 );
or ( n6580 , n6578 , n6579 );
buf ( n6581 , n5342 );
or ( n6582 , n6580 , n6581 );
buf ( n6583 , n5343 );
or ( n6584 , n6582 , n6583 );
buf ( n6585 , n5344 );
or ( n6586 , n6584 , n6585 );
buf ( n6587 , n5345 );
or ( n6588 , n6586 , n6587 );
buf ( n6589 , n5346 );
or ( n6590 , n6588 , n6589 );
buf ( n6591 , n5347 );
or ( n6592 , n6590 , n6591 );
buf ( n6593 , n5348 );
or ( n6594 , n6592 , n6593 );
buf ( n6595 , n5349 );
or ( n6596 , n6594 , n6595 );
buf ( n6597 , n5350 );
or ( n6598 , n6596 , n6597 );
buf ( n6599 , n5351 );
or ( n6600 , n6598 , n6599 );
buf ( n6601 , n5352 );
or ( n6602 , n6600 , n6601 );
buf ( n6603 , n5353 );
or ( n6604 , n6602 , n6603 );
buf ( n6605 , n5354 );
or ( n6606 , n6604 , n6605 );
buf ( n6607 , n5355 );
or ( n6608 , n6606 , n6607 );
buf ( n6609 , n5356 );
or ( n6610 , n6608 , n6609 );
buf ( n6611 , n5357 );
or ( n6612 , n6610 , n6611 );
buf ( n6613 , n5358 );
or ( n6614 , n6612 , n6613 );
buf ( n6615 , n5359 );
or ( n6616 , n6614 , n6615 );
buf ( n6617 , n5360 );
or ( n6618 , n6616 , n6617 );
buf ( n6619 , n5361 );
or ( n6620 , n6618 , n6619 );
buf ( n6621 , n5362 );
or ( n6622 , n6620 , n6621 );
buf ( n6623 , n5363 );
or ( n6624 , n6622 , n6623 );
buf ( n6625 , n5364 );
or ( n6626 , n6624 , n6625 );
buf ( n6627 , n5365 );
or ( n6628 , n6626 , n6627 );
buf ( n6629 , n5366 );
or ( n6630 , n6628 , n6629 );
buf ( n6631 , n5367 );
or ( n6632 , n6630 , n6631 );
buf ( n6633 , n5368 );
or ( n6634 , n6632 , n6633 );
buf ( n6635 , n5369 );
or ( n6636 , n6634 , n6635 );
buf ( n6637 , n5370 );
or ( n6638 , n6636 , n6637 );
buf ( n6639 , n5371 );
or ( n6640 , n6638 , n6639 );
buf ( n6641 , n5372 );
or ( n6642 , n6640 , n6641 );
buf ( n6643 , n5373 );
or ( n6644 , n6642 , n6643 );
buf ( n6645 , n5374 );
or ( n6646 , n6644 , n6645 );
buf ( n6647 , n5375 );
or ( n6648 , n6646 , n6647 );
buf ( n6649 , n5376 );
or ( n6650 , n6648 , n6649 );
buf ( n6651 , n5377 );
or ( n6652 , n6650 , n6651 );
buf ( n6653 , n5378 );
or ( n6654 , n6652 , n6653 );
buf ( n6655 , n5379 );
or ( n6656 , n6654 , n6655 );
buf ( n6657 , n5380 );
or ( n6658 , n6656 , n6657 );
buf ( n6659 , n5381 );
or ( n6660 , n6658 , n6659 );
buf ( n6661 , n5382 );
or ( n6662 , n6660 , n6661 );
buf ( n6663 , n5383 );
or ( n6664 , n6662 , n6663 );
buf ( n6665 , n5384 );
or ( n6666 , n6664 , n6665 );
buf ( n6667 , n5385 );
or ( n6668 , n6666 , n6667 );
buf ( n6669 , n5386 );
or ( n6670 , n6668 , n6669 );
buf ( n6671 , n5387 );
or ( n6672 , n6670 , n6671 );
buf ( n6673 , n5388 );
or ( n6674 , n6672 , n6673 );
buf ( n6675 , n5389 );
or ( n6676 , n6674 , n6675 );
buf ( n6677 , n5390 );
or ( n6678 , n6676 , n6677 );
buf ( n6679 , n5391 );
or ( n6680 , n6678 , n6679 );
buf ( n6681 , n5392 );
or ( n6682 , n6680 , n6681 );
buf ( n6683 , n5393 );
or ( n6684 , n6682 , n6683 );
buf ( n6685 , n5394 );
or ( n6686 , n6684 , n6685 );
buf ( n6687 , n5395 );
or ( n6688 , n6686 , n6687 );
buf ( n6689 , n5396 );
or ( n6690 , n6688 , n6689 );
buf ( n6691 , n5397 );
or ( n6692 , n6690 , n6691 );
buf ( n6693 , n5398 );
or ( n6694 , n6692 , n6693 );
buf ( n6695 , n5399 );
or ( n6696 , n6694 , n6695 );
buf ( n6697 , n5400 );
or ( n6698 , n6696 , n6697 );
buf ( n6699 , n5401 );
or ( n6700 , n6698 , n6699 );
buf ( n6701 , n5402 );
or ( n6702 , n6700 , n6701 );
buf ( n6703 , n5403 );
or ( n6704 , n6702 , n6703 );
buf ( n6705 , n5404 );
or ( n6706 , n6704 , n6705 );
buf ( n6707 , n5405 );
or ( n6708 , n6706 , n6707 );
buf ( n6709 , n5406 );
or ( n6710 , n6708 , n6709 );
buf ( n6711 , n5407 );
or ( n6712 , n6710 , n6711 );
buf ( n6713 , n5408 );
or ( n6714 , n6712 , n6713 );
buf ( n6715 , n5409 );
or ( n6716 , n6714 , n6715 );
buf ( n6717 , n5410 );
or ( n6718 , n6716 , n6717 );
buf ( n6719 , n5411 );
or ( n6720 , n6718 , n6719 );
buf ( n6721 , n5412 );
or ( n6722 , n6720 , n6721 );
buf ( n6723 , n5413 );
or ( n6724 , n6722 , n6723 );
buf ( n6725 , n5414 );
or ( n6726 , n6724 , n6725 );
buf ( n6727 , n5415 );
or ( n6728 , n6726 , n6727 );
buf ( n6729 , n5416 );
or ( n6730 , n6728 , n6729 );
buf ( n6731 , n5417 );
or ( n6732 , n6730 , n6731 );
buf ( n6733 , n5418 );
or ( n6734 , n6732 , n6733 );
buf ( n6735 , n5419 );
or ( n6736 , n6734 , n6735 );
buf ( n6737 , n5420 );
or ( n6738 , n6736 , n6737 );
buf ( n6739 , n5421 );
or ( n6740 , n6738 , n6739 );
buf ( n6741 , n5422 );
or ( n6742 , n6740 , n6741 );
buf ( n6743 , n5423 );
or ( n6744 , n6742 , n6743 );
buf ( n6745 , n5424 );
or ( n6746 , n6744 , n6745 );
buf ( n6747 , n5425 );
or ( n6748 , n6746 , n6747 );
buf ( n6749 , n5426 );
or ( n6750 , n6748 , n6749 );
buf ( n6751 , n5427 );
or ( n6752 , n6750 , n6751 );
buf ( n6753 , n5428 );
or ( n6754 , n6752 , n6753 );
buf ( n6755 , n5429 );
or ( n6756 , n6754 , n6755 );
buf ( n6757 , n5430 );
or ( n6758 , n6756 , n6757 );
buf ( n6759 , n5431 );
or ( n6760 , n6758 , n6759 );
buf ( n6761 , n5432 );
or ( n6762 , n6760 , n6761 );
buf ( n6763 , n5433 );
or ( n6764 , n6762 , n6763 );
buf ( n6765 , n5434 );
or ( n6766 , n6764 , n6765 );
buf ( n6767 , n5435 );
or ( n6768 , n6766 , n6767 );
buf ( n6769 , n5436 );
or ( n6770 , n6768 , n6769 );
buf ( n6771 , n5437 );
or ( n6772 , n6770 , n6771 );
buf ( n6773 , n5438 );
or ( n6774 , n6772 , n6773 );
buf ( n6775 , n5439 );
or ( n6776 , n6774 , n6775 );
buf ( n6777 , n5440 );
or ( n6778 , n6776 , n6777 );
buf ( n6779 , n5441 );
or ( n6780 , n6778 , n6779 );
buf ( n6781 , n5442 );
or ( n6782 , n6780 , n6781 );
buf ( n6783 , n5443 );
or ( n6784 , n6782 , n6783 );
buf ( n6785 , n5444 );
or ( n6786 , n6784 , n6785 );
buf ( n6787 , n5445 );
or ( n6788 , n6786 , n6787 );
buf ( n6789 , n5446 );
or ( n6790 , n6788 , n6789 );
buf ( n6791 , n5447 );
or ( n6792 , n6790 , n6791 );
buf ( n6793 , n5448 );
or ( n6794 , n6792 , n6793 );
buf ( n6795 , n5449 );
or ( n6796 , n6794 , n6795 );
buf ( n6797 , n5450 );
or ( n6798 , n6796 , n6797 );
buf ( n6799 , n5451 );
or ( n6800 , n6798 , n6799 );
buf ( n6801 , n5452 );
or ( n6802 , n6800 , n6801 );
buf ( n6803 , n5453 );
or ( n6804 , n6802 , n6803 );
buf ( n6805 , n5454 );
or ( n6806 , n6804 , n6805 );
buf ( n6807 , n5455 );
or ( n6808 , n6806 , n6807 );
buf ( n6809 , n5456 );
or ( n6810 , n6808 , n6809 );
buf ( n6811 , n5457 );
or ( n6812 , n6810 , n6811 );
buf ( n6813 , n5458 );
or ( n6814 , n6812 , n6813 );
buf ( n6815 , n5459 );
or ( n6816 , n6814 , n6815 );
buf ( n6817 , n5460 );
or ( n6818 , n6816 , n6817 );
buf ( n6819 , n5461 );
or ( n6820 , n6818 , n6819 );
buf ( n6821 , n5462 );
or ( n6822 , n6820 , n6821 );
buf ( n6823 , n5463 );
or ( n6824 , n6822 , n6823 );
buf ( n6825 , n5464 );
or ( n6826 , n6824 , n6825 );
buf ( n6827 , n5465 );
or ( n6828 , n6826 , n6827 );
buf ( n6829 , n5466 );
or ( n6830 , n6828 , n6829 );
buf ( n6831 , n5467 );
or ( n6832 , n6830 , n6831 );
buf ( n6833 , n5468 );
or ( n6834 , n6832 , n6833 );
buf ( n6835 , n5469 );
or ( n6836 , n6834 , n6835 );
buf ( n6837 , n5470 );
or ( n6838 , n6836 , n6837 );
buf ( n6839 , n5471 );
or ( n6840 , n6838 , n6839 );
buf ( n6841 , n5472 );
or ( n6842 , n6840 , n6841 );
buf ( n6843 , n5473 );
or ( n6844 , n6842 , n6843 );
buf ( n6845 , n5474 );
or ( n6846 , n6844 , n6845 );
buf ( n6847 , n5475 );
or ( n6848 , n6846 , n6847 );
buf ( n6849 , n5476 );
or ( n6850 , n6848 , n6849 );
buf ( n6851 , n5477 );
or ( n6852 , n6850 , n6851 );
buf ( n6853 , n5478 );
or ( n6854 , n6852 , n6853 );
buf ( n6855 , n5479 );
or ( n6856 , n6854 , n6855 );
buf ( n6857 , n5480 );
or ( n6858 , n6856 , n6857 );
buf ( n6859 , n5481 );
or ( n6860 , n6858 , n6859 );
buf ( n6861 , n5482 );
or ( n6862 , n6860 , n6861 );
buf ( n6863 , n5483 );
or ( n6864 , n6862 , n6863 );
buf ( n6865 , n5484 );
or ( n6866 , n6864 , n6865 );
buf ( n6867 , n5485 );
or ( n6868 , n6866 , n6867 );
buf ( n6869 , n5486 );
or ( n6870 , n6868 , n6869 );
buf ( n6871 , n5487 );
or ( n6872 , n6870 , n6871 );
buf ( n6873 , n5488 );
or ( n6874 , n6872 , n6873 );
buf ( n6875 , n5489 );
or ( n6876 , n6874 , n6875 );
buf ( n6877 , n5490 );
or ( n6878 , n6876 , n6877 );
buf ( n6879 , n5491 );
or ( n6880 , n6878 , n6879 );
buf ( n6881 , n5492 );
or ( n6882 , n6880 , n6881 );
buf ( n6883 , n5493 );
or ( n6884 , n6882 , n6883 );
buf ( n6885 , n5494 );
or ( n6886 , n6884 , n6885 );
buf ( n6887 , n5495 );
or ( n6888 , n6886 , n6887 );
buf ( n6889 , n5496 );
or ( n6890 , n6888 , n6889 );
buf ( n6891 , n5497 );
or ( n6892 , n6890 , n6891 );
buf ( n6893 , n5498 );
or ( n6894 , n6892 , n6893 );
buf ( n6895 , n5499 );
or ( n6896 , n6894 , n6895 );
buf ( n6897 , n5500 );
or ( n6898 , n6896 , n6897 );
buf ( n6899 , n5501 );
or ( n6900 , n6898 , n6899 );
buf ( n6901 , n5502 );
or ( n6902 , n6900 , n6901 );
buf ( n6903 , n5503 );
or ( n6904 , n6902 , n6903 );
buf ( n6905 , n5504 );
or ( n6906 , n6904 , n6905 );
buf ( n6907 , n5505 );
or ( n6908 , n6906 , n6907 );
buf ( n6909 , n5506 );
or ( n6910 , n6908 , n6909 );
buf ( n6911 , n5507 );
or ( n6912 , n6910 , n6911 );
buf ( n6913 , n5508 );
or ( n6914 , n6912 , n6913 );
buf ( n6915 , n5509 );
or ( n6916 , n6914 , n6915 );
buf ( n6917 , n5510 );
or ( n6918 , n6916 , n6917 );
buf ( n6919 , n5511 );
or ( n6920 , n6918 , n6919 );
buf ( n6921 , n5512 );
or ( n6922 , n6920 , n6921 );
buf ( n6923 , n5513 );
or ( n6924 , n6922 , n6923 );
buf ( n6925 , n5514 );
or ( n6926 , n6924 , n6925 );
buf ( n6927 , n5515 );
or ( n6928 , n6926 , n6927 );
buf ( n6929 , n5516 );
or ( n6930 , n6928 , n6929 );
buf ( n6931 , n5517 );
or ( n6932 , n6930 , n6931 );
buf ( n6933 , n5518 );
or ( n6934 , n6932 , n6933 );
buf ( n6935 , n5519 );
or ( n6936 , n6934 , n6935 );
buf ( n6937 , n5520 );
or ( n6938 , n6936 , n6937 );
buf ( n6939 , n5521 );
or ( n6940 , n6938 , n6939 );
buf ( n6941 , n5522 );
or ( n6942 , n6940 , n6941 );
buf ( n6943 , n5523 );
or ( n6944 , n6942 , n6943 );
buf ( n6945 , n5524 );
or ( n6946 , n6944 , n6945 );
buf ( n6947 , n5525 );
or ( n6948 , n6946 , n6947 );
buf ( n6949 , n5526 );
or ( n6950 , n6948 , n6949 );
buf ( n6951 , n5527 );
or ( n6952 , n6950 , n6951 );
buf ( n6953 , n5528 );
or ( n6954 , n6952 , n6953 );
buf ( n6955 , n5529 );
or ( n6956 , n6954 , n6955 );
buf ( n6957 , n5530 );
or ( n6958 , n6956 , n6957 );
buf ( n6959 , n5531 );
or ( n6960 , n6958 , n6959 );
buf ( n6961 , n5532 );
or ( n6962 , n6960 , n6961 );
buf ( n6963 , n5533 );
or ( n6964 , n6962 , n6963 );
buf ( n6965 , n5534 );
or ( n6966 , n6964 , n6965 );
buf ( n6967 , n5535 );
or ( n6968 , n6966 , n6967 );
buf ( n6969 , n5536 );
or ( n6970 , n6968 , n6969 );
buf ( n6971 , n5537 );
or ( n6972 , n6970 , n6971 );
buf ( n6973 , n5538 );
or ( n6974 , n6972 , n6973 );
buf ( n6975 , n5539 );
or ( n6976 , n6974 , n6975 );
buf ( n6977 , n5540 );
or ( n6978 , n6976 , n6977 );
buf ( n6979 , n5541 );
or ( n6980 , n6978 , n6979 );
buf ( n6981 , n5542 );
or ( n6982 , n6980 , n6981 );
buf ( n6983 , n5543 );
or ( n6984 , n6982 , n6983 );
buf ( n6985 , n5544 );
or ( n6986 , n6984 , n6985 );
buf ( n6987 , n5545 );
or ( n6988 , n6986 , n6987 );
buf ( n6989 , n5546 );
or ( n6990 , n6988 , n6989 );
buf ( n6991 , n5547 );
or ( n6992 , n6990 , n6991 );
buf ( n6993 , n5548 );
or ( n6994 , n6992 , n6993 );
buf ( n6995 , n5549 );
or ( n6996 , n6994 , n6995 );
buf ( n6997 , n5550 );
or ( n6998 , n6996 , n6997 );
buf ( n6999 , n5551 );
or ( n7000 , n6998 , n6999 );
buf ( n7001 , n5552 );
or ( n7002 , n7000 , n7001 );
buf ( n7003 , n5553 );
or ( n7004 , n7002 , n7003 );
buf ( n7005 , n5554 );
or ( n7006 , n7004 , n7005 );
buf ( n7007 , n5555 );
or ( n7008 , n7006 , n7007 );
buf ( n7009 , n5556 );
or ( n7010 , n7008 , n7009 );
buf ( n7011 , n5557 );
or ( n7012 , n7010 , n7011 );
buf ( n7013 , n5558 );
or ( n7014 , n7012 , n7013 );
buf ( n7015 , n5559 );
or ( n7016 , n7014 , n7015 );
buf ( n7017 , n5560 );
or ( n7018 , n7016 , n7017 );
buf ( n7019 , n5561 );
or ( n7020 , n7018 , n7019 );
buf ( n7021 , n5562 );
or ( n7022 , n7020 , n7021 );
buf ( n7023 , n5563 );
or ( n7024 , n7022 , n7023 );
buf ( n7025 , n5564 );
or ( n7026 , n7024 , n7025 );
buf ( n7027 , n5565 );
or ( n7028 , n7026 , n7027 );
buf ( n7029 , n5566 );
or ( n7030 , n7028 , n7029 );
buf ( n7031 , n5567 );
or ( n7032 , n7030 , n7031 );
buf ( n7033 , n5568 );
or ( n7034 , n7032 , n7033 );
buf ( n7035 , n5569 );
or ( n7036 , n7034 , n7035 );
buf ( n7037 , n5570 );
or ( n7038 , n7036 , n7037 );
buf ( n7039 , n5571 );
or ( n7040 , n7038 , n7039 );
buf ( n7041 , n5572 );
or ( n7042 , n7040 , n7041 );
buf ( n7043 , n5573 );
or ( n7044 , n7042 , n7043 );
buf ( n7045 , n5574 );
or ( n7046 , n7044 , n7045 );
buf ( n7047 , n5575 );
or ( n7048 , n7046 , n7047 );
buf ( n7049 , n5576 );
or ( n7050 , n7048 , n7049 );
buf ( n7051 , n5577 );
or ( n7052 , n7050 , n7051 );
buf ( n7053 , n5578 );
or ( n7054 , n7052 , n7053 );
buf ( n7055 , n5579 );
or ( n7056 , n7054 , n7055 );
buf ( n7057 , n5580 );
or ( n7058 , n7056 , n7057 );
buf ( n7059 , n5581 );
or ( n7060 , n7058 , n7059 );
buf ( n7061 , n5582 );
or ( n7062 , n7060 , n7061 );
buf ( n7063 , n5583 );
or ( n7064 , n7062 , n7063 );
buf ( n7065 , n5584 );
or ( n7066 , n7064 , n7065 );
buf ( n7067 , n5585 );
or ( n7068 , n7066 , n7067 );
buf ( n7069 , n5586 );
or ( n7070 , n7068 , n7069 );
buf ( n7071 , n5587 );
or ( n7072 , n7070 , n7071 );
buf ( n7073 , n5588 );
or ( n7074 , n7072 , n7073 );
buf ( n7075 , n5589 );
or ( n7076 , n7074 , n7075 );
buf ( n7077 , n5590 );
or ( n7078 , n7076 , n7077 );
buf ( n7079 , n5591 );
or ( n7080 , n7078 , n7079 );
buf ( n7081 , n5592 );
or ( n7082 , n7080 , n7081 );
buf ( n7083 , n5593 );
or ( n7084 , n7082 , n7083 );
buf ( n7085 , n5594 );
or ( n7086 , n7084 , n7085 );
buf ( n7087 , n5595 );
or ( n7088 , n7086 , n7087 );
buf ( n7089 , n5596 );
or ( n7090 , n7088 , n7089 );
buf ( n7091 , n5597 );
or ( n7092 , n7090 , n7091 );
buf ( n7093 , n5598 );
or ( n7094 , n7092 , n7093 );
buf ( n7095 , n5599 );
or ( n7096 , n7094 , n7095 );
buf ( n7097 , n5600 );
or ( n7098 , n7096 , n7097 );
buf ( n7099 , n5601 );
or ( n7100 , n7098 , n7099 );
buf ( n7101 , n5602 );
or ( n7102 , n7100 , n7101 );
buf ( n7103 , n5603 );
or ( n7104 , n7102 , n7103 );
buf ( n7105 , n5604 );
or ( n7106 , n7104 , n7105 );
buf ( n7107 , n5605 );
or ( n7108 , n7106 , n7107 );
buf ( n7109 , n5606 );
or ( n7110 , n7108 , n7109 );
buf ( n7111 , n5607 );
or ( n7112 , n7110 , n7111 );
buf ( n7113 , n5608 );
or ( n7114 , n7112 , n7113 );
buf ( n7115 , n5609 );
or ( n7116 , n7114 , n7115 );
buf ( n7117 , n5610 );
or ( n7118 , n7116 , n7117 );
buf ( n7119 , n5611 );
or ( n7120 , n7118 , n7119 );
buf ( n7121 , n5612 );
or ( n7122 , n7120 , n7121 );
buf ( n7123 , n5613 );
or ( n7124 , n7122 , n7123 );
buf ( n7125 , n5614 );
or ( n7126 , n7124 , n7125 );
buf ( n7127 , n5615 );
or ( n7128 , n7126 , n7127 );
buf ( n7129 , n5616 );
or ( n7130 , n7128 , n7129 );
buf ( n7131 , n5617 );
or ( n7132 , n7130 , n7131 );
buf ( n7133 , n5618 );
or ( n7134 , n7132 , n7133 );
buf ( n7135 , n5619 );
or ( n7136 , n7134 , n7135 );
buf ( n7137 , n5620 );
or ( n7138 , n7136 , n7137 );
buf ( n7139 , n5621 );
or ( n7140 , n7138 , n7139 );
buf ( n7141 , n5622 );
or ( n7142 , n7140 , n7141 );
buf ( n7143 , n5623 );
or ( n7144 , n7142 , n7143 );
buf ( n7145 , n5624 );
or ( n7146 , n7144 , n7145 );
buf ( n7147 , n5625 );
or ( n7148 , n7146 , n7147 );
buf ( n7149 , n5626 );
or ( n7150 , n7148 , n7149 );
buf ( n7151 , n5627 );
or ( n7152 , n7150 , n7151 );
buf ( n7153 , n5628 );
or ( n7154 , n7152 , n7153 );
buf ( n7155 , n5629 );
or ( n7156 , n7154 , n7155 );
buf ( n7157 , n5630 );
or ( n7158 , n7156 , n7157 );
buf ( n7159 , n5631 );
or ( n7160 , n7158 , n7159 );
buf ( n7161 , n5632 );
or ( n7162 , n7160 , n7161 );
buf ( n7163 , n5633 );
or ( n7164 , n7162 , n7163 );
buf ( n7165 , n5634 );
or ( n7166 , n7164 , n7165 );
buf ( n7167 , n5635 );
or ( n7168 , n7166 , n7167 );
buf ( n7169 , n5636 );
or ( n7170 , n7168 , n7169 );
buf ( n7171 , n5637 );
or ( n7172 , n7170 , n7171 );
buf ( n7173 , n5638 );
or ( n7174 , n7172 , n7173 );
buf ( n7175 , n5639 );
or ( n7176 , n7174 , n7175 );
buf ( n7177 , n5640 );
or ( n7178 , n7176 , n7177 );
buf ( n7179 , n5641 );
or ( n7180 , n7178 , n7179 );
buf ( n7181 , n5642 );
or ( n7182 , n7180 , n7181 );
buf ( n7183 , n5643 );
or ( n7184 , n7182 , n7183 );
buf ( n7185 , n5644 );
or ( n7186 , n7184 , n7185 );
buf ( n7187 , n5645 );
or ( n7188 , n7186 , n7187 );
buf ( n7189 , n5646 );
or ( n7190 , n7188 , n7189 );
buf ( n7191 , n5647 );
or ( n7192 , n7190 , n7191 );
buf ( n7193 , n5648 );
or ( n7194 , n7192 , n7193 );
buf ( n7195 , n5649 );
or ( n7196 , n7194 , n7195 );
buf ( n7197 , n5650 );
or ( n7198 , n7196 , n7197 );
buf ( n7199 , n5651 );
or ( n7200 , n7198 , n7199 );
buf ( n7201 , n5652 );
or ( n7202 , n7200 , n7201 );
buf ( n7203 , n5653 );
or ( n7204 , n7202 , n7203 );
buf ( n7205 , n5654 );
or ( n7206 , n7204 , n7205 );
buf ( n7207 , n5655 );
or ( n7208 , n7206 , n7207 );
buf ( n7209 , n5656 );
or ( n7210 , n7208 , n7209 );
buf ( n7211 , n5657 );
or ( n7212 , n7210 , n7211 );
buf ( n7213 , n5658 );
or ( n7214 , n7212 , n7213 );
buf ( n7215 , n5659 );
or ( n7216 , n7214 , n7215 );
buf ( n7217 , n5660 );
or ( n7218 , n7216 , n7217 );
buf ( n7219 , n5661 );
or ( n7220 , n7218 , n7219 );
buf ( n7221 , n5662 );
or ( n7222 , n7220 , n7221 );
buf ( n7223 , n5663 );
or ( n7224 , n7222 , n7223 );
buf ( n7225 , n5664 );
or ( n7226 , n7224 , n7225 );
buf ( n7227 , n5665 );
or ( n7228 , n7226 , n7227 );
buf ( n7229 , n5666 );
or ( n7230 , n7228 , n7229 );
buf ( n7231 , n5667 );
or ( n7232 , n7230 , n7231 );
buf ( n7233 , n5668 );
or ( n7234 , n7232 , n7233 );
buf ( n7235 , n5669 );
or ( n7236 , n7234 , n7235 );
buf ( n7237 , n5670 );
or ( n7238 , n7236 , n7237 );
buf ( n7239 , n5671 );
or ( n7240 , n7238 , n7239 );
buf ( n7241 , n5672 );
or ( n7242 , n7240 , n7241 );
buf ( n7243 , n5673 );
or ( n7244 , n7242 , n7243 );
buf ( n7245 , n5674 );
or ( n7246 , n7244 , n7245 );
buf ( n7247 , n5675 );
or ( n7248 , n7246 , n7247 );
buf ( n7249 , n5676 );
or ( n7250 , n7248 , n7249 );
buf ( n7251 , n5677 );
or ( n7252 , n7250 , n7251 );
buf ( n7253 , n5678 );
or ( n7254 , n7252 , n7253 );
buf ( n7255 , n5679 );
or ( n7256 , n7254 , n7255 );
buf ( n7257 , n5680 );
or ( n7258 , n7256 , n7257 );
buf ( n7259 , n5681 );
or ( n7260 , n7258 , n7259 );
buf ( n7261 , n5682 );
or ( n7262 , n7260 , n7261 );
buf ( n7263 , n5683 );
or ( n7264 , n7262 , n7263 );
buf ( n7265 , n5684 );
or ( n7266 , n7264 , n7265 );
buf ( n7267 , n5685 );
or ( n7268 , n7266 , n7267 );
buf ( n7269 , n5686 );
or ( n7270 , n7268 , n7269 );
buf ( n7271 , n5687 );
or ( n7272 , n7270 , n7271 );
buf ( n7273 , n5688 );
or ( n7274 , n7272 , n7273 );
buf ( n7275 , n5689 );
or ( n7276 , n7274 , n7275 );
buf ( n7277 , n5690 );
or ( n7278 , n7276 , n7277 );
buf ( n7279 , n5691 );
or ( n7280 , n7278 , n7279 );
buf ( n7281 , n5692 );
or ( n7282 , n7280 , n7281 );
buf ( n7283 , n5693 );
or ( n7284 , n7282 , n7283 );
buf ( n7285 , n5694 );
or ( n7286 , n7284 , n7285 );
buf ( n7287 , n5695 );
or ( n7288 , n7286 , n7287 );
buf ( n7289 , n5696 );
or ( n7290 , n7288 , n7289 );
buf ( n7291 , n5697 );
or ( n7292 , n7290 , n7291 );
buf ( n7293 , n5698 );
or ( n7294 , n7292 , n7293 );
buf ( n7295 , n5699 );
or ( n7296 , n7294 , n7295 );
buf ( n7297 , n5700 );
or ( n7298 , n7296 , n7297 );
buf ( n7299 , n5701 );
or ( n7300 , n7298 , n7299 );
buf ( n7301 , n5702 );
or ( n7302 , n7300 , n7301 );
buf ( n7303 , n5703 );
or ( n7304 , n7302 , n7303 );
buf ( n7305 , n5704 );
or ( n7306 , n7304 , n7305 );
buf ( n7307 , n5705 );
or ( n7308 , n7306 , n7307 );
buf ( n7309 , n5706 );
or ( n7310 , n7308 , n7309 );
buf ( n7311 , n5707 );
or ( n7312 , n7310 , n7311 );
buf ( n7313 , n5708 );
or ( n7314 , n7312 , n7313 );
buf ( n7315 , n5709 );
or ( n7316 , n7314 , n7315 );
buf ( n7317 , n5710 );
or ( n7318 , n7316 , n7317 );
buf ( n7319 , n5711 );
or ( n7320 , n7318 , n7319 );
buf ( n7321 , n5712 );
or ( n7322 , n7320 , n7321 );
buf ( n7323 , n5713 );
or ( n7324 , n7322 , n7323 );
buf ( n7325 , n5714 );
or ( n7326 , n7324 , n7325 );
buf ( n7327 , n5715 );
or ( n7328 , n7326 , n7327 );
buf ( n7329 , n5716 );
or ( n7330 , n7328 , n7329 );
buf ( n7331 , n5717 );
or ( n7332 , n7330 , n7331 );
buf ( n7333 , n5718 );
or ( n7334 , n7332 , n7333 );
buf ( n7335 , n5719 );
or ( n7336 , n7334 , n7335 );
buf ( n7337 , n5720 );
or ( n7338 , n7336 , n7337 );
buf ( n7339 , n5721 );
or ( n7340 , n7338 , n7339 );
buf ( n7341 , n5722 );
or ( n7342 , n7340 , n7341 );
buf ( n7343 , n5723 );
or ( n7344 , n7342 , n7343 );
buf ( n7345 , n5724 );
or ( n7346 , n7344 , n7345 );
buf ( n7347 , n5725 );
or ( n7348 , n7346 , n7347 );
buf ( n7349 , n5726 );
or ( n7350 , n7348 , n7349 );
buf ( n7351 , n5727 );
or ( n7352 , n7350 , n7351 );
buf ( n7353 , n5728 );
or ( n7354 , n7352 , n7353 );
buf ( n7355 , n5729 );
or ( n7356 , n7354 , n7355 );
buf ( n7357 , n5730 );
or ( n7358 , n7356 , n7357 );
buf ( n7359 , n5731 );
or ( n7360 , n7358 , n7359 );
buf ( n7361 , n5732 );
or ( n7362 , n7360 , n7361 );
buf ( n7363 , n5733 );
or ( n7364 , n7362 , n7363 );
buf ( n7365 , n5734 );
or ( n7366 , n7364 , n7365 );
buf ( n7367 , n5735 );
or ( n7368 , n7366 , n7367 );
buf ( n7369 , n5736 );
or ( n7370 , n7368 , n7369 );
buf ( n7371 , n5737 );
or ( n7372 , n7370 , n7371 );
buf ( n7373 , n5738 );
or ( n7374 , n7372 , n7373 );
buf ( n7375 , n5739 );
or ( n7376 , n7374 , n7375 );
buf ( n7377 , n5740 );
or ( n7378 , n7376 , n7377 );
buf ( n7379 , n5741 );
or ( n7380 , n7378 , n7379 );
buf ( n7381 , n5742 );
or ( n7382 , n7380 , n7381 );
buf ( n7383 , n5743 );
or ( n7384 , n7382 , n7383 );
buf ( n7385 , n5744 );
or ( n7386 , n7384 , n7385 );
buf ( n7387 , n5745 );
or ( n7388 , n7386 , n7387 );
buf ( n7389 , n5746 );
or ( n7390 , n7388 , n7389 );
buf ( n7391 , n5747 );
or ( n7392 , n7390 , n7391 );
buf ( n7393 , n5748 );
or ( n7394 , n7392 , n7393 );
buf ( n7395 , n5749 );
or ( n7396 , n7394 , n7395 );
buf ( n7397 , n5750 );
or ( n7398 , n7396 , n7397 );
buf ( n7399 , n5751 );
or ( n7400 , n7398 , n7399 );
buf ( n7401 , n5752 );
or ( n7402 , n7400 , n7401 );
buf ( n7403 , n5753 );
or ( n7404 , n7402 , n7403 );
buf ( n7405 , n5754 );
or ( n7406 , n7404 , n7405 );
buf ( n7407 , n5755 );
or ( n7408 , n7406 , n7407 );
buf ( n7409 , n5756 );
or ( n7410 , n7408 , n7409 );
buf ( n7411 , n5757 );
or ( n7412 , n7410 , n7411 );
buf ( n7413 , n5758 );
or ( n7414 , n7412 , n7413 );
buf ( n7415 , n5759 );
or ( n7416 , n7414 , n7415 );
buf ( n7417 , n5760 );
or ( n7418 , n7416 , n7417 );
buf ( n7419 , n5761 );
or ( n7420 , n7418 , n7419 );
buf ( n7421 , n5762 );
or ( n7422 , n7420 , n7421 );
buf ( n7423 , n5763 );
or ( n7424 , n7422 , n7423 );
buf ( n7425 , n5764 );
or ( n7426 , n7424 , n7425 );
buf ( n7427 , n5765 );
or ( n7428 , n7426 , n7427 );
buf ( n7429 , n5766 );
or ( n7430 , n7428 , n7429 );
buf ( n7431 , n5767 );
or ( n7432 , n7430 , n7431 );
buf ( n7433 , n5768 );
or ( n7434 , n7432 , n7433 );
buf ( n7435 , n5769 );
or ( n7436 , n7434 , n7435 );
buf ( n7437 , n5770 );
or ( n7438 , n7436 , n7437 );
buf ( n7439 , n5771 );
or ( n7440 , n7438 , n7439 );
buf ( n7441 , n5772 );
or ( n7442 , n7440 , n7441 );
buf ( n7443 , n5773 );
or ( n7444 , n7442 , n7443 );
buf ( n7445 , n5774 );
or ( n7446 , n7444 , n7445 );
buf ( n7447 , n5775 );
or ( n7448 , n7446 , n7447 );
buf ( n7449 , n5776 );
or ( n7450 , n7448 , n7449 );
buf ( n7451 , n5777 );
or ( n7452 , n7450 , n7451 );
buf ( n7453 , n5778 );
or ( n7454 , n7452 , n7453 );
buf ( n7455 , n5779 );
or ( n7456 , n7454 , n7455 );
buf ( n7457 , n5780 );
or ( n7458 , n7456 , n7457 );
buf ( n7459 , n5781 );
or ( n7460 , n7458 , n7459 );
buf ( n7461 , n5782 );
or ( n7462 , n7460 , n7461 );
buf ( n7463 , n5783 );
or ( n7464 , n7462 , n7463 );
buf ( n7465 , n5784 );
or ( n7466 , n7464 , n7465 );
buf ( n7467 , n5785 );
or ( n7468 , n7466 , n7467 );
buf ( n7469 , n5786 );
or ( n7470 , n7468 , n7469 );
buf ( n7471 , n5787 );
or ( n7472 , n7470 , n7471 );
buf ( n7473 , n5788 );
or ( n7474 , n7472 , n7473 );
buf ( n7475 , n5789 );
or ( n7476 , n7474 , n7475 );
buf ( n7477 , n5790 );
or ( n7478 , n7476 , n7477 );
buf ( n7479 , n5791 );
or ( n7480 , n7478 , n7479 );
buf ( n7481 , n5792 );
or ( n7482 , n7480 , n7481 );
buf ( n7483 , n5793 );
or ( n7484 , n7482 , n7483 );
buf ( n7485 , n5794 );
or ( n7486 , n7484 , n7485 );
buf ( n7487 , n5795 );
or ( n7488 , n7486 , n7487 );
buf ( n7489 , n5796 );
or ( n7490 , n7488 , n7489 );
buf ( n7491 , n5797 );
or ( n7492 , n7490 , n7491 );
buf ( n7493 , n5798 );
or ( n7494 , n7492 , n7493 );
buf ( n7495 , n5799 );
or ( n7496 , n7494 , n7495 );
buf ( n7497 , n5800 );
or ( n7498 , n7496 , n7497 );
buf ( n7499 , n5801 );
or ( n7500 , n7498 , n7499 );
buf ( n7501 , n5802 );
or ( n7502 , n7500 , n7501 );
buf ( n7503 , n5803 );
or ( n7504 , n7502 , n7503 );
buf ( n7505 , n5804 );
or ( n7506 , n7504 , n7505 );
buf ( n7507 , n5805 );
or ( n7508 , n7506 , n7507 );
buf ( n7509 , n5806 );
or ( n7510 , n7508 , n7509 );
buf ( n7511 , n5807 );
or ( n7512 , n7510 , n7511 );
buf ( n7513 , n5808 );
or ( n7514 , n7512 , n7513 );
buf ( n7515 , n5809 );
or ( n7516 , n7514 , n7515 );
buf ( n7517 , n5810 );
or ( n7518 , n7516 , n7517 );
buf ( n7519 , n5811 );
or ( n7520 , n7518 , n7519 );
buf ( n7521 , n5812 );
or ( n7522 , n7520 , n7521 );
buf ( n7523 , n5813 );
or ( n7524 , n7522 , n7523 );
buf ( n7525 , n5814 );
or ( n7526 , n7524 , n7525 );
buf ( n7527 , n5815 );
or ( n7528 , n7526 , n7527 );
buf ( n7529 , n5816 );
or ( n7530 , n7528 , n7529 );
buf ( n7531 , n5817 );
or ( n7532 , n7530 , n7531 );
buf ( n7533 , n5818 );
or ( n7534 , n7532 , n7533 );
buf ( n7535 , n5819 );
or ( n7536 , n7534 , n7535 );
buf ( n7537 , n5820 );
or ( n7538 , n7536 , n7537 );
buf ( n7539 , n5821 );
or ( n7540 , n7538 , n7539 );
buf ( n7541 , n5822 );
or ( n7542 , n7540 , n7541 );
buf ( n7543 , n5823 );
or ( n7544 , n7542 , n7543 );
buf ( n7545 , n5824 );
or ( n7546 , n7544 , n7545 );
buf ( n7547 , n5825 );
or ( n7548 , n7546 , n7547 );
buf ( n7549 , n5826 );
or ( n7550 , n7548 , n7549 );
buf ( n7551 , n5827 );
or ( n7552 , n7550 , n7551 );
buf ( n7553 , n5828 );
or ( n7554 , n7552 , n7553 );
buf ( n7555 , n5829 );
or ( n7556 , n7554 , n7555 );
buf ( n7557 , n5830 );
or ( n7558 , n7556 , n7557 );
buf ( n7559 , n5831 );
or ( n7560 , n7558 , n7559 );
buf ( n7561 , n5832 );
or ( n7562 , n7560 , n7561 );
buf ( n7563 , n5833 );
or ( n7564 , n7562 , n7563 );
buf ( n7565 , n5834 );
or ( n7566 , n7564 , n7565 );
buf ( n7567 , n5835 );
or ( n7568 , n7566 , n7567 );
buf ( n7569 , n5836 );
or ( n7570 , n7568 , n7569 );
buf ( n7571 , n5837 );
or ( n7572 , n7570 , n7571 );
buf ( n7573 , n5838 );
or ( n7574 , n7572 , n7573 );
buf ( n7575 , n5839 );
or ( n7576 , n7574 , n7575 );
buf ( n7577 , n5840 );
or ( n7578 , n7576 , n7577 );
buf ( n7579 , n5841 );
or ( n7580 , n7578 , n7579 );
buf ( n7581 , n5842 );
or ( n7582 , n7580 , n7581 );
buf ( n7583 , n5843 );
or ( n7584 , n7582 , n7583 );
buf ( n7585 , n5844 );
or ( n7586 , n7584 , n7585 );
buf ( n7587 , n5845 );
or ( n7588 , n7586 , n7587 );
buf ( n7589 , n5846 );
or ( n7590 , n7588 , n7589 );
buf ( n7591 , n5847 );
or ( n7592 , n7590 , n7591 );
buf ( n7593 , n5848 );
or ( n7594 , n7592 , n7593 );
buf ( n7595 , n5849 );
or ( n7596 , n7594 , n7595 );
buf ( n7597 , n5850 );
or ( n7598 , n7596 , n7597 );
buf ( n7599 , n5851 );
or ( n7600 , n7598 , n7599 );
buf ( n7601 , n5852 );
or ( n7602 , n7600 , n7601 );
buf ( n7603 , n5853 );
or ( n7604 , n7602 , n7603 );
buf ( n7605 , n5854 );
or ( n7606 , n7604 , n7605 );
buf ( n7607 , n5855 );
or ( n7608 , n7606 , n7607 );
buf ( n7609 , n5856 );
or ( n7610 , n7608 , n7609 );
buf ( n7611 , n5857 );
or ( n7612 , n7610 , n7611 );
buf ( n7613 , n5858 );
or ( n7614 , n7612 , n7613 );
buf ( n7615 , n5859 );
or ( n7616 , n7614 , n7615 );
buf ( n7617 , n5860 );
or ( n7618 , n7616 , n7617 );
buf ( n7619 , n5861 );
or ( n7620 , n7618 , n7619 );
buf ( n7621 , n5862 );
or ( n7622 , n7620 , n7621 );
buf ( n7623 , n5863 );
or ( n7624 , n7622 , n7623 );
buf ( n7625 , n5864 );
or ( n7626 , n7624 , n7625 );
buf ( n7627 , n5865 );
or ( n7628 , n7626 , n7627 );
buf ( n7629 , n5866 );
or ( n7630 , n7628 , n7629 );
buf ( n7631 , n5867 );
or ( n7632 , n7630 , n7631 );
buf ( n7633 , n5868 );
or ( n7634 , n7632 , n7633 );
buf ( n7635 , n5869 );
or ( n7636 , n7634 , n7635 );
buf ( n7637 , n5870 );
or ( n7638 , n7636 , n7637 );
buf ( n7639 , n5871 );
or ( n7640 , n7638 , n7639 );
buf ( n7641 , n5872 );
or ( n7642 , n7640 , n7641 );
buf ( n7643 , n5873 );
or ( n7644 , n7642 , n7643 );
buf ( n7645 , n5874 );
or ( n7646 , n7644 , n7645 );
buf ( n7647 , n5875 );
or ( n7648 , n7646 , n7647 );
buf ( n7649 , n5876 );
or ( n7650 , n7648 , n7649 );
buf ( n7651 , n5877 );
or ( n7652 , n7650 , n7651 );
buf ( n7653 , n5878 );
or ( n7654 , n7652 , n7653 );
buf ( n7655 , n5879 );
or ( n7656 , n7654 , n7655 );
buf ( n7657 , n5880 );
or ( n7658 , n7656 , n7657 );
buf ( n7659 , n5881 );
or ( n7660 , n7658 , n7659 );
buf ( n7661 , n5882 );
or ( n7662 , n7660 , n7661 );
buf ( n7663 , n5883 );
or ( n7664 , n7662 , n7663 );
buf ( n7665 , n5884 );
or ( n7666 , n7664 , n7665 );
buf ( n7667 , n5885 );
or ( n7668 , n7666 , n7667 );
buf ( n7669 , n5886 );
or ( n7670 , n7668 , n7669 );
buf ( n7671 , n5887 );
or ( n7672 , n7670 , n7671 );
buf ( n7673 , n5888 );
or ( n7674 , n7672 , n7673 );
buf ( n7675 , n5889 );
or ( n7676 , n7674 , n7675 );
buf ( n7677 , n5890 );
or ( n7678 , n7676 , n7677 );
buf ( n7679 , n5891 );
or ( n7680 , n7678 , n7679 );
buf ( n7681 , n5892 );
or ( n7682 , n7680 , n7681 );
buf ( n7683 , n5893 );
or ( n7684 , n7682 , n7683 );
buf ( n7685 , n5894 );
or ( n7686 , n7684 , n7685 );
buf ( n7687 , n5895 );
or ( n7688 , n7686 , n7687 );
buf ( n7689 , n5896 );
or ( n7690 , n7688 , n7689 );
buf ( n7691 , n5897 );
or ( n7692 , n7690 , n7691 );
buf ( n7693 , n5898 );
or ( n7694 , n7692 , n7693 );
buf ( n7695 , n5899 );
or ( n7696 , n7694 , n7695 );
buf ( n7697 , n5900 );
or ( n7698 , n7696 , n7697 );
buf ( n7699 , n5901 );
or ( n7700 , n7698 , n7699 );
buf ( n7701 , n5902 );
or ( n7702 , n7700 , n7701 );
buf ( n7703 , n5903 );
or ( n7704 , n7702 , n7703 );
buf ( n7705 , n5904 );
or ( n7706 , n7704 , n7705 );
buf ( n7707 , n5905 );
or ( n7708 , n7706 , n7707 );
buf ( n7709 , n5906 );
or ( n7710 , n7708 , n7709 );
buf ( n7711 , n5907 );
or ( n7712 , n7710 , n7711 );
buf ( n7713 , n5908 );
or ( n7714 , n7712 , n7713 );
buf ( n7715 , n5909 );
or ( n7716 , n7714 , n7715 );
buf ( n7717 , n5910 );
or ( n7718 , n7716 , n7717 );
buf ( n7719 , n5911 );
or ( n7720 , n7718 , n7719 );
buf ( n7721 , n5912 );
or ( n7722 , n7720 , n7721 );
buf ( n7723 , n5913 );
or ( n7724 , n7722 , n7723 );
buf ( n7725 , n5914 );
or ( n7726 , n7724 , n7725 );
buf ( n7727 , n5915 );
or ( n7728 , n7726 , n7727 );
buf ( n7729 , n5916 );
or ( n7730 , n7728 , n7729 );
buf ( n7731 , n5917 );
or ( n7732 , n7730 , n7731 );
buf ( n7733 , n5918 );
or ( n7734 , n7732 , n7733 );
buf ( n7735 , n5919 );
or ( n7736 , n7734 , n7735 );
buf ( n7737 , n5920 );
or ( n7738 , n7736 , n7737 );
buf ( n7739 , n5921 );
or ( n7740 , n7738 , n7739 );
buf ( n7741 , n5922 );
or ( n7742 , n7740 , n7741 );
buf ( n7743 , n5923 );
or ( n7744 , n7742 , n7743 );
buf ( n7745 , n5924 );
or ( n7746 , n7744 , n7745 );
buf ( n7747 , n5925 );
or ( n7748 , n7746 , n7747 );
buf ( n7749 , n5926 );
or ( n7750 , n7748 , n7749 );
buf ( n7751 , n5927 );
or ( n7752 , n7750 , n7751 );
buf ( n7753 , n5928 );
or ( n7754 , n7752 , n7753 );
buf ( n7755 , n5929 );
or ( n7756 , n7754 , n7755 );
buf ( n7757 , n5930 );
or ( n7758 , n7756 , n7757 );
buf ( n7759 , n5931 );
or ( n7760 , n7758 , n7759 );
buf ( n7761 , n5932 );
or ( n7762 , n7760 , n7761 );
buf ( n7763 , n5933 );
or ( n7764 , n7762 , n7763 );
buf ( n7765 , n5934 );
or ( n7766 , n7764 , n7765 );
buf ( n7767 , n5935 );
or ( n7768 , n7766 , n7767 );
buf ( n7769 , n5936 );
or ( n7770 , n7768 , n7769 );
buf ( n7771 , n5937 );
or ( n7772 , n7770 , n7771 );
buf ( n7773 , n5938 );
or ( n7774 , n7772 , n7773 );
buf ( n7775 , n5939 );
or ( n7776 , n7774 , n7775 );
buf ( n7777 , n5940 );
or ( n7778 , n7776 , n7777 );
buf ( n7779 , n5941 );
or ( n7780 , n7778 , n7779 );
buf ( n7781 , n5942 );
or ( n7782 , n7780 , n7781 );
buf ( n7783 , n5943 );
or ( n7784 , n7782 , n7783 );
buf ( n7785 , n5944 );
or ( n7786 , n7784 , n7785 );
buf ( n7787 , n5945 );
or ( n7788 , n7786 , n7787 );
buf ( n7789 , n5946 );
or ( n7790 , n7788 , n7789 );
buf ( n7791 , n5947 );
or ( n7792 , n7790 , n7791 );
buf ( n7793 , n5948 );
or ( n7794 , n7792 , n7793 );
buf ( n7795 , n5949 );
or ( n7796 , n7794 , n7795 );
buf ( n7797 , n5950 );
or ( n7798 , n7796 , n7797 );
buf ( n7799 , n5951 );
or ( n7800 , n7798 , n7799 );
buf ( n7801 , n5952 );
or ( n7802 , n7800 , n7801 );
buf ( n7803 , n5953 );
or ( n7804 , n7802 , n7803 );
buf ( n7805 , n5954 );
or ( n7806 , n7804 , n7805 );
buf ( n7807 , n5955 );
or ( n7808 , n7806 , n7807 );
buf ( n7809 , n5956 );
or ( n7810 , n7808 , n7809 );
buf ( n7811 , n5957 );
or ( n7812 , n7810 , n7811 );
buf ( n7813 , n5958 );
or ( n7814 , n7812 , n7813 );
buf ( n7815 , n5959 );
or ( n7816 , n7814 , n7815 );
buf ( n7817 , n5960 );
or ( n7818 , n7816 , n7817 );
buf ( n7819 , n5961 );
or ( n7820 , n7818 , n7819 );
buf ( n7821 , n5962 );
or ( n7822 , n7820 , n7821 );
buf ( n7823 , n5963 );
or ( n7824 , n7822 , n7823 );
buf ( n7825 , n5964 );
or ( n7826 , n7824 , n7825 );
buf ( n7827 , n5965 );
or ( n7828 , n7826 , n7827 );
buf ( n7829 , n5966 );
or ( n7830 , n7828 , n7829 );
buf ( n7831 , n5967 );
or ( n7832 , n7830 , n7831 );
buf ( n7833 , n5968 );
or ( n7834 , n7832 , n7833 );
buf ( n7835 , n5969 );
or ( n7836 , n7834 , n7835 );
buf ( n7837 , n5970 );
or ( n7838 , n7836 , n7837 );
buf ( n7839 , n5971 );
or ( n7840 , n7838 , n7839 );
buf ( n7841 , n5972 );
or ( n7842 , n7840 , n7841 );
buf ( n7843 , n5973 );
or ( n7844 , n7842 , n7843 );
buf ( n7845 , n5974 );
or ( n7846 , n7844 , n7845 );
buf ( n7847 , n5975 );
or ( n7848 , n7846 , n7847 );
buf ( n7849 , n5976 );
or ( n7850 , n7848 , n7849 );
buf ( n7851 , n5977 );
or ( n7852 , n7850 , n7851 );
buf ( n7853 , n5978 );
or ( n7854 , n7852 , n7853 );
buf ( n7855 , n5979 );
or ( n7856 , n7854 , n7855 );
buf ( n7857 , n5980 );
or ( n7858 , n7856 , n7857 );
buf ( n7859 , n5981 );
or ( n7860 , n7858 , n7859 );
buf ( n7861 , n5982 );
or ( n7862 , n7860 , n7861 );
buf ( n7863 , n5983 );
or ( n7864 , n7862 , n7863 );
buf ( n7865 , n5984 );
or ( n7866 , n7864 , n7865 );
buf ( n7867 , n5985 );
or ( n7868 , n7866 , n7867 );
buf ( n7869 , n5986 );
or ( n7870 , n7868 , n7869 );
buf ( n7871 , n5987 );
or ( n7872 , n7870 , n7871 );
buf ( n7873 , n5988 );
or ( n7874 , n7872 , n7873 );
buf ( n7875 , n5989 );
or ( n7876 , n7874 , n7875 );
buf ( n7877 , n5990 );
or ( n7878 , n7876 , n7877 );
buf ( n7879 , n5991 );
or ( n7880 , n7878 , n7879 );
buf ( n7881 , n5992 );
or ( n7882 , n7880 , n7881 );
buf ( n7883 , n5993 );
or ( n7884 , n7882 , n7883 );
buf ( n7885 , n5994 );
or ( n7886 , n7884 , n7885 );
buf ( n7887 , n5995 );
or ( n7888 , n7886 , n7887 );
buf ( n7889 , n5996 );
or ( n7890 , n7888 , n7889 );
buf ( n7891 , n5997 );
or ( n7892 , n7890 , n7891 );
buf ( n7893 , n5998 );
or ( n7894 , n7892 , n7893 );
buf ( n7895 , n5999 );
or ( n7896 , n7894 , n7895 );
buf ( n7897 , n6000 );
or ( n7898 , n7896 , n7897 );
buf ( n7899 , n6001 );
or ( n7900 , n7898 , n7899 );
buf ( n7901 , n6002 );
or ( n7902 , n7900 , n7901 );
buf ( n7903 , n6003 );
or ( n7904 , n7902 , n7903 );
buf ( n7905 , n6004 );
or ( n7906 , n7904 , n7905 );
buf ( n7907 , n6005 );
or ( n7908 , n7906 , n7907 );
buf ( n7909 , n6006 );
or ( n7910 , n7908 , n7909 );
buf ( n7911 , n6007 );
or ( n7912 , n7910 , n7911 );
buf ( n7913 , n6008 );
or ( n7914 , n7912 , n7913 );
buf ( n7915 , n6009 );
or ( n7916 , n7914 , n7915 );
buf ( n7917 , n6010 );
or ( n7918 , n7916 , n7917 );
buf ( n7919 , n6011 );
or ( n7920 , n7918 , n7919 );
buf ( n7921 , n6012 );
or ( n7922 , n7920 , n7921 );
buf ( n7923 , n6013 );
or ( n7924 , n7922 , n7923 );
buf ( n7925 , n6014 );
or ( n7926 , n7924 , n7925 );
buf ( n7927 , n6015 );
or ( n7928 , n7926 , n7927 );
buf ( n7929 , n6016 );
or ( n7930 , n7928 , n7929 );
buf ( n7931 , n6017 );
or ( n7932 , n7930 , n7931 );
buf ( n7933 , n6018 );
or ( n7934 , n7932 , n7933 );
buf ( n7935 , n6019 );
or ( n7936 , n7934 , n7935 );
buf ( n7937 , n6020 );
or ( n7938 , n7936 , n7937 );
buf ( n7939 , n6021 );
or ( n7940 , n7938 , n7939 );
buf ( n7941 , n6022 );
or ( n7942 , n7940 , n7941 );
buf ( n7943 , n6023 );
or ( n7944 , n7942 , n7943 );
buf ( n7945 , n6024 );
or ( n7946 , n7944 , n7945 );
buf ( n7947 , n6025 );
or ( n7948 , n7946 , n7947 );
buf ( n7949 , n6026 );
or ( n7950 , n7948 , n7949 );
buf ( n7951 , n6027 );
or ( n7952 , n7950 , n7951 );
buf ( n7953 , n6028 );
or ( n7954 , n7952 , n7953 );
buf ( n7955 , n6029 );
or ( n7956 , n7954 , n7955 );
buf ( n7957 , n6030 );
or ( n7958 , n7956 , n7957 );
buf ( n7959 , n6031 );
or ( n7960 , n7958 , n7959 );
buf ( n7961 , n6032 );
or ( n7962 , n7960 , n7961 );
buf ( n7963 , n6033 );
or ( n7964 , n7962 , n7963 );
buf ( n7965 , n6034 );
or ( n7966 , n7964 , n7965 );
buf ( n7967 , n6035 );
or ( n7968 , n7966 , n7967 );
buf ( n7969 , n6036 );
or ( n7970 , n7968 , n7969 );
buf ( n7971 , n6037 );
or ( n7972 , n7970 , n7971 );
buf ( n7973 , n6038 );
or ( n7974 , n7972 , n7973 );
buf ( n7975 , n6039 );
or ( n7976 , n7974 , n7975 );
buf ( n7977 , n6040 );
or ( n7978 , n7976 , n7977 );
buf ( n7979 , n6041 );
or ( n7980 , n7978 , n7979 );
buf ( n7981 , n6042 );
or ( n7982 , n7980 , n7981 );
buf ( n7983 , n6043 );
or ( n7984 , n7982 , n7983 );
buf ( n7985 , n6044 );
or ( n7986 , n7984 , n7985 );
buf ( n7987 , n6045 );
or ( n7988 , n7986 , n7987 );
buf ( n7989 , n6046 );
or ( n7990 , n7988 , n7989 );
buf ( n7991 , n6047 );
or ( n7992 , n7990 , n7991 );
buf ( n7993 , n6048 );
or ( n7994 , n7992 , n7993 );
buf ( n7995 , n6049 );
or ( n7996 , n7994 , n7995 );
buf ( n7997 , n6050 );
or ( n7998 , n7996 , n7997 );
buf ( n7999 , n6051 );
or ( n8000 , n7998 , n7999 );
buf ( n8001 , n6052 );
or ( n8002 , n8000 , n8001 );
buf ( n8003 , n6053 );
or ( n8004 , n8002 , n8003 );
buf ( n8005 , n6054 );
or ( n8006 , n8004 , n8005 );
buf ( n8007 , n6055 );
or ( n8008 , n8006 , n8007 );
buf ( n8009 , n6056 );
or ( n8010 , n8008 , n8009 );
buf ( n8011 , n6057 );
or ( n8012 , n8010 , n8011 );
buf ( n8013 , n6058 );
or ( n8014 , n8012 , n8013 );
buf ( n8015 , n6059 );
or ( n8016 , n8014 , n8015 );
buf ( n8017 , n6060 );
or ( n8018 , n8016 , n8017 );
buf ( n8019 , n6061 );
or ( n8020 , n8018 , n8019 );
buf ( n8021 , n6062 );
or ( n8022 , n8020 , n8021 );
buf ( n8023 , n6063 );
or ( n8024 , n8022 , n8023 );
buf ( n8025 , n6064 );
or ( n8026 , n8024 , n8025 );
buf ( n8027 , n6065 );
or ( n8028 , n8026 , n8027 );
buf ( n8029 , n6066 );
or ( n8030 , n8028 , n8029 );
buf ( n8031 , n6067 );
or ( n8032 , n8030 , n8031 );
buf ( n8033 , n6068 );
or ( n8034 , n8032 , n8033 );
buf ( n8035 , n6069 );
or ( n8036 , n8034 , n8035 );
buf ( n8037 , n6070 );
or ( n8038 , n8036 , n8037 );
buf ( n8039 , n6071 );
or ( n8040 , n8038 , n8039 );
buf ( n8041 , n6072 );
or ( n8042 , n8040 , n8041 );
buf ( n8043 , n6073 );
or ( n8044 , n8042 , n8043 );
buf ( n8045 , n6074 );
or ( n8046 , n8044 , n8045 );
buf ( n8047 , n6075 );
or ( n8048 , n8046 , n8047 );
buf ( n8049 , n6076 );
or ( n8050 , n8048 , n8049 );
buf ( n8051 , n6077 );
or ( n8052 , n8050 , n8051 );
buf ( n8053 , n6078 );
or ( n8054 , n8052 , n8053 );
buf ( n8055 , n6079 );
or ( n8056 , n8054 , n8055 );
buf ( n8057 , n6080 );
or ( n8058 , n8056 , n8057 );
buf ( n8059 , n6081 );
or ( n8060 , n8058 , n8059 );
buf ( n8061 , n6082 );
or ( n8062 , n8060 , n8061 );
buf ( n8063 , n6083 );
or ( n8064 , n8062 , n8063 );
buf ( n8065 , n6084 );
or ( n8066 , n8064 , n8065 );
buf ( n8067 , n6085 );
or ( n8068 , n8066 , n8067 );
buf ( n8069 , n6086 );
or ( n8070 , n8068 , n8069 );
buf ( n8071 , n6087 );
or ( n8072 , n8070 , n8071 );
buf ( n8073 , n6088 );
or ( n8074 , n8072 , n8073 );
buf ( n8075 , n6089 );
or ( n8076 , n8074 , n8075 );
buf ( n8077 , n6090 );
or ( n8078 , n8076 , n8077 );
buf ( n8079 , n6091 );
or ( n8080 , n8078 , n8079 );
buf ( n8081 , n6092 );
or ( n8082 , n8080 , n8081 );
buf ( n8083 , n6093 );
or ( n8084 , n8082 , n8083 );
buf ( n8085 , n6094 );
or ( n8086 , n8084 , n8085 );
buf ( n8087 , n6095 );
or ( n8088 , n8086 , n8087 );
buf ( n8089 , n6096 );
or ( n8090 , n8088 , n8089 );
buf ( n8091 , n6097 );
or ( n8092 , n8090 , n8091 );
buf ( n8093 , n6098 );
or ( n8094 , n8092 , n8093 );
buf ( n8095 , n6099 );
or ( n8096 , n8094 , n8095 );
buf ( n8097 , n6100 );
or ( n8098 , n8096 , n8097 );
buf ( n8099 , n6101 );
or ( n8100 , n8098 , n8099 );
buf ( n8101 , n6102 );
or ( n8102 , n8100 , n8101 );
buf ( n8103 , n6103 );
or ( n8104 , n8102 , n8103 );
buf ( n8105 , n6104 );
or ( n8106 , n8104 , n8105 );
buf ( n8107 , n6105 );
or ( n8108 , n8106 , n8107 );
buf ( n8109 , n6106 );
or ( n8110 , n8108 , n8109 );
buf ( n8111 , n6107 );
or ( n8112 , n8110 , n8111 );
buf ( n8113 , n6108 );
or ( n8114 , n8112 , n8113 );
buf ( n8115 , n6109 );
or ( n8116 , n8114 , n8115 );
buf ( n8117 , n6110 );
or ( n8118 , n8116 , n8117 );
buf ( n8119 , n6111 );
or ( n8120 , n8118 , n8119 );
buf ( n8121 , n6112 );
or ( n8122 , n8120 , n8121 );
buf ( n8123 , n6113 );
or ( n8124 , n8122 , n8123 );
buf ( n8125 , n6114 );
or ( n8126 , n8124 , n8125 );
buf ( n8127 , n6115 );
or ( n8128 , n8126 , n8127 );
buf ( n8129 , n5092 );
buf ( n8130 , n6116 );
xor ( n8131 , n8129 , n8130 );
or ( n8132 , n8128 , n8131 );
buf ( n8133 , n6117 );
or ( n8134 , n8132 , n8133 );
buf ( n8135 , n5094 );
buf ( n8136 , n6118 );
xor ( n8137 , n8135 , n8136 );
or ( n8138 , n8134 , n8137 );
buf ( n8139 , n6119 );
or ( n8140 , n8138 , n8139 );
buf ( n8141 , n6120 );
or ( n8142 , n8140 , n8141 );
buf ( n8143 , n5097 );
buf ( n8144 , n6121 );
xor ( n8145 , n8143 , n8144 );
or ( n8146 , n8142 , n8145 );
buf ( n8147 , n6122 );
or ( n8148 , n8146 , n8147 );
buf ( n8149 , n5099 );
buf ( n8150 , n6123 );
xor ( n8151 , n8149 , n8150 );
or ( n8152 , n8148 , n8151 );
buf ( n8153 , n5100 );
buf ( n8154 , n6124 );
xor ( n8155 , n8153 , n8154 );
or ( n8156 , n8152 , n8155 );
buf ( n8157 , n6125 );
or ( n8158 , n8156 , n8157 );
buf ( n8159 , n6126 );
or ( n8160 , n8158 , n8159 );
buf ( n8161 , n5103 );
buf ( n8162 , n6127 );
xor ( n8163 , n8161 , n8162 );
or ( n8164 , n8160 , n8163 );
buf ( n8165 , n6128 );
or ( n8166 , n8164 , n8165 );
buf ( n8167 , n6129 );
or ( n8168 , n8166 , n8167 );
buf ( n8169 , n6130 );
or ( n8170 , n8168 , n8169 );
buf ( n8171 , n5107 );
buf ( n8172 , n6131 );
xor ( n8173 , n8171 , n8172 );
or ( n8174 , n8170 , n8173 );
buf ( n8175 , n6132 );
or ( n8176 , n8174 , n8175 );
buf ( n8177 , n6133 );
or ( n8178 , n8176 , n8177 );
buf ( n8179 , n6134 );
or ( n8180 , n8178 , n8179 );
buf ( n8181 , n5111 );
buf ( n8182 , n6135 );
xor ( n8183 , n8181 , n8182 );
or ( n8184 , n8180 , n8183 );
buf ( n8185 , n5112 );
buf ( n8186 , n6136 );
xor ( n8187 , n8185 , n8186 );
or ( n8188 , n8184 , n8187 );
buf ( n8189 , n6137 );
or ( n8190 , n8188 , n8189 );
buf ( n8191 , n5114 );
buf ( n8192 , n6138 );
xor ( n8193 , n8191 , n8192 );
or ( n8194 , n8190 , n8193 );
buf ( n8195 , n6139 );
or ( n8196 , n8194 , n8195 );
buf ( n8197 , n6140 );
or ( n8198 , n8196 , n8197 );
buf ( n8199 , n6141 );
or ( n8200 , n8198 , n8199 );
buf ( n8201 , n5118 );
buf ( n8202 , n6142 );
xor ( n8203 , n8201 , n8202 );
or ( n8204 , n8200 , n8203 );
buf ( n8205 , n5119 );
buf ( n8206 , n6143 );
xor ( n8207 , n8205 , n8206 );
or ( n8208 , n8204 , n8207 );
buf ( n8209 , n6144 );
or ( n8210 , n8208 , n8209 );
buf ( n8211 , n5121 );
buf ( n8212 , n6145 );
xor ( n8213 , n8211 , n8212 );
or ( n8214 , n8210 , n8213 );
buf ( n8215 , n5122 );
buf ( n8216 , n6146 );
xor ( n8217 , n8215 , n8216 );
or ( n8218 , n8214 , n8217 );
buf ( n8219 , n6147 );
or ( n8220 , n8218 , n8219 );
buf ( n8221 , n5124 );
buf ( n8222 , n6148 );
xor ( n8223 , n8221 , n8222 );
or ( n8224 , n8220 , n8223 );
buf ( n8225 , n5125 );
buf ( n8226 , n6149 );
xor ( n8227 , n8225 , n8226 );
or ( n8228 , n8224 , n8227 );
buf ( n8229 , n8228 );
buf ( n8230 , n8229 );
buf ( n8231 , n4102 );
buf ( n8232 , n5126 );
xor ( n8233 , n8231 , n8232 );
buf ( n8234 , n4103 );
buf ( n8235 , n5127 );
xor ( n8236 , n8234 , n8235 );
or ( n8237 , n8233 , n8236 );
buf ( n8238 , n4104 );
buf ( n8239 , n5128 );
xor ( n8240 , n8238 , n8239 );
or ( n8241 , n8237 , n8240 );
buf ( n8242 , n4105 );
buf ( n8243 , n5129 );
xor ( n8244 , n8242 , n8243 );
or ( n8245 , n8241 , n8244 );
buf ( n8246 , n4106 );
buf ( n8247 , n5130 );
xor ( n8248 , n8246 , n8247 );
or ( n8249 , n8245 , n8248 );
buf ( n8250 , n4107 );
buf ( n8251 , n5131 );
xor ( n8252 , n8250 , n8251 );
or ( n8253 , n8249 , n8252 );
buf ( n8254 , n4108 );
buf ( n8255 , n5132 );
xor ( n8256 , n8254 , n8255 );
or ( n8257 , n8253 , n8256 );
buf ( n8258 , n4109 );
buf ( n8259 , n5133 );
xor ( n8260 , n8258 , n8259 );
or ( n8261 , n8257 , n8260 );
buf ( n8262 , n4110 );
buf ( n8263 , n5134 );
xor ( n8264 , n8262 , n8263 );
or ( n8265 , n8261 , n8264 );
buf ( n8266 , n4111 );
buf ( n8267 , n5135 );
xor ( n8268 , n8266 , n8267 );
or ( n8269 , n8265 , n8268 );
buf ( n8270 , n4112 );
buf ( n8271 , n5136 );
xor ( n8272 , n8270 , n8271 );
or ( n8273 , n8269 , n8272 );
buf ( n8274 , n4113 );
buf ( n8275 , n5137 );
xor ( n8276 , n8274 , n8275 );
or ( n8277 , n8273 , n8276 );
buf ( n8278 , n4114 );
buf ( n8279 , n5138 );
xor ( n8280 , n8278 , n8279 );
or ( n8281 , n8277 , n8280 );
buf ( n8282 , n4115 );
buf ( n8283 , n5139 );
xor ( n8284 , n8282 , n8283 );
or ( n8285 , n8281 , n8284 );
buf ( n8286 , n4116 );
buf ( n8287 , n5140 );
xor ( n8288 , n8286 , n8287 );
or ( n8289 , n8285 , n8288 );
buf ( n8290 , n4117 );
buf ( n8291 , n5141 );
xor ( n8292 , n8290 , n8291 );
or ( n8293 , n8289 , n8292 );
buf ( n8294 , n4118 );
buf ( n8295 , n5142 );
xor ( n8296 , n8294 , n8295 );
or ( n8297 , n8293 , n8296 );
buf ( n8298 , n4119 );
buf ( n8299 , n5143 );
xor ( n8300 , n8298 , n8299 );
or ( n8301 , n8297 , n8300 );
buf ( n8302 , n4120 );
buf ( n8303 , n5144 );
xor ( n8304 , n8302 , n8303 );
or ( n8305 , n8301 , n8304 );
buf ( n8306 , n4121 );
buf ( n8307 , n5145 );
xor ( n8308 , n8306 , n8307 );
or ( n8309 , n8305 , n8308 );
buf ( n8310 , n4122 );
buf ( n8311 , n5146 );
xor ( n8312 , n8310 , n8311 );
or ( n8313 , n8309 , n8312 );
buf ( n8314 , n4123 );
buf ( n8315 , n5147 );
xor ( n8316 , n8314 , n8315 );
or ( n8317 , n8313 , n8316 );
buf ( n8318 , n4124 );
buf ( n8319 , n5148 );
xor ( n8320 , n8318 , n8319 );
or ( n8321 , n8317 , n8320 );
buf ( n8322 , n4125 );
buf ( n8323 , n5149 );
xor ( n8324 , n8322 , n8323 );
or ( n8325 , n8321 , n8324 );
buf ( n8326 , n4126 );
buf ( n8327 , n5150 );
xor ( n8328 , n8326 , n8327 );
or ( n8329 , n8325 , n8328 );
buf ( n8330 , n4127 );
buf ( n8331 , n5151 );
xor ( n8332 , n8330 , n8331 );
or ( n8333 , n8329 , n8332 );
buf ( n8334 , n4128 );
buf ( n8335 , n5152 );
xor ( n8336 , n8334 , n8335 );
or ( n8337 , n8333 , n8336 );
buf ( n8338 , n4129 );
buf ( n8339 , n5153 );
xor ( n8340 , n8338 , n8339 );
or ( n8341 , n8337 , n8340 );
buf ( n8342 , n4130 );
buf ( n8343 , n5154 );
xor ( n8344 , n8342 , n8343 );
or ( n8345 , n8341 , n8344 );
buf ( n8346 , n4131 );
buf ( n8347 , n5155 );
xor ( n8348 , n8346 , n8347 );
or ( n8349 , n8345 , n8348 );
buf ( n8350 , n4132 );
buf ( n8351 , n5156 );
xor ( n8352 , n8350 , n8351 );
or ( n8353 , n8349 , n8352 );
buf ( n8354 , n4133 );
buf ( n8355 , n5157 );
xor ( n8356 , n8354 , n8355 );
or ( n8357 , n8353 , n8356 );
buf ( n8358 , n4134 );
buf ( n8359 , n5158 );
xor ( n8360 , n8358 , n8359 );
or ( n8361 , n8357 , n8360 );
buf ( n8362 , n4135 );
buf ( n8363 , n5159 );
xor ( n8364 , n8362 , n8363 );
or ( n8365 , n8361 , n8364 );
buf ( n8366 , n4136 );
buf ( n8367 , n5160 );
xor ( n8368 , n8366 , n8367 );
or ( n8369 , n8365 , n8368 );
buf ( n8370 , n4137 );
buf ( n8371 , n5161 );
xor ( n8372 , n8370 , n8371 );
or ( n8373 , n8369 , n8372 );
buf ( n8374 , n4138 );
buf ( n8375 , n5162 );
xor ( n8376 , n8374 , n8375 );
or ( n8377 , n8373 , n8376 );
buf ( n8378 , n4139 );
buf ( n8379 , n5163 );
xor ( n8380 , n8378 , n8379 );
or ( n8381 , n8377 , n8380 );
buf ( n8382 , n4140 );
buf ( n8383 , n5164 );
xor ( n8384 , n8382 , n8383 );
or ( n8385 , n8381 , n8384 );
buf ( n8386 , n4141 );
buf ( n8387 , n5165 );
xor ( n8388 , n8386 , n8387 );
or ( n8389 , n8385 , n8388 );
buf ( n8390 , n4142 );
buf ( n8391 , n5166 );
xor ( n8392 , n8390 , n8391 );
or ( n8393 , n8389 , n8392 );
buf ( n8394 , n4143 );
buf ( n8395 , n5167 );
xor ( n8396 , n8394 , n8395 );
or ( n8397 , n8393 , n8396 );
buf ( n8398 , n4144 );
buf ( n8399 , n5168 );
xor ( n8400 , n8398 , n8399 );
or ( n8401 , n8397 , n8400 );
buf ( n8402 , n4145 );
buf ( n8403 , n5169 );
xor ( n8404 , n8402 , n8403 );
or ( n8405 , n8401 , n8404 );
buf ( n8406 , n4146 );
buf ( n8407 , n5170 );
xor ( n8408 , n8406 , n8407 );
or ( n8409 , n8405 , n8408 );
buf ( n8410 , n4147 );
buf ( n8411 , n5171 );
xor ( n8412 , n8410 , n8411 );
or ( n8413 , n8409 , n8412 );
buf ( n8414 , n4148 );
buf ( n8415 , n5172 );
xor ( n8416 , n8414 , n8415 );
or ( n8417 , n8413 , n8416 );
buf ( n8418 , n4149 );
buf ( n8419 , n5173 );
xor ( n8420 , n8418 , n8419 );
or ( n8421 , n8417 , n8420 );
buf ( n8422 , n4150 );
buf ( n8423 , n5174 );
xor ( n8424 , n8422 , n8423 );
or ( n8425 , n8421 , n8424 );
buf ( n8426 , n4151 );
buf ( n8427 , n5175 );
xor ( n8428 , n8426 , n8427 );
or ( n8429 , n8425 , n8428 );
buf ( n8430 , n4152 );
buf ( n8431 , n5176 );
xor ( n8432 , n8430 , n8431 );
or ( n8433 , n8429 , n8432 );
buf ( n8434 , n4153 );
buf ( n8435 , n5177 );
xor ( n8436 , n8434 , n8435 );
or ( n8437 , n8433 , n8436 );
buf ( n8438 , n4154 );
buf ( n8439 , n5178 );
xor ( n8440 , n8438 , n8439 );
or ( n8441 , n8437 , n8440 );
buf ( n8442 , n4155 );
buf ( n8443 , n5179 );
xor ( n8444 , n8442 , n8443 );
or ( n8445 , n8441 , n8444 );
buf ( n8446 , n4156 );
buf ( n8447 , n5180 );
xor ( n8448 , n8446 , n8447 );
or ( n8449 , n8445 , n8448 );
buf ( n8450 , n4157 );
buf ( n8451 , n5181 );
xor ( n8452 , n8450 , n8451 );
or ( n8453 , n8449 , n8452 );
buf ( n8454 , n4158 );
buf ( n8455 , n5182 );
xor ( n8456 , n8454 , n8455 );
or ( n8457 , n8453 , n8456 );
buf ( n8458 , n4159 );
buf ( n8459 , n5183 );
xor ( n8460 , n8458 , n8459 );
or ( n8461 , n8457 , n8460 );
buf ( n8462 , n4160 );
buf ( n8463 , n5184 );
xor ( n8464 , n8462 , n8463 );
or ( n8465 , n8461 , n8464 );
buf ( n8466 , n4161 );
buf ( n8467 , n5185 );
xor ( n8468 , n8466 , n8467 );
or ( n8469 , n8465 , n8468 );
buf ( n8470 , n4162 );
buf ( n8471 , n5186 );
xor ( n8472 , n8470 , n8471 );
or ( n8473 , n8469 , n8472 );
buf ( n8474 , n4163 );
buf ( n8475 , n5187 );
xor ( n8476 , n8474 , n8475 );
or ( n8477 , n8473 , n8476 );
buf ( n8478 , n4164 );
buf ( n8479 , n5188 );
xor ( n8480 , n8478 , n8479 );
or ( n8481 , n8477 , n8480 );
buf ( n8482 , n4165 );
buf ( n8483 , n5189 );
xor ( n8484 , n8482 , n8483 );
or ( n8485 , n8481 , n8484 );
buf ( n8486 , n4166 );
buf ( n8487 , n5190 );
xor ( n8488 , n8486 , n8487 );
or ( n8489 , n8485 , n8488 );
buf ( n8490 , n4167 );
buf ( n8491 , n5191 );
xor ( n8492 , n8490 , n8491 );
or ( n8493 , n8489 , n8492 );
buf ( n8494 , n4168 );
buf ( n8495 , n5192 );
xor ( n8496 , n8494 , n8495 );
or ( n8497 , n8493 , n8496 );
buf ( n8498 , n4169 );
buf ( n8499 , n5193 );
xor ( n8500 , n8498 , n8499 );
or ( n8501 , n8497 , n8500 );
buf ( n8502 , n4170 );
buf ( n8503 , n5194 );
xor ( n8504 , n8502 , n8503 );
or ( n8505 , n8501 , n8504 );
buf ( n8506 , n4171 );
buf ( n8507 , n5195 );
xor ( n8508 , n8506 , n8507 );
or ( n8509 , n8505 , n8508 );
buf ( n8510 , n4172 );
buf ( n8511 , n5196 );
xor ( n8512 , n8510 , n8511 );
or ( n8513 , n8509 , n8512 );
buf ( n8514 , n4173 );
buf ( n8515 , n5197 );
xor ( n8516 , n8514 , n8515 );
or ( n8517 , n8513 , n8516 );
buf ( n8518 , n4174 );
buf ( n8519 , n5198 );
xor ( n8520 , n8518 , n8519 );
or ( n8521 , n8517 , n8520 );
buf ( n8522 , n4175 );
buf ( n8523 , n5199 );
xor ( n8524 , n8522 , n8523 );
or ( n8525 , n8521 , n8524 );
buf ( n8526 , n4176 );
buf ( n8527 , n5200 );
xor ( n8528 , n8526 , n8527 );
or ( n8529 , n8525 , n8528 );
buf ( n8530 , n4177 );
buf ( n8531 , n5201 );
xor ( n8532 , n8530 , n8531 );
or ( n8533 , n8529 , n8532 );
buf ( n8534 , n4178 );
buf ( n8535 , n5202 );
xor ( n8536 , n8534 , n8535 );
or ( n8537 , n8533 , n8536 );
buf ( n8538 , n4179 );
buf ( n8539 , n5203 );
xor ( n8540 , n8538 , n8539 );
or ( n8541 , n8537 , n8540 );
buf ( n8542 , n4180 );
buf ( n8543 , n5204 );
xor ( n8544 , n8542 , n8543 );
or ( n8545 , n8541 , n8544 );
buf ( n8546 , n4181 );
buf ( n8547 , n5205 );
xor ( n8548 , n8546 , n8547 );
or ( n8549 , n8545 , n8548 );
buf ( n8550 , n4182 );
buf ( n8551 , n5206 );
xor ( n8552 , n8550 , n8551 );
or ( n8553 , n8549 , n8552 );
buf ( n8554 , n4183 );
buf ( n8555 , n5207 );
xor ( n8556 , n8554 , n8555 );
or ( n8557 , n8553 , n8556 );
buf ( n8558 , n4184 );
buf ( n8559 , n5208 );
xor ( n8560 , n8558 , n8559 );
or ( n8561 , n8557 , n8560 );
buf ( n8562 , n4185 );
buf ( n8563 , n5209 );
xor ( n8564 , n8562 , n8563 );
or ( n8565 , n8561 , n8564 );
buf ( n8566 , n4186 );
buf ( n8567 , n5210 );
xor ( n8568 , n8566 , n8567 );
or ( n8569 , n8565 , n8568 );
buf ( n8570 , n4187 );
buf ( n8571 , n5211 );
xor ( n8572 , n8570 , n8571 );
or ( n8573 , n8569 , n8572 );
buf ( n8574 , n4188 );
buf ( n8575 , n5212 );
xor ( n8576 , n8574 , n8575 );
or ( n8577 , n8573 , n8576 );
buf ( n8578 , n4189 );
buf ( n8579 , n5213 );
xor ( n8580 , n8578 , n8579 );
or ( n8581 , n8577 , n8580 );
buf ( n8582 , n4190 );
buf ( n8583 , n5214 );
xor ( n8584 , n8582 , n8583 );
or ( n8585 , n8581 , n8584 );
buf ( n8586 , n4191 );
buf ( n8587 , n5215 );
xor ( n8588 , n8586 , n8587 );
or ( n8589 , n8585 , n8588 );
buf ( n8590 , n4192 );
buf ( n8591 , n5216 );
xor ( n8592 , n8590 , n8591 );
or ( n8593 , n8589 , n8592 );
buf ( n8594 , n4193 );
buf ( n8595 , n5217 );
xor ( n8596 , n8594 , n8595 );
or ( n8597 , n8593 , n8596 );
buf ( n8598 , n4194 );
buf ( n8599 , n5218 );
xor ( n8600 , n8598 , n8599 );
or ( n8601 , n8597 , n8600 );
buf ( n8602 , n4195 );
buf ( n8603 , n5219 );
xor ( n8604 , n8602 , n8603 );
or ( n8605 , n8601 , n8604 );
buf ( n8606 , n4196 );
buf ( n8607 , n5220 );
xor ( n8608 , n8606 , n8607 );
or ( n8609 , n8605 , n8608 );
buf ( n8610 , n4197 );
buf ( n8611 , n5221 );
xor ( n8612 , n8610 , n8611 );
or ( n8613 , n8609 , n8612 );
buf ( n8614 , n4198 );
buf ( n8615 , n5222 );
xor ( n8616 , n8614 , n8615 );
or ( n8617 , n8613 , n8616 );
buf ( n8618 , n4199 );
buf ( n8619 , n5223 );
xor ( n8620 , n8618 , n8619 );
or ( n8621 , n8617 , n8620 );
buf ( n8622 , n4200 );
buf ( n8623 , n5224 );
xor ( n8624 , n8622 , n8623 );
or ( n8625 , n8621 , n8624 );
buf ( n8626 , n4201 );
buf ( n8627 , n5225 );
xor ( n8628 , n8626 , n8627 );
or ( n8629 , n8625 , n8628 );
buf ( n8630 , n4202 );
buf ( n8631 , n5226 );
xor ( n8632 , n8630 , n8631 );
or ( n8633 , n8629 , n8632 );
buf ( n8634 , n4203 );
buf ( n8635 , n5227 );
xor ( n8636 , n8634 , n8635 );
or ( n8637 , n8633 , n8636 );
buf ( n8638 , n4204 );
buf ( n8639 , n5228 );
xor ( n8640 , n8638 , n8639 );
or ( n8641 , n8637 , n8640 );
buf ( n8642 , n4205 );
buf ( n8643 , n5229 );
xor ( n8644 , n8642 , n8643 );
or ( n8645 , n8641 , n8644 );
buf ( n8646 , n4206 );
buf ( n8647 , n5230 );
xor ( n8648 , n8646 , n8647 );
or ( n8649 , n8645 , n8648 );
buf ( n8650 , n4207 );
buf ( n8651 , n5231 );
xor ( n8652 , n8650 , n8651 );
or ( n8653 , n8649 , n8652 );
buf ( n8654 , n4208 );
buf ( n8655 , n5232 );
xor ( n8656 , n8654 , n8655 );
or ( n8657 , n8653 , n8656 );
buf ( n8658 , n4209 );
buf ( n8659 , n5233 );
xor ( n8660 , n8658 , n8659 );
or ( n8661 , n8657 , n8660 );
buf ( n8662 , n4210 );
buf ( n8663 , n5234 );
xor ( n8664 , n8662 , n8663 );
or ( n8665 , n8661 , n8664 );
buf ( n8666 , n4211 );
buf ( n8667 , n5235 );
xor ( n8668 , n8666 , n8667 );
or ( n8669 , n8665 , n8668 );
buf ( n8670 , n4212 );
buf ( n8671 , n5236 );
xor ( n8672 , n8670 , n8671 );
or ( n8673 , n8669 , n8672 );
buf ( n8674 , n4213 );
buf ( n8675 , n5237 );
xor ( n8676 , n8674 , n8675 );
or ( n8677 , n8673 , n8676 );
buf ( n8678 , n4214 );
buf ( n8679 , n5238 );
xor ( n8680 , n8678 , n8679 );
or ( n8681 , n8677 , n8680 );
buf ( n8682 , n4215 );
buf ( n8683 , n5239 );
xor ( n8684 , n8682 , n8683 );
or ( n8685 , n8681 , n8684 );
buf ( n8686 , n4216 );
buf ( n8687 , n5240 );
xor ( n8688 , n8686 , n8687 );
or ( n8689 , n8685 , n8688 );
buf ( n8690 , n4217 );
buf ( n8691 , n5241 );
xor ( n8692 , n8690 , n8691 );
or ( n8693 , n8689 , n8692 );
buf ( n8694 , n4218 );
buf ( n8695 , n5242 );
xor ( n8696 , n8694 , n8695 );
or ( n8697 , n8693 , n8696 );
buf ( n8698 , n4219 );
buf ( n8699 , n5243 );
xor ( n8700 , n8698 , n8699 );
or ( n8701 , n8697 , n8700 );
buf ( n8702 , n4220 );
buf ( n8703 , n5244 );
xor ( n8704 , n8702 , n8703 );
or ( n8705 , n8701 , n8704 );
buf ( n8706 , n4221 );
buf ( n8707 , n5245 );
xor ( n8708 , n8706 , n8707 );
or ( n8709 , n8705 , n8708 );
buf ( n8710 , n4222 );
buf ( n8711 , n5246 );
xor ( n8712 , n8710 , n8711 );
or ( n8713 , n8709 , n8712 );
buf ( n8714 , n4223 );
buf ( n8715 , n5247 );
xor ( n8716 , n8714 , n8715 );
or ( n8717 , n8713 , n8716 );
buf ( n8718 , n4224 );
buf ( n8719 , n5248 );
xor ( n8720 , n8718 , n8719 );
or ( n8721 , n8717 , n8720 );
buf ( n8722 , n4225 );
buf ( n8723 , n5249 );
xor ( n8724 , n8722 , n8723 );
or ( n8725 , n8721 , n8724 );
buf ( n8726 , n4226 );
buf ( n8727 , n5250 );
xor ( n8728 , n8726 , n8727 );
or ( n8729 , n8725 , n8728 );
buf ( n8730 , n4227 );
buf ( n8731 , n5251 );
xor ( n8732 , n8730 , n8731 );
or ( n8733 , n8729 , n8732 );
buf ( n8734 , n4228 );
buf ( n8735 , n5252 );
xor ( n8736 , n8734 , n8735 );
or ( n8737 , n8733 , n8736 );
buf ( n8738 , n4229 );
buf ( n8739 , n5253 );
xor ( n8740 , n8738 , n8739 );
or ( n8741 , n8737 , n8740 );
buf ( n8742 , n4230 );
buf ( n8743 , n5254 );
xor ( n8744 , n8742 , n8743 );
or ( n8745 , n8741 , n8744 );
buf ( n8746 , n4231 );
buf ( n8747 , n5255 );
xor ( n8748 , n8746 , n8747 );
or ( n8749 , n8745 , n8748 );
buf ( n8750 , n4232 );
buf ( n8751 , n5256 );
xor ( n8752 , n8750 , n8751 );
or ( n8753 , n8749 , n8752 );
buf ( n8754 , n4233 );
buf ( n8755 , n5257 );
xor ( n8756 , n8754 , n8755 );
or ( n8757 , n8753 , n8756 );
buf ( n8758 , n4234 );
buf ( n8759 , n5258 );
xor ( n8760 , n8758 , n8759 );
or ( n8761 , n8757 , n8760 );
buf ( n8762 , n4235 );
buf ( n8763 , n5259 );
xor ( n8764 , n8762 , n8763 );
or ( n8765 , n8761 , n8764 );
buf ( n8766 , n4236 );
buf ( n8767 , n5260 );
xor ( n8768 , n8766 , n8767 );
or ( n8769 , n8765 , n8768 );
buf ( n8770 , n4237 );
buf ( n8771 , n5261 );
xor ( n8772 , n8770 , n8771 );
or ( n8773 , n8769 , n8772 );
buf ( n8774 , n4238 );
buf ( n8775 , n5262 );
xor ( n8776 , n8774 , n8775 );
or ( n8777 , n8773 , n8776 );
buf ( n8778 , n4239 );
buf ( n8779 , n5263 );
xor ( n8780 , n8778 , n8779 );
or ( n8781 , n8777 , n8780 );
buf ( n8782 , n4240 );
buf ( n8783 , n5264 );
xor ( n8784 , n8782 , n8783 );
or ( n8785 , n8781 , n8784 );
buf ( n8786 , n4241 );
buf ( n8787 , n5265 );
xor ( n8788 , n8786 , n8787 );
or ( n8789 , n8785 , n8788 );
buf ( n8790 , n4242 );
buf ( n8791 , n5266 );
xor ( n8792 , n8790 , n8791 );
or ( n8793 , n8789 , n8792 );
buf ( n8794 , n4243 );
buf ( n8795 , n5267 );
xor ( n8796 , n8794 , n8795 );
or ( n8797 , n8793 , n8796 );
buf ( n8798 , n4244 );
buf ( n8799 , n5268 );
xor ( n8800 , n8798 , n8799 );
or ( n8801 , n8797 , n8800 );
buf ( n8802 , n4245 );
buf ( n8803 , n5269 );
xor ( n8804 , n8802 , n8803 );
or ( n8805 , n8801 , n8804 );
buf ( n8806 , n4246 );
buf ( n8807 , n5270 );
xor ( n8808 , n8806 , n8807 );
or ( n8809 , n8805 , n8808 );
buf ( n8810 , n4247 );
buf ( n8811 , n5271 );
xor ( n8812 , n8810 , n8811 );
or ( n8813 , n8809 , n8812 );
buf ( n8814 , n4248 );
buf ( n8815 , n5272 );
xor ( n8816 , n8814 , n8815 );
or ( n8817 , n8813 , n8816 );
buf ( n8818 , n4249 );
buf ( n8819 , n5273 );
xor ( n8820 , n8818 , n8819 );
or ( n8821 , n8817 , n8820 );
buf ( n8822 , n4250 );
buf ( n8823 , n5274 );
xor ( n8824 , n8822 , n8823 );
or ( n8825 , n8821 , n8824 );
buf ( n8826 , n4251 );
buf ( n8827 , n5275 );
xor ( n8828 , n8826 , n8827 );
or ( n8829 , n8825 , n8828 );
buf ( n8830 , n4252 );
buf ( n8831 , n5276 );
xor ( n8832 , n8830 , n8831 );
or ( n8833 , n8829 , n8832 );
buf ( n8834 , n4253 );
buf ( n8835 , n5277 );
xor ( n8836 , n8834 , n8835 );
or ( n8837 , n8833 , n8836 );
buf ( n8838 , n4254 );
buf ( n8839 , n5278 );
xor ( n8840 , n8838 , n8839 );
or ( n8841 , n8837 , n8840 );
buf ( n8842 , n4255 );
buf ( n8843 , n5279 );
xor ( n8844 , n8842 , n8843 );
or ( n8845 , n8841 , n8844 );
buf ( n8846 , n4256 );
buf ( n8847 , n5280 );
xor ( n8848 , n8846 , n8847 );
or ( n8849 , n8845 , n8848 );
buf ( n8850 , n4257 );
buf ( n8851 , n5281 );
xor ( n8852 , n8850 , n8851 );
or ( n8853 , n8849 , n8852 );
buf ( n8854 , n4258 );
buf ( n8855 , n5282 );
xor ( n8856 , n8854 , n8855 );
or ( n8857 , n8853 , n8856 );
buf ( n8858 , n4259 );
buf ( n8859 , n5283 );
xor ( n8860 , n8858 , n8859 );
or ( n8861 , n8857 , n8860 );
buf ( n8862 , n4260 );
buf ( n8863 , n5284 );
xor ( n8864 , n8862 , n8863 );
or ( n8865 , n8861 , n8864 );
buf ( n8866 , n4261 );
buf ( n8867 , n5285 );
xor ( n8868 , n8866 , n8867 );
or ( n8869 , n8865 , n8868 );
buf ( n8870 , n4262 );
buf ( n8871 , n5286 );
xor ( n8872 , n8870 , n8871 );
or ( n8873 , n8869 , n8872 );
buf ( n8874 , n4263 );
buf ( n8875 , n5287 );
xor ( n8876 , n8874 , n8875 );
or ( n8877 , n8873 , n8876 );
buf ( n8878 , n4264 );
buf ( n8879 , n5288 );
xor ( n8880 , n8878 , n8879 );
or ( n8881 , n8877 , n8880 );
buf ( n8882 , n4265 );
buf ( n8883 , n5289 );
xor ( n8884 , n8882 , n8883 );
or ( n8885 , n8881 , n8884 );
buf ( n8886 , n4266 );
buf ( n8887 , n5290 );
xor ( n8888 , n8886 , n8887 );
or ( n8889 , n8885 , n8888 );
buf ( n8890 , n4267 );
buf ( n8891 , n5291 );
xor ( n8892 , n8890 , n8891 );
or ( n8893 , n8889 , n8892 );
buf ( n8894 , n4268 );
buf ( n8895 , n5292 );
xor ( n8896 , n8894 , n8895 );
or ( n8897 , n8893 , n8896 );
buf ( n8898 , n4269 );
buf ( n8899 , n5293 );
xor ( n8900 , n8898 , n8899 );
or ( n8901 , n8897 , n8900 );
buf ( n8902 , n4270 );
buf ( n8903 , n5294 );
xor ( n8904 , n8902 , n8903 );
or ( n8905 , n8901 , n8904 );
buf ( n8906 , n4271 );
buf ( n8907 , n5295 );
xor ( n8908 , n8906 , n8907 );
or ( n8909 , n8905 , n8908 );
buf ( n8910 , n4272 );
buf ( n8911 , n5296 );
xor ( n8912 , n8910 , n8911 );
or ( n8913 , n8909 , n8912 );
buf ( n8914 , n4273 );
buf ( n8915 , n5297 );
xor ( n8916 , n8914 , n8915 );
or ( n8917 , n8913 , n8916 );
buf ( n8918 , n4274 );
buf ( n8919 , n5298 );
xor ( n8920 , n8918 , n8919 );
or ( n8921 , n8917 , n8920 );
buf ( n8922 , n4275 );
buf ( n8923 , n5299 );
xor ( n8924 , n8922 , n8923 );
or ( n8925 , n8921 , n8924 );
buf ( n8926 , n4276 );
buf ( n8927 , n5300 );
xor ( n8928 , n8926 , n8927 );
or ( n8929 , n8925 , n8928 );
buf ( n8930 , n4277 );
buf ( n8931 , n5301 );
xor ( n8932 , n8930 , n8931 );
or ( n8933 , n8929 , n8932 );
buf ( n8934 , n4278 );
buf ( n8935 , n5302 );
xor ( n8936 , n8934 , n8935 );
or ( n8937 , n8933 , n8936 );
buf ( n8938 , n4279 );
buf ( n8939 , n5303 );
xor ( n8940 , n8938 , n8939 );
or ( n8941 , n8937 , n8940 );
buf ( n8942 , n4280 );
buf ( n8943 , n5304 );
xor ( n8944 , n8942 , n8943 );
or ( n8945 , n8941 , n8944 );
buf ( n8946 , n4281 );
buf ( n8947 , n5305 );
xor ( n8948 , n8946 , n8947 );
or ( n8949 , n8945 , n8948 );
buf ( n8950 , n4282 );
buf ( n8951 , n5306 );
xor ( n8952 , n8950 , n8951 );
or ( n8953 , n8949 , n8952 );
buf ( n8954 , n4283 );
buf ( n8955 , n5307 );
xor ( n8956 , n8954 , n8955 );
or ( n8957 , n8953 , n8956 );
buf ( n8958 , n4284 );
buf ( n8959 , n5308 );
xor ( n8960 , n8958 , n8959 );
or ( n8961 , n8957 , n8960 );
buf ( n8962 , n4285 );
buf ( n8963 , n5309 );
xor ( n8964 , n8962 , n8963 );
or ( n8965 , n8961 , n8964 );
buf ( n8966 , n4286 );
buf ( n8967 , n5310 );
xor ( n8968 , n8966 , n8967 );
or ( n8969 , n8965 , n8968 );
buf ( n8970 , n4287 );
buf ( n8971 , n5311 );
xor ( n8972 , n8970 , n8971 );
or ( n8973 , n8969 , n8972 );
buf ( n8974 , n4288 );
buf ( n8975 , n5312 );
xor ( n8976 , n8974 , n8975 );
or ( n8977 , n8973 , n8976 );
buf ( n8978 , n4289 );
buf ( n8979 , n5313 );
xor ( n8980 , n8978 , n8979 );
or ( n8981 , n8977 , n8980 );
buf ( n8982 , n4290 );
buf ( n8983 , n5314 );
xor ( n8984 , n8982 , n8983 );
or ( n8985 , n8981 , n8984 );
buf ( n8986 , n4291 );
buf ( n8987 , n5315 );
xor ( n8988 , n8986 , n8987 );
or ( n8989 , n8985 , n8988 );
buf ( n8990 , n4292 );
buf ( n8991 , n5316 );
xor ( n8992 , n8990 , n8991 );
or ( n8993 , n8989 , n8992 );
buf ( n8994 , n4293 );
buf ( n8995 , n5317 );
xor ( n8996 , n8994 , n8995 );
or ( n8997 , n8993 , n8996 );
buf ( n8998 , n4294 );
buf ( n8999 , n5318 );
xor ( n9000 , n8998 , n8999 );
or ( n9001 , n8997 , n9000 );
buf ( n9002 , n4295 );
buf ( n9003 , n5319 );
xor ( n9004 , n9002 , n9003 );
or ( n9005 , n9001 , n9004 );
buf ( n9006 , n4296 );
buf ( n9007 , n5320 );
xor ( n9008 , n9006 , n9007 );
or ( n9009 , n9005 , n9008 );
buf ( n9010 , n4297 );
buf ( n9011 , n5321 );
xor ( n9012 , n9010 , n9011 );
or ( n9013 , n9009 , n9012 );
buf ( n9014 , n4298 );
buf ( n9015 , n5322 );
xor ( n9016 , n9014 , n9015 );
or ( n9017 , n9013 , n9016 );
buf ( n9018 , n4299 );
buf ( n9019 , n5323 );
xor ( n9020 , n9018 , n9019 );
or ( n9021 , n9017 , n9020 );
buf ( n9022 , n4300 );
buf ( n9023 , n5324 );
xor ( n9024 , n9022 , n9023 );
or ( n9025 , n9021 , n9024 );
buf ( n9026 , n4301 );
buf ( n9027 , n5325 );
xor ( n9028 , n9026 , n9027 );
or ( n9029 , n9025 , n9028 );
buf ( n9030 , n4302 );
buf ( n9031 , n5326 );
xor ( n9032 , n9030 , n9031 );
or ( n9033 , n9029 , n9032 );
buf ( n9034 , n4303 );
buf ( n9035 , n5327 );
xor ( n9036 , n9034 , n9035 );
or ( n9037 , n9033 , n9036 );
buf ( n9038 , n4304 );
buf ( n9039 , n5328 );
xor ( n9040 , n9038 , n9039 );
or ( n9041 , n9037 , n9040 );
buf ( n9042 , n4305 );
buf ( n9043 , n5329 );
xor ( n9044 , n9042 , n9043 );
or ( n9045 , n9041 , n9044 );
buf ( n9046 , n4306 );
buf ( n9047 , n5330 );
xor ( n9048 , n9046 , n9047 );
or ( n9049 , n9045 , n9048 );
buf ( n9050 , n4307 );
buf ( n9051 , n5331 );
xor ( n9052 , n9050 , n9051 );
or ( n9053 , n9049 , n9052 );
buf ( n9054 , n4308 );
buf ( n9055 , n5332 );
xor ( n9056 , n9054 , n9055 );
or ( n9057 , n9053 , n9056 );
buf ( n9058 , n4309 );
buf ( n9059 , n5333 );
xor ( n9060 , n9058 , n9059 );
or ( n9061 , n9057 , n9060 );
buf ( n9062 , n4310 );
buf ( n9063 , n5334 );
xor ( n9064 , n9062 , n9063 );
or ( n9065 , n9061 , n9064 );
buf ( n9066 , n4311 );
buf ( n9067 , n5335 );
xor ( n9068 , n9066 , n9067 );
or ( n9069 , n9065 , n9068 );
buf ( n9070 , n4312 );
buf ( n9071 , n5336 );
xor ( n9072 , n9070 , n9071 );
or ( n9073 , n9069 , n9072 );
buf ( n9074 , n4313 );
buf ( n9075 , n5337 );
xor ( n9076 , n9074 , n9075 );
or ( n9077 , n9073 , n9076 );
buf ( n9078 , n4314 );
buf ( n9079 , n5338 );
xor ( n9080 , n9078 , n9079 );
or ( n9081 , n9077 , n9080 );
buf ( n9082 , n4315 );
buf ( n9083 , n5339 );
xor ( n9084 , n9082 , n9083 );
or ( n9085 , n9081 , n9084 );
buf ( n9086 , n4316 );
buf ( n9087 , n5340 );
xor ( n9088 , n9086 , n9087 );
or ( n9089 , n9085 , n9088 );
buf ( n9090 , n4317 );
buf ( n9091 , n5341 );
xor ( n9092 , n9090 , n9091 );
or ( n9093 , n9089 , n9092 );
buf ( n9094 , n4318 );
buf ( n9095 , n5342 );
xor ( n9096 , n9094 , n9095 );
or ( n9097 , n9093 , n9096 );
buf ( n9098 , n4319 );
buf ( n9099 , n5343 );
xor ( n9100 , n9098 , n9099 );
or ( n9101 , n9097 , n9100 );
buf ( n9102 , n4320 );
buf ( n9103 , n5344 );
xor ( n9104 , n9102 , n9103 );
or ( n9105 , n9101 , n9104 );
buf ( n9106 , n4321 );
buf ( n9107 , n5345 );
xor ( n9108 , n9106 , n9107 );
or ( n9109 , n9105 , n9108 );
buf ( n9110 , n4322 );
buf ( n9111 , n5346 );
xor ( n9112 , n9110 , n9111 );
or ( n9113 , n9109 , n9112 );
buf ( n9114 , n4323 );
buf ( n9115 , n5347 );
xor ( n9116 , n9114 , n9115 );
or ( n9117 , n9113 , n9116 );
buf ( n9118 , n4324 );
buf ( n9119 , n5348 );
xor ( n9120 , n9118 , n9119 );
or ( n9121 , n9117 , n9120 );
buf ( n9122 , n4325 );
buf ( n9123 , n5349 );
xor ( n9124 , n9122 , n9123 );
or ( n9125 , n9121 , n9124 );
buf ( n9126 , n4326 );
buf ( n9127 , n5350 );
xor ( n9128 , n9126 , n9127 );
or ( n9129 , n9125 , n9128 );
buf ( n9130 , n4327 );
buf ( n9131 , n5351 );
xor ( n9132 , n9130 , n9131 );
or ( n9133 , n9129 , n9132 );
buf ( n9134 , n4328 );
buf ( n9135 , n5352 );
xor ( n9136 , n9134 , n9135 );
or ( n9137 , n9133 , n9136 );
buf ( n9138 , n4329 );
buf ( n9139 , n5353 );
xor ( n9140 , n9138 , n9139 );
or ( n9141 , n9137 , n9140 );
buf ( n9142 , n4330 );
buf ( n9143 , n5354 );
xor ( n9144 , n9142 , n9143 );
or ( n9145 , n9141 , n9144 );
buf ( n9146 , n4331 );
buf ( n9147 , n5355 );
xor ( n9148 , n9146 , n9147 );
or ( n9149 , n9145 , n9148 );
buf ( n9150 , n4332 );
buf ( n9151 , n5356 );
xor ( n9152 , n9150 , n9151 );
or ( n9153 , n9149 , n9152 );
buf ( n9154 , n4333 );
buf ( n9155 , n5357 );
xor ( n9156 , n9154 , n9155 );
or ( n9157 , n9153 , n9156 );
buf ( n9158 , n4334 );
buf ( n9159 , n5358 );
xor ( n9160 , n9158 , n9159 );
or ( n9161 , n9157 , n9160 );
buf ( n9162 , n4335 );
buf ( n9163 , n5359 );
xor ( n9164 , n9162 , n9163 );
or ( n9165 , n9161 , n9164 );
buf ( n9166 , n4336 );
buf ( n9167 , n5360 );
xor ( n9168 , n9166 , n9167 );
or ( n9169 , n9165 , n9168 );
buf ( n9170 , n4337 );
buf ( n9171 , n5361 );
xor ( n9172 , n9170 , n9171 );
or ( n9173 , n9169 , n9172 );
buf ( n9174 , n4338 );
buf ( n9175 , n5362 );
xor ( n9176 , n9174 , n9175 );
or ( n9177 , n9173 , n9176 );
buf ( n9178 , n4339 );
buf ( n9179 , n5363 );
xor ( n9180 , n9178 , n9179 );
or ( n9181 , n9177 , n9180 );
buf ( n9182 , n4340 );
buf ( n9183 , n5364 );
xor ( n9184 , n9182 , n9183 );
or ( n9185 , n9181 , n9184 );
buf ( n9186 , n4341 );
buf ( n9187 , n5365 );
xor ( n9188 , n9186 , n9187 );
or ( n9189 , n9185 , n9188 );
buf ( n9190 , n4342 );
buf ( n9191 , n5366 );
xor ( n9192 , n9190 , n9191 );
or ( n9193 , n9189 , n9192 );
buf ( n9194 , n4343 );
buf ( n9195 , n5367 );
xor ( n9196 , n9194 , n9195 );
or ( n9197 , n9193 , n9196 );
buf ( n9198 , n4344 );
buf ( n9199 , n5368 );
xor ( n9200 , n9198 , n9199 );
or ( n9201 , n9197 , n9200 );
buf ( n9202 , n4345 );
buf ( n9203 , n5369 );
xor ( n9204 , n9202 , n9203 );
or ( n9205 , n9201 , n9204 );
buf ( n9206 , n4346 );
buf ( n9207 , n5370 );
xor ( n9208 , n9206 , n9207 );
or ( n9209 , n9205 , n9208 );
buf ( n9210 , n4347 );
buf ( n9211 , n5371 );
xor ( n9212 , n9210 , n9211 );
or ( n9213 , n9209 , n9212 );
buf ( n9214 , n4348 );
buf ( n9215 , n5372 );
xor ( n9216 , n9214 , n9215 );
or ( n9217 , n9213 , n9216 );
buf ( n9218 , n4349 );
buf ( n9219 , n5373 );
xor ( n9220 , n9218 , n9219 );
or ( n9221 , n9217 , n9220 );
buf ( n9222 , n4350 );
buf ( n9223 , n5374 );
xor ( n9224 , n9222 , n9223 );
or ( n9225 , n9221 , n9224 );
buf ( n9226 , n4351 );
buf ( n9227 , n5375 );
xor ( n9228 , n9226 , n9227 );
or ( n9229 , n9225 , n9228 );
buf ( n9230 , n4352 );
buf ( n9231 , n5376 );
xor ( n9232 , n9230 , n9231 );
or ( n9233 , n9229 , n9232 );
buf ( n9234 , n4353 );
buf ( n9235 , n5377 );
xor ( n9236 , n9234 , n9235 );
or ( n9237 , n9233 , n9236 );
buf ( n9238 , n4354 );
buf ( n9239 , n5378 );
xor ( n9240 , n9238 , n9239 );
or ( n9241 , n9237 , n9240 );
buf ( n9242 , n4355 );
buf ( n9243 , n5379 );
xor ( n9244 , n9242 , n9243 );
or ( n9245 , n9241 , n9244 );
buf ( n9246 , n4356 );
buf ( n9247 , n5380 );
xor ( n9248 , n9246 , n9247 );
or ( n9249 , n9245 , n9248 );
buf ( n9250 , n4357 );
buf ( n9251 , n5381 );
xor ( n9252 , n9250 , n9251 );
or ( n9253 , n9249 , n9252 );
buf ( n9254 , n4358 );
buf ( n9255 , n5382 );
xor ( n9256 , n9254 , n9255 );
or ( n9257 , n9253 , n9256 );
buf ( n9258 , n4359 );
buf ( n9259 , n5383 );
xor ( n9260 , n9258 , n9259 );
or ( n9261 , n9257 , n9260 );
buf ( n9262 , n4360 );
buf ( n9263 , n5384 );
xor ( n9264 , n9262 , n9263 );
or ( n9265 , n9261 , n9264 );
buf ( n9266 , n4361 );
buf ( n9267 , n5385 );
xor ( n9268 , n9266 , n9267 );
or ( n9269 , n9265 , n9268 );
buf ( n9270 , n4362 );
buf ( n9271 , n5386 );
xor ( n9272 , n9270 , n9271 );
or ( n9273 , n9269 , n9272 );
buf ( n9274 , n4363 );
buf ( n9275 , n5387 );
xor ( n9276 , n9274 , n9275 );
or ( n9277 , n9273 , n9276 );
buf ( n9278 , n4364 );
buf ( n9279 , n5388 );
xor ( n9280 , n9278 , n9279 );
or ( n9281 , n9277 , n9280 );
buf ( n9282 , n4365 );
buf ( n9283 , n5389 );
xor ( n9284 , n9282 , n9283 );
or ( n9285 , n9281 , n9284 );
buf ( n9286 , n4366 );
buf ( n9287 , n5390 );
xor ( n9288 , n9286 , n9287 );
or ( n9289 , n9285 , n9288 );
buf ( n9290 , n4367 );
buf ( n9291 , n5391 );
xor ( n9292 , n9290 , n9291 );
or ( n9293 , n9289 , n9292 );
buf ( n9294 , n4368 );
buf ( n9295 , n5392 );
xor ( n9296 , n9294 , n9295 );
or ( n9297 , n9293 , n9296 );
buf ( n9298 , n4369 );
buf ( n9299 , n5393 );
xor ( n9300 , n9298 , n9299 );
or ( n9301 , n9297 , n9300 );
buf ( n9302 , n4370 );
buf ( n9303 , n5394 );
xor ( n9304 , n9302 , n9303 );
or ( n9305 , n9301 , n9304 );
buf ( n9306 , n4371 );
buf ( n9307 , n5395 );
xor ( n9308 , n9306 , n9307 );
or ( n9309 , n9305 , n9308 );
buf ( n9310 , n4372 );
buf ( n9311 , n5396 );
xor ( n9312 , n9310 , n9311 );
or ( n9313 , n9309 , n9312 );
buf ( n9314 , n4373 );
buf ( n9315 , n5397 );
xor ( n9316 , n9314 , n9315 );
or ( n9317 , n9313 , n9316 );
buf ( n9318 , n4374 );
buf ( n9319 , n5398 );
xor ( n9320 , n9318 , n9319 );
or ( n9321 , n9317 , n9320 );
buf ( n9322 , n4375 );
buf ( n9323 , n5399 );
xor ( n9324 , n9322 , n9323 );
or ( n9325 , n9321 , n9324 );
buf ( n9326 , n4376 );
buf ( n9327 , n5400 );
xor ( n9328 , n9326 , n9327 );
or ( n9329 , n9325 , n9328 );
buf ( n9330 , n4377 );
buf ( n9331 , n5401 );
xor ( n9332 , n9330 , n9331 );
or ( n9333 , n9329 , n9332 );
buf ( n9334 , n4378 );
buf ( n9335 , n5402 );
xor ( n9336 , n9334 , n9335 );
or ( n9337 , n9333 , n9336 );
buf ( n9338 , n4379 );
buf ( n9339 , n5403 );
xor ( n9340 , n9338 , n9339 );
or ( n9341 , n9337 , n9340 );
buf ( n9342 , n4380 );
buf ( n9343 , n5404 );
xor ( n9344 , n9342 , n9343 );
or ( n9345 , n9341 , n9344 );
buf ( n9346 , n4381 );
buf ( n9347 , n5405 );
xor ( n9348 , n9346 , n9347 );
or ( n9349 , n9345 , n9348 );
buf ( n9350 , n4382 );
buf ( n9351 , n5406 );
xor ( n9352 , n9350 , n9351 );
or ( n9353 , n9349 , n9352 );
buf ( n9354 , n4383 );
buf ( n9355 , n5407 );
xor ( n9356 , n9354 , n9355 );
or ( n9357 , n9353 , n9356 );
buf ( n9358 , n4384 );
buf ( n9359 , n5408 );
xor ( n9360 , n9358 , n9359 );
or ( n9361 , n9357 , n9360 );
buf ( n9362 , n4385 );
buf ( n9363 , n5409 );
xor ( n9364 , n9362 , n9363 );
or ( n9365 , n9361 , n9364 );
buf ( n9366 , n4386 );
buf ( n9367 , n5410 );
xor ( n9368 , n9366 , n9367 );
or ( n9369 , n9365 , n9368 );
buf ( n9370 , n4387 );
buf ( n9371 , n5411 );
xor ( n9372 , n9370 , n9371 );
or ( n9373 , n9369 , n9372 );
buf ( n9374 , n4388 );
buf ( n9375 , n5412 );
xor ( n9376 , n9374 , n9375 );
or ( n9377 , n9373 , n9376 );
buf ( n9378 , n4389 );
buf ( n9379 , n5413 );
xor ( n9380 , n9378 , n9379 );
or ( n9381 , n9377 , n9380 );
buf ( n9382 , n4390 );
buf ( n9383 , n5414 );
xor ( n9384 , n9382 , n9383 );
or ( n9385 , n9381 , n9384 );
buf ( n9386 , n4391 );
buf ( n9387 , n5415 );
xor ( n9388 , n9386 , n9387 );
or ( n9389 , n9385 , n9388 );
buf ( n9390 , n4392 );
buf ( n9391 , n5416 );
xor ( n9392 , n9390 , n9391 );
or ( n9393 , n9389 , n9392 );
buf ( n9394 , n4393 );
buf ( n9395 , n5417 );
xor ( n9396 , n9394 , n9395 );
or ( n9397 , n9393 , n9396 );
buf ( n9398 , n4394 );
buf ( n9399 , n5418 );
xor ( n9400 , n9398 , n9399 );
or ( n9401 , n9397 , n9400 );
buf ( n9402 , n4395 );
buf ( n9403 , n5419 );
xor ( n9404 , n9402 , n9403 );
or ( n9405 , n9401 , n9404 );
buf ( n9406 , n4396 );
buf ( n9407 , n5420 );
xor ( n9408 , n9406 , n9407 );
or ( n9409 , n9405 , n9408 );
buf ( n9410 , n4397 );
buf ( n9411 , n5421 );
xor ( n9412 , n9410 , n9411 );
or ( n9413 , n9409 , n9412 );
buf ( n9414 , n4398 );
buf ( n9415 , n5422 );
xor ( n9416 , n9414 , n9415 );
or ( n9417 , n9413 , n9416 );
buf ( n9418 , n4399 );
buf ( n9419 , n5423 );
xor ( n9420 , n9418 , n9419 );
or ( n9421 , n9417 , n9420 );
buf ( n9422 , n4400 );
buf ( n9423 , n5424 );
xor ( n9424 , n9422 , n9423 );
or ( n9425 , n9421 , n9424 );
buf ( n9426 , n4401 );
buf ( n9427 , n5425 );
xor ( n9428 , n9426 , n9427 );
or ( n9429 , n9425 , n9428 );
buf ( n9430 , n4402 );
buf ( n9431 , n5426 );
xor ( n9432 , n9430 , n9431 );
or ( n9433 , n9429 , n9432 );
buf ( n9434 , n4403 );
buf ( n9435 , n5427 );
xor ( n9436 , n9434 , n9435 );
or ( n9437 , n9433 , n9436 );
buf ( n9438 , n4404 );
buf ( n9439 , n5428 );
xor ( n9440 , n9438 , n9439 );
or ( n9441 , n9437 , n9440 );
buf ( n9442 , n4405 );
buf ( n9443 , n5429 );
xor ( n9444 , n9442 , n9443 );
or ( n9445 , n9441 , n9444 );
buf ( n9446 , n4406 );
buf ( n9447 , n5430 );
xor ( n9448 , n9446 , n9447 );
or ( n9449 , n9445 , n9448 );
buf ( n9450 , n4407 );
buf ( n9451 , n5431 );
xor ( n9452 , n9450 , n9451 );
or ( n9453 , n9449 , n9452 );
buf ( n9454 , n4408 );
buf ( n9455 , n5432 );
xor ( n9456 , n9454 , n9455 );
or ( n9457 , n9453 , n9456 );
buf ( n9458 , n4409 );
buf ( n9459 , n5433 );
xor ( n9460 , n9458 , n9459 );
or ( n9461 , n9457 , n9460 );
buf ( n9462 , n4410 );
buf ( n9463 , n5434 );
xor ( n9464 , n9462 , n9463 );
or ( n9465 , n9461 , n9464 );
buf ( n9466 , n4411 );
buf ( n9467 , n5435 );
xor ( n9468 , n9466 , n9467 );
or ( n9469 , n9465 , n9468 );
buf ( n9470 , n4412 );
buf ( n9471 , n5436 );
xor ( n9472 , n9470 , n9471 );
or ( n9473 , n9469 , n9472 );
buf ( n9474 , n4413 );
buf ( n9475 , n5437 );
xor ( n9476 , n9474 , n9475 );
or ( n9477 , n9473 , n9476 );
buf ( n9478 , n4414 );
buf ( n9479 , n5438 );
xor ( n9480 , n9478 , n9479 );
or ( n9481 , n9477 , n9480 );
buf ( n9482 , n4415 );
buf ( n9483 , n5439 );
xor ( n9484 , n9482 , n9483 );
or ( n9485 , n9481 , n9484 );
buf ( n9486 , n4416 );
buf ( n9487 , n5440 );
xor ( n9488 , n9486 , n9487 );
or ( n9489 , n9485 , n9488 );
buf ( n9490 , n4417 );
buf ( n9491 , n5441 );
xor ( n9492 , n9490 , n9491 );
or ( n9493 , n9489 , n9492 );
buf ( n9494 , n4418 );
buf ( n9495 , n5442 );
xor ( n9496 , n9494 , n9495 );
or ( n9497 , n9493 , n9496 );
buf ( n9498 , n4419 );
buf ( n9499 , n5443 );
xor ( n9500 , n9498 , n9499 );
or ( n9501 , n9497 , n9500 );
buf ( n9502 , n4420 );
buf ( n9503 , n5444 );
xor ( n9504 , n9502 , n9503 );
or ( n9505 , n9501 , n9504 );
buf ( n9506 , n4421 );
buf ( n9507 , n5445 );
xor ( n9508 , n9506 , n9507 );
or ( n9509 , n9505 , n9508 );
buf ( n9510 , n4422 );
buf ( n9511 , n5446 );
xor ( n9512 , n9510 , n9511 );
or ( n9513 , n9509 , n9512 );
buf ( n9514 , n4423 );
buf ( n9515 , n5447 );
xor ( n9516 , n9514 , n9515 );
or ( n9517 , n9513 , n9516 );
buf ( n9518 , n4424 );
buf ( n9519 , n5448 );
xor ( n9520 , n9518 , n9519 );
or ( n9521 , n9517 , n9520 );
buf ( n9522 , n4425 );
buf ( n9523 , n5449 );
xor ( n9524 , n9522 , n9523 );
or ( n9525 , n9521 , n9524 );
buf ( n9526 , n4426 );
buf ( n9527 , n5450 );
xor ( n9528 , n9526 , n9527 );
or ( n9529 , n9525 , n9528 );
buf ( n9530 , n4427 );
buf ( n9531 , n5451 );
xor ( n9532 , n9530 , n9531 );
or ( n9533 , n9529 , n9532 );
buf ( n9534 , n4428 );
buf ( n9535 , n5452 );
xor ( n9536 , n9534 , n9535 );
or ( n9537 , n9533 , n9536 );
buf ( n9538 , n4429 );
buf ( n9539 , n5453 );
xor ( n9540 , n9538 , n9539 );
or ( n9541 , n9537 , n9540 );
buf ( n9542 , n4430 );
buf ( n9543 , n5454 );
xor ( n9544 , n9542 , n9543 );
or ( n9545 , n9541 , n9544 );
buf ( n9546 , n4431 );
buf ( n9547 , n5455 );
xor ( n9548 , n9546 , n9547 );
or ( n9549 , n9545 , n9548 );
buf ( n9550 , n4432 );
buf ( n9551 , n5456 );
xor ( n9552 , n9550 , n9551 );
or ( n9553 , n9549 , n9552 );
buf ( n9554 , n4433 );
buf ( n9555 , n5457 );
xor ( n9556 , n9554 , n9555 );
or ( n9557 , n9553 , n9556 );
buf ( n9558 , n4434 );
buf ( n9559 , n5458 );
xor ( n9560 , n9558 , n9559 );
or ( n9561 , n9557 , n9560 );
buf ( n9562 , n4435 );
buf ( n9563 , n5459 );
xor ( n9564 , n9562 , n9563 );
or ( n9565 , n9561 , n9564 );
buf ( n9566 , n4436 );
buf ( n9567 , n5460 );
xor ( n9568 , n9566 , n9567 );
or ( n9569 , n9565 , n9568 );
buf ( n9570 , n4437 );
buf ( n9571 , n5461 );
xor ( n9572 , n9570 , n9571 );
or ( n9573 , n9569 , n9572 );
buf ( n9574 , n4438 );
buf ( n9575 , n5462 );
xor ( n9576 , n9574 , n9575 );
or ( n9577 , n9573 , n9576 );
buf ( n9578 , n4439 );
buf ( n9579 , n5463 );
xor ( n9580 , n9578 , n9579 );
or ( n9581 , n9577 , n9580 );
buf ( n9582 , n4440 );
buf ( n9583 , n5464 );
xor ( n9584 , n9582 , n9583 );
or ( n9585 , n9581 , n9584 );
buf ( n9586 , n4441 );
buf ( n9587 , n5465 );
xor ( n9588 , n9586 , n9587 );
or ( n9589 , n9585 , n9588 );
buf ( n9590 , n4442 );
buf ( n9591 , n5466 );
xor ( n9592 , n9590 , n9591 );
or ( n9593 , n9589 , n9592 );
buf ( n9594 , n4443 );
buf ( n9595 , n5467 );
xor ( n9596 , n9594 , n9595 );
or ( n9597 , n9593 , n9596 );
buf ( n9598 , n4444 );
buf ( n9599 , n5468 );
xor ( n9600 , n9598 , n9599 );
or ( n9601 , n9597 , n9600 );
buf ( n9602 , n4445 );
buf ( n9603 , n5469 );
xor ( n9604 , n9602 , n9603 );
or ( n9605 , n9601 , n9604 );
buf ( n9606 , n4446 );
buf ( n9607 , n5470 );
xor ( n9608 , n9606 , n9607 );
or ( n9609 , n9605 , n9608 );
buf ( n9610 , n4447 );
buf ( n9611 , n5471 );
xor ( n9612 , n9610 , n9611 );
or ( n9613 , n9609 , n9612 );
buf ( n9614 , n4448 );
buf ( n9615 , n5472 );
xor ( n9616 , n9614 , n9615 );
or ( n9617 , n9613 , n9616 );
buf ( n9618 , n4449 );
buf ( n9619 , n5473 );
xor ( n9620 , n9618 , n9619 );
or ( n9621 , n9617 , n9620 );
buf ( n9622 , n4450 );
buf ( n9623 , n5474 );
xor ( n9624 , n9622 , n9623 );
or ( n9625 , n9621 , n9624 );
buf ( n9626 , n4451 );
buf ( n9627 , n5475 );
xor ( n9628 , n9626 , n9627 );
or ( n9629 , n9625 , n9628 );
buf ( n9630 , n4452 );
buf ( n9631 , n5476 );
xor ( n9632 , n9630 , n9631 );
or ( n9633 , n9629 , n9632 );
buf ( n9634 , n4453 );
buf ( n9635 , n5477 );
xor ( n9636 , n9634 , n9635 );
or ( n9637 , n9633 , n9636 );
buf ( n9638 , n4454 );
buf ( n9639 , n5478 );
xor ( n9640 , n9638 , n9639 );
or ( n9641 , n9637 , n9640 );
buf ( n9642 , n4455 );
buf ( n9643 , n5479 );
xor ( n9644 , n9642 , n9643 );
or ( n9645 , n9641 , n9644 );
buf ( n9646 , n4456 );
buf ( n9647 , n5480 );
xor ( n9648 , n9646 , n9647 );
or ( n9649 , n9645 , n9648 );
buf ( n9650 , n4457 );
buf ( n9651 , n5481 );
xor ( n9652 , n9650 , n9651 );
or ( n9653 , n9649 , n9652 );
buf ( n9654 , n4458 );
buf ( n9655 , n5482 );
xor ( n9656 , n9654 , n9655 );
or ( n9657 , n9653 , n9656 );
buf ( n9658 , n4459 );
buf ( n9659 , n5483 );
xor ( n9660 , n9658 , n9659 );
or ( n9661 , n9657 , n9660 );
buf ( n9662 , n4460 );
buf ( n9663 , n5484 );
xor ( n9664 , n9662 , n9663 );
or ( n9665 , n9661 , n9664 );
buf ( n9666 , n4461 );
buf ( n9667 , n5485 );
xor ( n9668 , n9666 , n9667 );
or ( n9669 , n9665 , n9668 );
buf ( n9670 , n4462 );
buf ( n9671 , n5486 );
xor ( n9672 , n9670 , n9671 );
or ( n9673 , n9669 , n9672 );
buf ( n9674 , n4463 );
buf ( n9675 , n5487 );
xor ( n9676 , n9674 , n9675 );
or ( n9677 , n9673 , n9676 );
buf ( n9678 , n4464 );
buf ( n9679 , n5488 );
xor ( n9680 , n9678 , n9679 );
or ( n9681 , n9677 , n9680 );
buf ( n9682 , n4465 );
buf ( n9683 , n5489 );
xor ( n9684 , n9682 , n9683 );
or ( n9685 , n9681 , n9684 );
buf ( n9686 , n4466 );
buf ( n9687 , n5490 );
xor ( n9688 , n9686 , n9687 );
or ( n9689 , n9685 , n9688 );
buf ( n9690 , n4467 );
buf ( n9691 , n5491 );
xor ( n9692 , n9690 , n9691 );
or ( n9693 , n9689 , n9692 );
buf ( n9694 , n4468 );
buf ( n9695 , n5492 );
xor ( n9696 , n9694 , n9695 );
or ( n9697 , n9693 , n9696 );
buf ( n9698 , n4469 );
buf ( n9699 , n5493 );
xor ( n9700 , n9698 , n9699 );
or ( n9701 , n9697 , n9700 );
buf ( n9702 , n4470 );
buf ( n9703 , n5494 );
xor ( n9704 , n9702 , n9703 );
or ( n9705 , n9701 , n9704 );
buf ( n9706 , n4471 );
buf ( n9707 , n5495 );
xor ( n9708 , n9706 , n9707 );
or ( n9709 , n9705 , n9708 );
buf ( n9710 , n4472 );
buf ( n9711 , n5496 );
xor ( n9712 , n9710 , n9711 );
or ( n9713 , n9709 , n9712 );
buf ( n9714 , n4473 );
buf ( n9715 , n5497 );
xor ( n9716 , n9714 , n9715 );
or ( n9717 , n9713 , n9716 );
buf ( n9718 , n4474 );
buf ( n9719 , n5498 );
xor ( n9720 , n9718 , n9719 );
or ( n9721 , n9717 , n9720 );
buf ( n9722 , n4475 );
buf ( n9723 , n5499 );
xor ( n9724 , n9722 , n9723 );
or ( n9725 , n9721 , n9724 );
buf ( n9726 , n4476 );
buf ( n9727 , n5500 );
xor ( n9728 , n9726 , n9727 );
or ( n9729 , n9725 , n9728 );
buf ( n9730 , n4477 );
buf ( n9731 , n5501 );
xor ( n9732 , n9730 , n9731 );
or ( n9733 , n9729 , n9732 );
buf ( n9734 , n4478 );
buf ( n9735 , n5502 );
xor ( n9736 , n9734 , n9735 );
or ( n9737 , n9733 , n9736 );
buf ( n9738 , n4479 );
buf ( n9739 , n5503 );
xor ( n9740 , n9738 , n9739 );
or ( n9741 , n9737 , n9740 );
buf ( n9742 , n4480 );
buf ( n9743 , n5504 );
xor ( n9744 , n9742 , n9743 );
or ( n9745 , n9741 , n9744 );
buf ( n9746 , n4481 );
buf ( n9747 , n5505 );
xor ( n9748 , n9746 , n9747 );
or ( n9749 , n9745 , n9748 );
buf ( n9750 , n4482 );
buf ( n9751 , n5506 );
xor ( n9752 , n9750 , n9751 );
or ( n9753 , n9749 , n9752 );
buf ( n9754 , n4483 );
buf ( n9755 , n5507 );
xor ( n9756 , n9754 , n9755 );
or ( n9757 , n9753 , n9756 );
buf ( n9758 , n4484 );
buf ( n9759 , n5508 );
xor ( n9760 , n9758 , n9759 );
or ( n9761 , n9757 , n9760 );
buf ( n9762 , n4485 );
buf ( n9763 , n5509 );
xor ( n9764 , n9762 , n9763 );
or ( n9765 , n9761 , n9764 );
buf ( n9766 , n4486 );
buf ( n9767 , n5510 );
xor ( n9768 , n9766 , n9767 );
or ( n9769 , n9765 , n9768 );
buf ( n9770 , n4487 );
buf ( n9771 , n5511 );
xor ( n9772 , n9770 , n9771 );
or ( n9773 , n9769 , n9772 );
buf ( n9774 , n4488 );
buf ( n9775 , n5512 );
xor ( n9776 , n9774 , n9775 );
or ( n9777 , n9773 , n9776 );
buf ( n9778 , n4489 );
buf ( n9779 , n5513 );
xor ( n9780 , n9778 , n9779 );
or ( n9781 , n9777 , n9780 );
buf ( n9782 , n4490 );
buf ( n9783 , n5514 );
xor ( n9784 , n9782 , n9783 );
or ( n9785 , n9781 , n9784 );
buf ( n9786 , n4491 );
buf ( n9787 , n5515 );
xor ( n9788 , n9786 , n9787 );
or ( n9789 , n9785 , n9788 );
buf ( n9790 , n4492 );
buf ( n9791 , n5516 );
xor ( n9792 , n9790 , n9791 );
or ( n9793 , n9789 , n9792 );
buf ( n9794 , n4493 );
buf ( n9795 , n5517 );
xor ( n9796 , n9794 , n9795 );
or ( n9797 , n9793 , n9796 );
buf ( n9798 , n4494 );
buf ( n9799 , n5518 );
xor ( n9800 , n9798 , n9799 );
or ( n9801 , n9797 , n9800 );
buf ( n9802 , n4495 );
buf ( n9803 , n5519 );
xor ( n9804 , n9802 , n9803 );
or ( n9805 , n9801 , n9804 );
buf ( n9806 , n4496 );
buf ( n9807 , n5520 );
xor ( n9808 , n9806 , n9807 );
or ( n9809 , n9805 , n9808 );
buf ( n9810 , n4497 );
buf ( n9811 , n5521 );
xor ( n9812 , n9810 , n9811 );
or ( n9813 , n9809 , n9812 );
buf ( n9814 , n4498 );
buf ( n9815 , n5522 );
xor ( n9816 , n9814 , n9815 );
or ( n9817 , n9813 , n9816 );
buf ( n9818 , n4499 );
buf ( n9819 , n5523 );
xor ( n9820 , n9818 , n9819 );
or ( n9821 , n9817 , n9820 );
buf ( n9822 , n4500 );
buf ( n9823 , n5524 );
xor ( n9824 , n9822 , n9823 );
or ( n9825 , n9821 , n9824 );
buf ( n9826 , n4501 );
buf ( n9827 , n5525 );
xor ( n9828 , n9826 , n9827 );
or ( n9829 , n9825 , n9828 );
buf ( n9830 , n4502 );
buf ( n9831 , n5526 );
xor ( n9832 , n9830 , n9831 );
or ( n9833 , n9829 , n9832 );
buf ( n9834 , n4503 );
buf ( n9835 , n5527 );
xor ( n9836 , n9834 , n9835 );
or ( n9837 , n9833 , n9836 );
buf ( n9838 , n4504 );
buf ( n9839 , n5528 );
xor ( n9840 , n9838 , n9839 );
or ( n9841 , n9837 , n9840 );
buf ( n9842 , n4505 );
buf ( n9843 , n5529 );
xor ( n9844 , n9842 , n9843 );
or ( n9845 , n9841 , n9844 );
buf ( n9846 , n4506 );
buf ( n9847 , n5530 );
xor ( n9848 , n9846 , n9847 );
or ( n9849 , n9845 , n9848 );
buf ( n9850 , n4507 );
buf ( n9851 , n5531 );
xor ( n9852 , n9850 , n9851 );
or ( n9853 , n9849 , n9852 );
buf ( n9854 , n4508 );
buf ( n9855 , n5532 );
xor ( n9856 , n9854 , n9855 );
or ( n9857 , n9853 , n9856 );
buf ( n9858 , n4509 );
buf ( n9859 , n5533 );
xor ( n9860 , n9858 , n9859 );
or ( n9861 , n9857 , n9860 );
buf ( n9862 , n4510 );
buf ( n9863 , n5534 );
xor ( n9864 , n9862 , n9863 );
or ( n9865 , n9861 , n9864 );
buf ( n9866 , n4511 );
buf ( n9867 , n5535 );
xor ( n9868 , n9866 , n9867 );
or ( n9869 , n9865 , n9868 );
buf ( n9870 , n4512 );
buf ( n9871 , n5536 );
xor ( n9872 , n9870 , n9871 );
or ( n9873 , n9869 , n9872 );
buf ( n9874 , n4513 );
buf ( n9875 , n5537 );
xor ( n9876 , n9874 , n9875 );
or ( n9877 , n9873 , n9876 );
buf ( n9878 , n4514 );
buf ( n9879 , n5538 );
xor ( n9880 , n9878 , n9879 );
or ( n9881 , n9877 , n9880 );
buf ( n9882 , n4515 );
buf ( n9883 , n5539 );
xor ( n9884 , n9882 , n9883 );
or ( n9885 , n9881 , n9884 );
buf ( n9886 , n4516 );
buf ( n9887 , n5540 );
xor ( n9888 , n9886 , n9887 );
or ( n9889 , n9885 , n9888 );
buf ( n9890 , n4517 );
buf ( n9891 , n5541 );
xor ( n9892 , n9890 , n9891 );
or ( n9893 , n9889 , n9892 );
buf ( n9894 , n4518 );
buf ( n9895 , n5542 );
xor ( n9896 , n9894 , n9895 );
or ( n9897 , n9893 , n9896 );
buf ( n9898 , n4519 );
buf ( n9899 , n5543 );
xor ( n9900 , n9898 , n9899 );
or ( n9901 , n9897 , n9900 );
buf ( n9902 , n4520 );
buf ( n9903 , n5544 );
xor ( n9904 , n9902 , n9903 );
or ( n9905 , n9901 , n9904 );
buf ( n9906 , n4521 );
buf ( n9907 , n5545 );
xor ( n9908 , n9906 , n9907 );
or ( n9909 , n9905 , n9908 );
buf ( n9910 , n4522 );
buf ( n9911 , n5546 );
xor ( n9912 , n9910 , n9911 );
or ( n9913 , n9909 , n9912 );
buf ( n9914 , n4523 );
buf ( n9915 , n5547 );
xor ( n9916 , n9914 , n9915 );
or ( n9917 , n9913 , n9916 );
buf ( n9918 , n4524 );
buf ( n9919 , n5548 );
xor ( n9920 , n9918 , n9919 );
or ( n9921 , n9917 , n9920 );
buf ( n9922 , n4525 );
buf ( n9923 , n5549 );
xor ( n9924 , n9922 , n9923 );
or ( n9925 , n9921 , n9924 );
buf ( n9926 , n4526 );
buf ( n9927 , n5550 );
xor ( n9928 , n9926 , n9927 );
or ( n9929 , n9925 , n9928 );
buf ( n9930 , n4527 );
buf ( n9931 , n5551 );
xor ( n9932 , n9930 , n9931 );
or ( n9933 , n9929 , n9932 );
buf ( n9934 , n4528 );
buf ( n9935 , n5552 );
xor ( n9936 , n9934 , n9935 );
or ( n9937 , n9933 , n9936 );
buf ( n9938 , n4529 );
buf ( n9939 , n5553 );
xor ( n9940 , n9938 , n9939 );
or ( n9941 , n9937 , n9940 );
buf ( n9942 , n4530 );
buf ( n9943 , n5554 );
xor ( n9944 , n9942 , n9943 );
or ( n9945 , n9941 , n9944 );
buf ( n9946 , n4531 );
buf ( n9947 , n5555 );
xor ( n9948 , n9946 , n9947 );
or ( n9949 , n9945 , n9948 );
buf ( n9950 , n4532 );
buf ( n9951 , n5556 );
xor ( n9952 , n9950 , n9951 );
or ( n9953 , n9949 , n9952 );
buf ( n9954 , n4533 );
buf ( n9955 , n5557 );
xor ( n9956 , n9954 , n9955 );
or ( n9957 , n9953 , n9956 );
buf ( n9958 , n4534 );
buf ( n9959 , n5558 );
xor ( n9960 , n9958 , n9959 );
or ( n9961 , n9957 , n9960 );
buf ( n9962 , n4535 );
buf ( n9963 , n5559 );
xor ( n9964 , n9962 , n9963 );
or ( n9965 , n9961 , n9964 );
buf ( n9966 , n4536 );
buf ( n9967 , n5560 );
xor ( n9968 , n9966 , n9967 );
or ( n9969 , n9965 , n9968 );
buf ( n9970 , n4537 );
buf ( n9971 , n5561 );
xor ( n9972 , n9970 , n9971 );
or ( n9973 , n9969 , n9972 );
buf ( n9974 , n4538 );
buf ( n9975 , n5562 );
xor ( n9976 , n9974 , n9975 );
or ( n9977 , n9973 , n9976 );
buf ( n9978 , n4539 );
buf ( n9979 , n5563 );
xor ( n9980 , n9978 , n9979 );
or ( n9981 , n9977 , n9980 );
buf ( n9982 , n4540 );
buf ( n9983 , n5564 );
xor ( n9984 , n9982 , n9983 );
or ( n9985 , n9981 , n9984 );
buf ( n9986 , n4541 );
buf ( n9987 , n5565 );
xor ( n9988 , n9986 , n9987 );
or ( n9989 , n9985 , n9988 );
buf ( n9990 , n4542 );
buf ( n9991 , n5566 );
xor ( n9992 , n9990 , n9991 );
or ( n9993 , n9989 , n9992 );
buf ( n9994 , n4543 );
buf ( n9995 , n5567 );
xor ( n9996 , n9994 , n9995 );
or ( n9997 , n9993 , n9996 );
buf ( n9998 , n4544 );
buf ( n9999 , n5568 );
xor ( n10000 , n9998 , n9999 );
or ( n10001 , n9997 , n10000 );
buf ( n10002 , n4545 );
buf ( n10003 , n5569 );
xor ( n10004 , n10002 , n10003 );
or ( n10005 , n10001 , n10004 );
buf ( n10006 , n4546 );
buf ( n10007 , n5570 );
xor ( n10008 , n10006 , n10007 );
or ( n10009 , n10005 , n10008 );
buf ( n10010 , n4547 );
buf ( n10011 , n5571 );
xor ( n10012 , n10010 , n10011 );
or ( n10013 , n10009 , n10012 );
buf ( n10014 , n4548 );
buf ( n10015 , n5572 );
xor ( n10016 , n10014 , n10015 );
or ( n10017 , n10013 , n10016 );
buf ( n10018 , n4549 );
buf ( n10019 , n5573 );
xor ( n10020 , n10018 , n10019 );
or ( n10021 , n10017 , n10020 );
buf ( n10022 , n4550 );
buf ( n10023 , n5574 );
xor ( n10024 , n10022 , n10023 );
or ( n10025 , n10021 , n10024 );
buf ( n10026 , n4551 );
buf ( n10027 , n5575 );
xor ( n10028 , n10026 , n10027 );
or ( n10029 , n10025 , n10028 );
buf ( n10030 , n4552 );
buf ( n10031 , n5576 );
xor ( n10032 , n10030 , n10031 );
or ( n10033 , n10029 , n10032 );
buf ( n10034 , n4553 );
buf ( n10035 , n5577 );
xor ( n10036 , n10034 , n10035 );
or ( n10037 , n10033 , n10036 );
buf ( n10038 , n4554 );
buf ( n10039 , n5578 );
xor ( n10040 , n10038 , n10039 );
or ( n10041 , n10037 , n10040 );
buf ( n10042 , n4555 );
buf ( n10043 , n5579 );
xor ( n10044 , n10042 , n10043 );
or ( n10045 , n10041 , n10044 );
buf ( n10046 , n4556 );
buf ( n10047 , n5580 );
xor ( n10048 , n10046 , n10047 );
or ( n10049 , n10045 , n10048 );
buf ( n10050 , n4557 );
buf ( n10051 , n5581 );
xor ( n10052 , n10050 , n10051 );
or ( n10053 , n10049 , n10052 );
buf ( n10054 , n4558 );
buf ( n10055 , n5582 );
xor ( n10056 , n10054 , n10055 );
or ( n10057 , n10053 , n10056 );
buf ( n10058 , n4559 );
buf ( n10059 , n5583 );
xor ( n10060 , n10058 , n10059 );
or ( n10061 , n10057 , n10060 );
buf ( n10062 , n4560 );
buf ( n10063 , n5584 );
xor ( n10064 , n10062 , n10063 );
or ( n10065 , n10061 , n10064 );
buf ( n10066 , n4561 );
buf ( n10067 , n5585 );
xor ( n10068 , n10066 , n10067 );
or ( n10069 , n10065 , n10068 );
buf ( n10070 , n4562 );
buf ( n10071 , n5586 );
xor ( n10072 , n10070 , n10071 );
or ( n10073 , n10069 , n10072 );
buf ( n10074 , n4563 );
buf ( n10075 , n5587 );
xor ( n10076 , n10074 , n10075 );
or ( n10077 , n10073 , n10076 );
buf ( n10078 , n4564 );
buf ( n10079 , n5588 );
xor ( n10080 , n10078 , n10079 );
or ( n10081 , n10077 , n10080 );
buf ( n10082 , n4565 );
buf ( n10083 , n5589 );
xor ( n10084 , n10082 , n10083 );
or ( n10085 , n10081 , n10084 );
buf ( n10086 , n4566 );
buf ( n10087 , n5590 );
xor ( n10088 , n10086 , n10087 );
or ( n10089 , n10085 , n10088 );
buf ( n10090 , n4567 );
buf ( n10091 , n5591 );
xor ( n10092 , n10090 , n10091 );
or ( n10093 , n10089 , n10092 );
buf ( n10094 , n4568 );
buf ( n10095 , n5592 );
xor ( n10096 , n10094 , n10095 );
or ( n10097 , n10093 , n10096 );
buf ( n10098 , n4569 );
buf ( n10099 , n5593 );
xor ( n10100 , n10098 , n10099 );
or ( n10101 , n10097 , n10100 );
buf ( n10102 , n4570 );
buf ( n10103 , n5594 );
xor ( n10104 , n10102 , n10103 );
or ( n10105 , n10101 , n10104 );
buf ( n10106 , n4571 );
buf ( n10107 , n5595 );
xor ( n10108 , n10106 , n10107 );
or ( n10109 , n10105 , n10108 );
buf ( n10110 , n4572 );
buf ( n10111 , n5596 );
xor ( n10112 , n10110 , n10111 );
or ( n10113 , n10109 , n10112 );
buf ( n10114 , n4573 );
buf ( n10115 , n5597 );
xor ( n10116 , n10114 , n10115 );
or ( n10117 , n10113 , n10116 );
buf ( n10118 , n4574 );
buf ( n10119 , n5598 );
xor ( n10120 , n10118 , n10119 );
or ( n10121 , n10117 , n10120 );
buf ( n10122 , n4575 );
buf ( n10123 , n5599 );
xor ( n10124 , n10122 , n10123 );
or ( n10125 , n10121 , n10124 );
buf ( n10126 , n4576 );
buf ( n10127 , n5600 );
xor ( n10128 , n10126 , n10127 );
or ( n10129 , n10125 , n10128 );
buf ( n10130 , n4577 );
buf ( n10131 , n5601 );
xor ( n10132 , n10130 , n10131 );
or ( n10133 , n10129 , n10132 );
buf ( n10134 , n4578 );
buf ( n10135 , n5602 );
xor ( n10136 , n10134 , n10135 );
or ( n10137 , n10133 , n10136 );
buf ( n10138 , n4579 );
buf ( n10139 , n5603 );
xor ( n10140 , n10138 , n10139 );
or ( n10141 , n10137 , n10140 );
buf ( n10142 , n4580 );
buf ( n10143 , n5604 );
xor ( n10144 , n10142 , n10143 );
or ( n10145 , n10141 , n10144 );
buf ( n10146 , n4581 );
buf ( n10147 , n5605 );
xor ( n10148 , n10146 , n10147 );
or ( n10149 , n10145 , n10148 );
buf ( n10150 , n4582 );
buf ( n10151 , n5606 );
xor ( n10152 , n10150 , n10151 );
or ( n10153 , n10149 , n10152 );
buf ( n10154 , n4583 );
buf ( n10155 , n5607 );
xor ( n10156 , n10154 , n10155 );
or ( n10157 , n10153 , n10156 );
buf ( n10158 , n4584 );
buf ( n10159 , n5608 );
xor ( n10160 , n10158 , n10159 );
or ( n10161 , n10157 , n10160 );
buf ( n10162 , n4585 );
buf ( n10163 , n5609 );
xor ( n10164 , n10162 , n10163 );
or ( n10165 , n10161 , n10164 );
buf ( n10166 , n4586 );
buf ( n10167 , n5610 );
xor ( n10168 , n10166 , n10167 );
or ( n10169 , n10165 , n10168 );
buf ( n10170 , n4587 );
buf ( n10171 , n5611 );
xor ( n10172 , n10170 , n10171 );
or ( n10173 , n10169 , n10172 );
buf ( n10174 , n4588 );
buf ( n10175 , n5612 );
xor ( n10176 , n10174 , n10175 );
or ( n10177 , n10173 , n10176 );
buf ( n10178 , n4589 );
buf ( n10179 , n5613 );
xor ( n10180 , n10178 , n10179 );
or ( n10181 , n10177 , n10180 );
buf ( n10182 , n4590 );
buf ( n10183 , n5614 );
xor ( n10184 , n10182 , n10183 );
or ( n10185 , n10181 , n10184 );
buf ( n10186 , n4591 );
buf ( n10187 , n5615 );
xor ( n10188 , n10186 , n10187 );
or ( n10189 , n10185 , n10188 );
buf ( n10190 , n4592 );
buf ( n10191 , n5616 );
xor ( n10192 , n10190 , n10191 );
or ( n10193 , n10189 , n10192 );
buf ( n10194 , n4593 );
buf ( n10195 , n5617 );
xor ( n10196 , n10194 , n10195 );
or ( n10197 , n10193 , n10196 );
buf ( n10198 , n4594 );
buf ( n10199 , n5618 );
xor ( n10200 , n10198 , n10199 );
or ( n10201 , n10197 , n10200 );
buf ( n10202 , n4595 );
buf ( n10203 , n5619 );
xor ( n10204 , n10202 , n10203 );
or ( n10205 , n10201 , n10204 );
buf ( n10206 , n4596 );
buf ( n10207 , n5620 );
xor ( n10208 , n10206 , n10207 );
or ( n10209 , n10205 , n10208 );
buf ( n10210 , n4597 );
buf ( n10211 , n5621 );
xor ( n10212 , n10210 , n10211 );
or ( n10213 , n10209 , n10212 );
buf ( n10214 , n4598 );
buf ( n10215 , n5622 );
xor ( n10216 , n10214 , n10215 );
or ( n10217 , n10213 , n10216 );
buf ( n10218 , n4599 );
buf ( n10219 , n5623 );
xor ( n10220 , n10218 , n10219 );
or ( n10221 , n10217 , n10220 );
buf ( n10222 , n4600 );
buf ( n10223 , n5624 );
xor ( n10224 , n10222 , n10223 );
or ( n10225 , n10221 , n10224 );
buf ( n10226 , n4601 );
buf ( n10227 , n5625 );
xor ( n10228 , n10226 , n10227 );
or ( n10229 , n10225 , n10228 );
buf ( n10230 , n4602 );
buf ( n10231 , n5626 );
xor ( n10232 , n10230 , n10231 );
or ( n10233 , n10229 , n10232 );
buf ( n10234 , n4603 );
buf ( n10235 , n5627 );
xor ( n10236 , n10234 , n10235 );
or ( n10237 , n10233 , n10236 );
buf ( n10238 , n4604 );
buf ( n10239 , n5628 );
xor ( n10240 , n10238 , n10239 );
or ( n10241 , n10237 , n10240 );
buf ( n10242 , n4605 );
buf ( n10243 , n5629 );
xor ( n10244 , n10242 , n10243 );
or ( n10245 , n10241 , n10244 );
buf ( n10246 , n4606 );
buf ( n10247 , n5630 );
xor ( n10248 , n10246 , n10247 );
or ( n10249 , n10245 , n10248 );
buf ( n10250 , n4607 );
buf ( n10251 , n5631 );
xor ( n10252 , n10250 , n10251 );
or ( n10253 , n10249 , n10252 );
buf ( n10254 , n4608 );
buf ( n10255 , n5632 );
xor ( n10256 , n10254 , n10255 );
or ( n10257 , n10253 , n10256 );
buf ( n10258 , n4609 );
buf ( n10259 , n5633 );
xor ( n10260 , n10258 , n10259 );
or ( n10261 , n10257 , n10260 );
buf ( n10262 , n4610 );
buf ( n10263 , n5634 );
xor ( n10264 , n10262 , n10263 );
or ( n10265 , n10261 , n10264 );
buf ( n10266 , n4611 );
buf ( n10267 , n5635 );
xor ( n10268 , n10266 , n10267 );
or ( n10269 , n10265 , n10268 );
buf ( n10270 , n4612 );
buf ( n10271 , n5636 );
xor ( n10272 , n10270 , n10271 );
or ( n10273 , n10269 , n10272 );
buf ( n10274 , n4613 );
buf ( n10275 , n5637 );
xor ( n10276 , n10274 , n10275 );
or ( n10277 , n10273 , n10276 );
buf ( n10278 , n4614 );
buf ( n10279 , n5638 );
xor ( n10280 , n10278 , n10279 );
or ( n10281 , n10277 , n10280 );
buf ( n10282 , n4615 );
buf ( n10283 , n5639 );
xor ( n10284 , n10282 , n10283 );
or ( n10285 , n10281 , n10284 );
buf ( n10286 , n4616 );
buf ( n10287 , n5640 );
xor ( n10288 , n10286 , n10287 );
or ( n10289 , n10285 , n10288 );
buf ( n10290 , n4617 );
buf ( n10291 , n5641 );
xor ( n10292 , n10290 , n10291 );
or ( n10293 , n10289 , n10292 );
buf ( n10294 , n4618 );
buf ( n10295 , n5642 );
xor ( n10296 , n10294 , n10295 );
or ( n10297 , n10293 , n10296 );
buf ( n10298 , n4619 );
buf ( n10299 , n5643 );
xor ( n10300 , n10298 , n10299 );
or ( n10301 , n10297 , n10300 );
buf ( n10302 , n4620 );
buf ( n10303 , n5644 );
xor ( n10304 , n10302 , n10303 );
or ( n10305 , n10301 , n10304 );
buf ( n10306 , n4621 );
buf ( n10307 , n5645 );
xor ( n10308 , n10306 , n10307 );
or ( n10309 , n10305 , n10308 );
buf ( n10310 , n4622 );
buf ( n10311 , n5646 );
xor ( n10312 , n10310 , n10311 );
or ( n10313 , n10309 , n10312 );
buf ( n10314 , n4623 );
buf ( n10315 , n5647 );
xor ( n10316 , n10314 , n10315 );
or ( n10317 , n10313 , n10316 );
buf ( n10318 , n4624 );
buf ( n10319 , n5648 );
xor ( n10320 , n10318 , n10319 );
or ( n10321 , n10317 , n10320 );
buf ( n10322 , n4625 );
buf ( n10323 , n5649 );
xor ( n10324 , n10322 , n10323 );
or ( n10325 , n10321 , n10324 );
buf ( n10326 , n4626 );
buf ( n10327 , n5650 );
xor ( n10328 , n10326 , n10327 );
or ( n10329 , n10325 , n10328 );
buf ( n10330 , n4627 );
buf ( n10331 , n5651 );
xor ( n10332 , n10330 , n10331 );
or ( n10333 , n10329 , n10332 );
buf ( n10334 , n4628 );
buf ( n10335 , n5652 );
xor ( n10336 , n10334 , n10335 );
or ( n10337 , n10333 , n10336 );
buf ( n10338 , n4629 );
buf ( n10339 , n5653 );
xor ( n10340 , n10338 , n10339 );
or ( n10341 , n10337 , n10340 );
buf ( n10342 , n4630 );
buf ( n10343 , n5654 );
xor ( n10344 , n10342 , n10343 );
or ( n10345 , n10341 , n10344 );
buf ( n10346 , n4631 );
buf ( n10347 , n5655 );
xor ( n10348 , n10346 , n10347 );
or ( n10349 , n10345 , n10348 );
buf ( n10350 , n4632 );
buf ( n10351 , n5656 );
xor ( n10352 , n10350 , n10351 );
or ( n10353 , n10349 , n10352 );
buf ( n10354 , n4633 );
buf ( n10355 , n5657 );
xor ( n10356 , n10354 , n10355 );
or ( n10357 , n10353 , n10356 );
buf ( n10358 , n4634 );
buf ( n10359 , n5658 );
xor ( n10360 , n10358 , n10359 );
or ( n10361 , n10357 , n10360 );
buf ( n10362 , n4635 );
buf ( n10363 , n5659 );
xor ( n10364 , n10362 , n10363 );
or ( n10365 , n10361 , n10364 );
buf ( n10366 , n4636 );
buf ( n10367 , n5660 );
xor ( n10368 , n10366 , n10367 );
or ( n10369 , n10365 , n10368 );
buf ( n10370 , n4637 );
buf ( n10371 , n5661 );
xor ( n10372 , n10370 , n10371 );
or ( n10373 , n10369 , n10372 );
buf ( n10374 , n4638 );
buf ( n10375 , n5662 );
xor ( n10376 , n10374 , n10375 );
or ( n10377 , n10373 , n10376 );
buf ( n10378 , n4639 );
buf ( n10379 , n5663 );
xor ( n10380 , n10378 , n10379 );
or ( n10381 , n10377 , n10380 );
buf ( n10382 , n4640 );
buf ( n10383 , n5664 );
xor ( n10384 , n10382 , n10383 );
or ( n10385 , n10381 , n10384 );
buf ( n10386 , n4641 );
buf ( n10387 , n5665 );
xor ( n10388 , n10386 , n10387 );
or ( n10389 , n10385 , n10388 );
buf ( n10390 , n4642 );
buf ( n10391 , n5666 );
xor ( n10392 , n10390 , n10391 );
or ( n10393 , n10389 , n10392 );
buf ( n10394 , n4643 );
buf ( n10395 , n5667 );
xor ( n10396 , n10394 , n10395 );
or ( n10397 , n10393 , n10396 );
buf ( n10398 , n4644 );
buf ( n10399 , n5668 );
xor ( n10400 , n10398 , n10399 );
or ( n10401 , n10397 , n10400 );
buf ( n10402 , n4645 );
buf ( n10403 , n5669 );
xor ( n10404 , n10402 , n10403 );
or ( n10405 , n10401 , n10404 );
buf ( n10406 , n4646 );
buf ( n10407 , n5670 );
xor ( n10408 , n10406 , n10407 );
or ( n10409 , n10405 , n10408 );
buf ( n10410 , n4647 );
buf ( n10411 , n5671 );
xor ( n10412 , n10410 , n10411 );
or ( n10413 , n10409 , n10412 );
buf ( n10414 , n4648 );
buf ( n10415 , n5672 );
xor ( n10416 , n10414 , n10415 );
or ( n10417 , n10413 , n10416 );
buf ( n10418 , n4649 );
buf ( n10419 , n5673 );
xor ( n10420 , n10418 , n10419 );
or ( n10421 , n10417 , n10420 );
buf ( n10422 , n4650 );
buf ( n10423 , n5674 );
xor ( n10424 , n10422 , n10423 );
or ( n10425 , n10421 , n10424 );
buf ( n10426 , n4651 );
buf ( n10427 , n5675 );
xor ( n10428 , n10426 , n10427 );
or ( n10429 , n10425 , n10428 );
buf ( n10430 , n4652 );
buf ( n10431 , n5676 );
xor ( n10432 , n10430 , n10431 );
or ( n10433 , n10429 , n10432 );
buf ( n10434 , n4653 );
buf ( n10435 , n5677 );
xor ( n10436 , n10434 , n10435 );
or ( n10437 , n10433 , n10436 );
buf ( n10438 , n4654 );
buf ( n10439 , n5678 );
xor ( n10440 , n10438 , n10439 );
or ( n10441 , n10437 , n10440 );
buf ( n10442 , n4655 );
buf ( n10443 , n5679 );
xor ( n10444 , n10442 , n10443 );
or ( n10445 , n10441 , n10444 );
buf ( n10446 , n4656 );
buf ( n10447 , n5680 );
xor ( n10448 , n10446 , n10447 );
or ( n10449 , n10445 , n10448 );
buf ( n10450 , n4657 );
buf ( n10451 , n5681 );
xor ( n10452 , n10450 , n10451 );
or ( n10453 , n10449 , n10452 );
buf ( n10454 , n4658 );
buf ( n10455 , n5682 );
xor ( n10456 , n10454 , n10455 );
or ( n10457 , n10453 , n10456 );
buf ( n10458 , n4659 );
buf ( n10459 , n5683 );
xor ( n10460 , n10458 , n10459 );
or ( n10461 , n10457 , n10460 );
buf ( n10462 , n4660 );
buf ( n10463 , n5684 );
xor ( n10464 , n10462 , n10463 );
or ( n10465 , n10461 , n10464 );
buf ( n10466 , n4661 );
buf ( n10467 , n5685 );
xor ( n10468 , n10466 , n10467 );
or ( n10469 , n10465 , n10468 );
buf ( n10470 , n4662 );
buf ( n10471 , n5686 );
xor ( n10472 , n10470 , n10471 );
or ( n10473 , n10469 , n10472 );
buf ( n10474 , n4663 );
buf ( n10475 , n5687 );
xor ( n10476 , n10474 , n10475 );
or ( n10477 , n10473 , n10476 );
buf ( n10478 , n4664 );
buf ( n10479 , n5688 );
xor ( n10480 , n10478 , n10479 );
or ( n10481 , n10477 , n10480 );
buf ( n10482 , n4665 );
buf ( n10483 , n5689 );
xor ( n10484 , n10482 , n10483 );
or ( n10485 , n10481 , n10484 );
buf ( n10486 , n4666 );
buf ( n10487 , n5690 );
xor ( n10488 , n10486 , n10487 );
or ( n10489 , n10485 , n10488 );
buf ( n10490 , n4667 );
buf ( n10491 , n5691 );
xor ( n10492 , n10490 , n10491 );
or ( n10493 , n10489 , n10492 );
buf ( n10494 , n4668 );
buf ( n10495 , n5692 );
xor ( n10496 , n10494 , n10495 );
or ( n10497 , n10493 , n10496 );
buf ( n10498 , n4669 );
buf ( n10499 , n5693 );
xor ( n10500 , n10498 , n10499 );
or ( n10501 , n10497 , n10500 );
buf ( n10502 , n4670 );
buf ( n10503 , n5694 );
xor ( n10504 , n10502 , n10503 );
or ( n10505 , n10501 , n10504 );
buf ( n10506 , n4671 );
buf ( n10507 , n5695 );
xor ( n10508 , n10506 , n10507 );
or ( n10509 , n10505 , n10508 );
buf ( n10510 , n4672 );
buf ( n10511 , n5696 );
xor ( n10512 , n10510 , n10511 );
or ( n10513 , n10509 , n10512 );
buf ( n10514 , n4673 );
buf ( n10515 , n5697 );
xor ( n10516 , n10514 , n10515 );
or ( n10517 , n10513 , n10516 );
buf ( n10518 , n4674 );
buf ( n10519 , n5698 );
xor ( n10520 , n10518 , n10519 );
or ( n10521 , n10517 , n10520 );
buf ( n10522 , n4675 );
buf ( n10523 , n5699 );
xor ( n10524 , n10522 , n10523 );
or ( n10525 , n10521 , n10524 );
buf ( n10526 , n4676 );
buf ( n10527 , n5700 );
xor ( n10528 , n10526 , n10527 );
or ( n10529 , n10525 , n10528 );
buf ( n10530 , n4677 );
buf ( n10531 , n5701 );
xor ( n10532 , n10530 , n10531 );
or ( n10533 , n10529 , n10532 );
buf ( n10534 , n4678 );
buf ( n10535 , n5702 );
xor ( n10536 , n10534 , n10535 );
or ( n10537 , n10533 , n10536 );
buf ( n10538 , n4679 );
buf ( n10539 , n5703 );
xor ( n10540 , n10538 , n10539 );
or ( n10541 , n10537 , n10540 );
buf ( n10542 , n4680 );
buf ( n10543 , n5704 );
xor ( n10544 , n10542 , n10543 );
or ( n10545 , n10541 , n10544 );
buf ( n10546 , n4681 );
buf ( n10547 , n5705 );
xor ( n10548 , n10546 , n10547 );
or ( n10549 , n10545 , n10548 );
buf ( n10550 , n4682 );
buf ( n10551 , n5706 );
xor ( n10552 , n10550 , n10551 );
or ( n10553 , n10549 , n10552 );
buf ( n10554 , n4683 );
buf ( n10555 , n5707 );
xor ( n10556 , n10554 , n10555 );
or ( n10557 , n10553 , n10556 );
buf ( n10558 , n4684 );
buf ( n10559 , n5708 );
xor ( n10560 , n10558 , n10559 );
or ( n10561 , n10557 , n10560 );
buf ( n10562 , n4685 );
buf ( n10563 , n5709 );
xor ( n10564 , n10562 , n10563 );
or ( n10565 , n10561 , n10564 );
buf ( n10566 , n4686 );
buf ( n10567 , n5710 );
xor ( n10568 , n10566 , n10567 );
or ( n10569 , n10565 , n10568 );
buf ( n10570 , n4687 );
buf ( n10571 , n5711 );
xor ( n10572 , n10570 , n10571 );
or ( n10573 , n10569 , n10572 );
buf ( n10574 , n4688 );
buf ( n10575 , n5712 );
xor ( n10576 , n10574 , n10575 );
or ( n10577 , n10573 , n10576 );
buf ( n10578 , n4689 );
buf ( n10579 , n5713 );
xor ( n10580 , n10578 , n10579 );
or ( n10581 , n10577 , n10580 );
buf ( n10582 , n4690 );
buf ( n10583 , n5714 );
xor ( n10584 , n10582 , n10583 );
or ( n10585 , n10581 , n10584 );
buf ( n10586 , n4691 );
buf ( n10587 , n5715 );
xor ( n10588 , n10586 , n10587 );
or ( n10589 , n10585 , n10588 );
buf ( n10590 , n4692 );
buf ( n10591 , n5716 );
xor ( n10592 , n10590 , n10591 );
or ( n10593 , n10589 , n10592 );
buf ( n10594 , n4693 );
buf ( n10595 , n5717 );
xor ( n10596 , n10594 , n10595 );
or ( n10597 , n10593 , n10596 );
buf ( n10598 , n4694 );
buf ( n10599 , n5718 );
xor ( n10600 , n10598 , n10599 );
or ( n10601 , n10597 , n10600 );
buf ( n10602 , n4695 );
buf ( n10603 , n5719 );
xor ( n10604 , n10602 , n10603 );
or ( n10605 , n10601 , n10604 );
buf ( n10606 , n4696 );
buf ( n10607 , n5720 );
xor ( n10608 , n10606 , n10607 );
or ( n10609 , n10605 , n10608 );
buf ( n10610 , n4697 );
buf ( n10611 , n5721 );
xor ( n10612 , n10610 , n10611 );
or ( n10613 , n10609 , n10612 );
buf ( n10614 , n4698 );
buf ( n10615 , n5722 );
xor ( n10616 , n10614 , n10615 );
or ( n10617 , n10613 , n10616 );
buf ( n10618 , n4699 );
buf ( n10619 , n5723 );
xor ( n10620 , n10618 , n10619 );
or ( n10621 , n10617 , n10620 );
buf ( n10622 , n4700 );
buf ( n10623 , n5724 );
xor ( n10624 , n10622 , n10623 );
or ( n10625 , n10621 , n10624 );
buf ( n10626 , n4701 );
buf ( n10627 , n5725 );
xor ( n10628 , n10626 , n10627 );
or ( n10629 , n10625 , n10628 );
buf ( n10630 , n4702 );
buf ( n10631 , n5726 );
xor ( n10632 , n10630 , n10631 );
or ( n10633 , n10629 , n10632 );
buf ( n10634 , n4703 );
buf ( n10635 , n5727 );
xor ( n10636 , n10634 , n10635 );
or ( n10637 , n10633 , n10636 );
buf ( n10638 , n4704 );
buf ( n10639 , n5728 );
xor ( n10640 , n10638 , n10639 );
or ( n10641 , n10637 , n10640 );
buf ( n10642 , n4705 );
buf ( n10643 , n5729 );
xor ( n10644 , n10642 , n10643 );
or ( n10645 , n10641 , n10644 );
buf ( n10646 , n4706 );
buf ( n10647 , n5730 );
xor ( n10648 , n10646 , n10647 );
or ( n10649 , n10645 , n10648 );
buf ( n10650 , n4707 );
buf ( n10651 , n5731 );
xor ( n10652 , n10650 , n10651 );
or ( n10653 , n10649 , n10652 );
buf ( n10654 , n4708 );
buf ( n10655 , n5732 );
xor ( n10656 , n10654 , n10655 );
or ( n10657 , n10653 , n10656 );
buf ( n10658 , n4709 );
buf ( n10659 , n5733 );
xor ( n10660 , n10658 , n10659 );
or ( n10661 , n10657 , n10660 );
buf ( n10662 , n4710 );
buf ( n10663 , n5734 );
xor ( n10664 , n10662 , n10663 );
or ( n10665 , n10661 , n10664 );
buf ( n10666 , n4711 );
buf ( n10667 , n5735 );
xor ( n10668 , n10666 , n10667 );
or ( n10669 , n10665 , n10668 );
buf ( n10670 , n4712 );
buf ( n10671 , n5736 );
xor ( n10672 , n10670 , n10671 );
or ( n10673 , n10669 , n10672 );
buf ( n10674 , n4713 );
buf ( n10675 , n5737 );
xor ( n10676 , n10674 , n10675 );
or ( n10677 , n10673 , n10676 );
buf ( n10678 , n4714 );
buf ( n10679 , n5738 );
xor ( n10680 , n10678 , n10679 );
or ( n10681 , n10677 , n10680 );
buf ( n10682 , n4715 );
buf ( n10683 , n5739 );
xor ( n10684 , n10682 , n10683 );
or ( n10685 , n10681 , n10684 );
buf ( n10686 , n4716 );
buf ( n10687 , n5740 );
xor ( n10688 , n10686 , n10687 );
or ( n10689 , n10685 , n10688 );
buf ( n10690 , n4717 );
buf ( n10691 , n5741 );
xor ( n10692 , n10690 , n10691 );
or ( n10693 , n10689 , n10692 );
buf ( n10694 , n4718 );
buf ( n10695 , n5742 );
xor ( n10696 , n10694 , n10695 );
or ( n10697 , n10693 , n10696 );
buf ( n10698 , n4719 );
buf ( n10699 , n5743 );
xor ( n10700 , n10698 , n10699 );
or ( n10701 , n10697 , n10700 );
buf ( n10702 , n4720 );
buf ( n10703 , n5744 );
xor ( n10704 , n10702 , n10703 );
or ( n10705 , n10701 , n10704 );
buf ( n10706 , n4721 );
buf ( n10707 , n5745 );
xor ( n10708 , n10706 , n10707 );
or ( n10709 , n10705 , n10708 );
buf ( n10710 , n4722 );
buf ( n10711 , n5746 );
xor ( n10712 , n10710 , n10711 );
or ( n10713 , n10709 , n10712 );
buf ( n10714 , n4723 );
buf ( n10715 , n5747 );
xor ( n10716 , n10714 , n10715 );
or ( n10717 , n10713 , n10716 );
buf ( n10718 , n4724 );
buf ( n10719 , n5748 );
xor ( n10720 , n10718 , n10719 );
or ( n10721 , n10717 , n10720 );
buf ( n10722 , n4725 );
buf ( n10723 , n5749 );
xor ( n10724 , n10722 , n10723 );
or ( n10725 , n10721 , n10724 );
buf ( n10726 , n4726 );
buf ( n10727 , n5750 );
xor ( n10728 , n10726 , n10727 );
or ( n10729 , n10725 , n10728 );
buf ( n10730 , n4727 );
buf ( n10731 , n5751 );
xor ( n10732 , n10730 , n10731 );
or ( n10733 , n10729 , n10732 );
buf ( n10734 , n4728 );
buf ( n10735 , n5752 );
xor ( n10736 , n10734 , n10735 );
or ( n10737 , n10733 , n10736 );
buf ( n10738 , n4729 );
buf ( n10739 , n5753 );
xor ( n10740 , n10738 , n10739 );
or ( n10741 , n10737 , n10740 );
buf ( n10742 , n4730 );
buf ( n10743 , n5754 );
xor ( n10744 , n10742 , n10743 );
or ( n10745 , n10741 , n10744 );
buf ( n10746 , n4731 );
buf ( n10747 , n5755 );
xor ( n10748 , n10746 , n10747 );
or ( n10749 , n10745 , n10748 );
buf ( n10750 , n4732 );
buf ( n10751 , n5756 );
xor ( n10752 , n10750 , n10751 );
or ( n10753 , n10749 , n10752 );
buf ( n10754 , n4733 );
buf ( n10755 , n5757 );
xor ( n10756 , n10754 , n10755 );
or ( n10757 , n10753 , n10756 );
buf ( n10758 , n4734 );
buf ( n10759 , n5758 );
xor ( n10760 , n10758 , n10759 );
or ( n10761 , n10757 , n10760 );
buf ( n10762 , n4735 );
buf ( n10763 , n5759 );
xor ( n10764 , n10762 , n10763 );
or ( n10765 , n10761 , n10764 );
buf ( n10766 , n4736 );
buf ( n10767 , n5760 );
xor ( n10768 , n10766 , n10767 );
or ( n10769 , n10765 , n10768 );
buf ( n10770 , n4737 );
buf ( n10771 , n5761 );
xor ( n10772 , n10770 , n10771 );
or ( n10773 , n10769 , n10772 );
buf ( n10774 , n4738 );
buf ( n10775 , n5762 );
xor ( n10776 , n10774 , n10775 );
or ( n10777 , n10773 , n10776 );
buf ( n10778 , n4739 );
buf ( n10779 , n5763 );
xor ( n10780 , n10778 , n10779 );
or ( n10781 , n10777 , n10780 );
buf ( n10782 , n4740 );
buf ( n10783 , n5764 );
xor ( n10784 , n10782 , n10783 );
or ( n10785 , n10781 , n10784 );
buf ( n10786 , n4741 );
buf ( n10787 , n5765 );
xor ( n10788 , n10786 , n10787 );
or ( n10789 , n10785 , n10788 );
buf ( n10790 , n4742 );
buf ( n10791 , n5766 );
xor ( n10792 , n10790 , n10791 );
or ( n10793 , n10789 , n10792 );
buf ( n10794 , n4743 );
buf ( n10795 , n5767 );
xor ( n10796 , n10794 , n10795 );
or ( n10797 , n10793 , n10796 );
buf ( n10798 , n4744 );
buf ( n10799 , n5768 );
xor ( n10800 , n10798 , n10799 );
or ( n10801 , n10797 , n10800 );
buf ( n10802 , n4745 );
buf ( n10803 , n5769 );
xor ( n10804 , n10802 , n10803 );
or ( n10805 , n10801 , n10804 );
buf ( n10806 , n4746 );
buf ( n10807 , n5770 );
xor ( n10808 , n10806 , n10807 );
or ( n10809 , n10805 , n10808 );
buf ( n10810 , n4747 );
buf ( n10811 , n5771 );
xor ( n10812 , n10810 , n10811 );
or ( n10813 , n10809 , n10812 );
buf ( n10814 , n4748 );
buf ( n10815 , n5772 );
xor ( n10816 , n10814 , n10815 );
or ( n10817 , n10813 , n10816 );
buf ( n10818 , n4749 );
buf ( n10819 , n5773 );
xor ( n10820 , n10818 , n10819 );
or ( n10821 , n10817 , n10820 );
buf ( n10822 , n4750 );
buf ( n10823 , n5774 );
xor ( n10824 , n10822 , n10823 );
or ( n10825 , n10821 , n10824 );
buf ( n10826 , n4751 );
buf ( n10827 , n5775 );
xor ( n10828 , n10826 , n10827 );
or ( n10829 , n10825 , n10828 );
buf ( n10830 , n4752 );
buf ( n10831 , n5776 );
xor ( n10832 , n10830 , n10831 );
or ( n10833 , n10829 , n10832 );
buf ( n10834 , n4753 );
buf ( n10835 , n5777 );
xor ( n10836 , n10834 , n10835 );
or ( n10837 , n10833 , n10836 );
buf ( n10838 , n4754 );
buf ( n10839 , n5778 );
xor ( n10840 , n10838 , n10839 );
or ( n10841 , n10837 , n10840 );
buf ( n10842 , n4755 );
buf ( n10843 , n5779 );
xor ( n10844 , n10842 , n10843 );
or ( n10845 , n10841 , n10844 );
buf ( n10846 , n4756 );
buf ( n10847 , n5780 );
xor ( n10848 , n10846 , n10847 );
or ( n10849 , n10845 , n10848 );
buf ( n10850 , n4757 );
buf ( n10851 , n5781 );
xor ( n10852 , n10850 , n10851 );
or ( n10853 , n10849 , n10852 );
buf ( n10854 , n4758 );
buf ( n10855 , n5782 );
xor ( n10856 , n10854 , n10855 );
or ( n10857 , n10853 , n10856 );
buf ( n10858 , n4759 );
buf ( n10859 , n5783 );
xor ( n10860 , n10858 , n10859 );
or ( n10861 , n10857 , n10860 );
buf ( n10862 , n4760 );
buf ( n10863 , n5784 );
xor ( n10864 , n10862 , n10863 );
or ( n10865 , n10861 , n10864 );
buf ( n10866 , n4761 );
buf ( n10867 , n5785 );
xor ( n10868 , n10866 , n10867 );
or ( n10869 , n10865 , n10868 );
buf ( n10870 , n4762 );
buf ( n10871 , n5786 );
xor ( n10872 , n10870 , n10871 );
or ( n10873 , n10869 , n10872 );
buf ( n10874 , n4763 );
buf ( n10875 , n5787 );
xor ( n10876 , n10874 , n10875 );
or ( n10877 , n10873 , n10876 );
buf ( n10878 , n4764 );
buf ( n10879 , n5788 );
xor ( n10880 , n10878 , n10879 );
or ( n10881 , n10877 , n10880 );
buf ( n10882 , n4765 );
buf ( n10883 , n5789 );
xor ( n10884 , n10882 , n10883 );
or ( n10885 , n10881 , n10884 );
buf ( n10886 , n4766 );
buf ( n10887 , n5790 );
xor ( n10888 , n10886 , n10887 );
or ( n10889 , n10885 , n10888 );
buf ( n10890 , n4767 );
buf ( n10891 , n5791 );
xor ( n10892 , n10890 , n10891 );
or ( n10893 , n10889 , n10892 );
buf ( n10894 , n4768 );
buf ( n10895 , n5792 );
xor ( n10896 , n10894 , n10895 );
or ( n10897 , n10893 , n10896 );
buf ( n10898 , n4769 );
buf ( n10899 , n5793 );
xor ( n10900 , n10898 , n10899 );
or ( n10901 , n10897 , n10900 );
buf ( n10902 , n4770 );
buf ( n10903 , n5794 );
xor ( n10904 , n10902 , n10903 );
or ( n10905 , n10901 , n10904 );
buf ( n10906 , n4771 );
buf ( n10907 , n5795 );
xor ( n10908 , n10906 , n10907 );
or ( n10909 , n10905 , n10908 );
buf ( n10910 , n4772 );
buf ( n10911 , n5796 );
xor ( n10912 , n10910 , n10911 );
or ( n10913 , n10909 , n10912 );
buf ( n10914 , n4773 );
buf ( n10915 , n5797 );
xor ( n10916 , n10914 , n10915 );
or ( n10917 , n10913 , n10916 );
buf ( n10918 , n4774 );
buf ( n10919 , n5798 );
xor ( n10920 , n10918 , n10919 );
or ( n10921 , n10917 , n10920 );
buf ( n10922 , n4775 );
buf ( n10923 , n5799 );
xor ( n10924 , n10922 , n10923 );
or ( n10925 , n10921 , n10924 );
buf ( n10926 , n4776 );
buf ( n10927 , n5800 );
xor ( n10928 , n10926 , n10927 );
or ( n10929 , n10925 , n10928 );
buf ( n10930 , n4777 );
buf ( n10931 , n5801 );
xor ( n10932 , n10930 , n10931 );
or ( n10933 , n10929 , n10932 );
buf ( n10934 , n4778 );
buf ( n10935 , n5802 );
xor ( n10936 , n10934 , n10935 );
or ( n10937 , n10933 , n10936 );
buf ( n10938 , n4779 );
buf ( n10939 , n5803 );
xor ( n10940 , n10938 , n10939 );
or ( n10941 , n10937 , n10940 );
buf ( n10942 , n4780 );
buf ( n10943 , n5804 );
xor ( n10944 , n10942 , n10943 );
or ( n10945 , n10941 , n10944 );
buf ( n10946 , n4781 );
buf ( n10947 , n5805 );
xor ( n10948 , n10946 , n10947 );
or ( n10949 , n10945 , n10948 );
buf ( n10950 , n4782 );
buf ( n10951 , n5806 );
xor ( n10952 , n10950 , n10951 );
or ( n10953 , n10949 , n10952 );
buf ( n10954 , n4783 );
buf ( n10955 , n5807 );
xor ( n10956 , n10954 , n10955 );
or ( n10957 , n10953 , n10956 );
buf ( n10958 , n4784 );
buf ( n10959 , n5808 );
xor ( n10960 , n10958 , n10959 );
or ( n10961 , n10957 , n10960 );
buf ( n10962 , n4785 );
buf ( n10963 , n5809 );
xor ( n10964 , n10962 , n10963 );
or ( n10965 , n10961 , n10964 );
buf ( n10966 , n4786 );
buf ( n10967 , n5810 );
xor ( n10968 , n10966 , n10967 );
or ( n10969 , n10965 , n10968 );
buf ( n10970 , n4787 );
buf ( n10971 , n5811 );
xor ( n10972 , n10970 , n10971 );
or ( n10973 , n10969 , n10972 );
buf ( n10974 , n4788 );
buf ( n10975 , n5812 );
xor ( n10976 , n10974 , n10975 );
or ( n10977 , n10973 , n10976 );
buf ( n10978 , n4789 );
buf ( n10979 , n5813 );
xor ( n10980 , n10978 , n10979 );
or ( n10981 , n10977 , n10980 );
buf ( n10982 , n4790 );
buf ( n10983 , n5814 );
xor ( n10984 , n10982 , n10983 );
or ( n10985 , n10981 , n10984 );
buf ( n10986 , n4791 );
buf ( n10987 , n5815 );
xor ( n10988 , n10986 , n10987 );
or ( n10989 , n10985 , n10988 );
buf ( n10990 , n4792 );
buf ( n10991 , n5816 );
xor ( n10992 , n10990 , n10991 );
or ( n10993 , n10989 , n10992 );
buf ( n10994 , n4793 );
buf ( n10995 , n5817 );
xor ( n10996 , n10994 , n10995 );
or ( n10997 , n10993 , n10996 );
buf ( n10998 , n4794 );
buf ( n10999 , n5818 );
xor ( n11000 , n10998 , n10999 );
or ( n11001 , n10997 , n11000 );
buf ( n11002 , n4795 );
buf ( n11003 , n5819 );
xor ( n11004 , n11002 , n11003 );
or ( n11005 , n11001 , n11004 );
buf ( n11006 , n4796 );
buf ( n11007 , n5820 );
xor ( n11008 , n11006 , n11007 );
or ( n11009 , n11005 , n11008 );
buf ( n11010 , n4797 );
buf ( n11011 , n5821 );
xor ( n11012 , n11010 , n11011 );
or ( n11013 , n11009 , n11012 );
buf ( n11014 , n4798 );
buf ( n11015 , n5822 );
xor ( n11016 , n11014 , n11015 );
or ( n11017 , n11013 , n11016 );
buf ( n11018 , n4799 );
buf ( n11019 , n5823 );
xor ( n11020 , n11018 , n11019 );
or ( n11021 , n11017 , n11020 );
buf ( n11022 , n4800 );
buf ( n11023 , n5824 );
xor ( n11024 , n11022 , n11023 );
or ( n11025 , n11021 , n11024 );
buf ( n11026 , n4801 );
buf ( n11027 , n5825 );
xor ( n11028 , n11026 , n11027 );
or ( n11029 , n11025 , n11028 );
buf ( n11030 , n4802 );
buf ( n11031 , n5826 );
xor ( n11032 , n11030 , n11031 );
or ( n11033 , n11029 , n11032 );
buf ( n11034 , n4803 );
buf ( n11035 , n5827 );
xor ( n11036 , n11034 , n11035 );
or ( n11037 , n11033 , n11036 );
buf ( n11038 , n4804 );
buf ( n11039 , n5828 );
xor ( n11040 , n11038 , n11039 );
or ( n11041 , n11037 , n11040 );
buf ( n11042 , n4805 );
buf ( n11043 , n5829 );
xor ( n11044 , n11042 , n11043 );
or ( n11045 , n11041 , n11044 );
buf ( n11046 , n4806 );
buf ( n11047 , n5830 );
xor ( n11048 , n11046 , n11047 );
or ( n11049 , n11045 , n11048 );
buf ( n11050 , n4807 );
buf ( n11051 , n5831 );
xor ( n11052 , n11050 , n11051 );
or ( n11053 , n11049 , n11052 );
buf ( n11054 , n4808 );
buf ( n11055 , n5832 );
xor ( n11056 , n11054 , n11055 );
or ( n11057 , n11053 , n11056 );
buf ( n11058 , n4809 );
buf ( n11059 , n5833 );
xor ( n11060 , n11058 , n11059 );
or ( n11061 , n11057 , n11060 );
buf ( n11062 , n4810 );
buf ( n11063 , n5834 );
xor ( n11064 , n11062 , n11063 );
or ( n11065 , n11061 , n11064 );
buf ( n11066 , n4811 );
buf ( n11067 , n5835 );
xor ( n11068 , n11066 , n11067 );
or ( n11069 , n11065 , n11068 );
buf ( n11070 , n4812 );
buf ( n11071 , n5836 );
xor ( n11072 , n11070 , n11071 );
or ( n11073 , n11069 , n11072 );
buf ( n11074 , n4813 );
buf ( n11075 , n5837 );
xor ( n11076 , n11074 , n11075 );
or ( n11077 , n11073 , n11076 );
buf ( n11078 , n4814 );
buf ( n11079 , n5838 );
xor ( n11080 , n11078 , n11079 );
or ( n11081 , n11077 , n11080 );
buf ( n11082 , n4815 );
buf ( n11083 , n5839 );
xor ( n11084 , n11082 , n11083 );
or ( n11085 , n11081 , n11084 );
buf ( n11086 , n4816 );
buf ( n11087 , n5840 );
xor ( n11088 , n11086 , n11087 );
or ( n11089 , n11085 , n11088 );
buf ( n11090 , n4817 );
buf ( n11091 , n5841 );
xor ( n11092 , n11090 , n11091 );
or ( n11093 , n11089 , n11092 );
buf ( n11094 , n4818 );
buf ( n11095 , n5842 );
xor ( n11096 , n11094 , n11095 );
or ( n11097 , n11093 , n11096 );
buf ( n11098 , n4819 );
buf ( n11099 , n5843 );
xor ( n11100 , n11098 , n11099 );
or ( n11101 , n11097 , n11100 );
buf ( n11102 , n4820 );
buf ( n11103 , n5844 );
xor ( n11104 , n11102 , n11103 );
or ( n11105 , n11101 , n11104 );
buf ( n11106 , n4821 );
buf ( n11107 , n5845 );
xor ( n11108 , n11106 , n11107 );
or ( n11109 , n11105 , n11108 );
buf ( n11110 , n4822 );
buf ( n11111 , n5846 );
xor ( n11112 , n11110 , n11111 );
or ( n11113 , n11109 , n11112 );
buf ( n11114 , n4823 );
buf ( n11115 , n5847 );
xor ( n11116 , n11114 , n11115 );
or ( n11117 , n11113 , n11116 );
buf ( n11118 , n4824 );
buf ( n11119 , n5848 );
xor ( n11120 , n11118 , n11119 );
or ( n11121 , n11117 , n11120 );
buf ( n11122 , n4825 );
buf ( n11123 , n5849 );
xor ( n11124 , n11122 , n11123 );
or ( n11125 , n11121 , n11124 );
buf ( n11126 , n4826 );
buf ( n11127 , n5850 );
xor ( n11128 , n11126 , n11127 );
or ( n11129 , n11125 , n11128 );
buf ( n11130 , n4827 );
buf ( n11131 , n5851 );
xor ( n11132 , n11130 , n11131 );
or ( n11133 , n11129 , n11132 );
buf ( n11134 , n4828 );
buf ( n11135 , n5852 );
xor ( n11136 , n11134 , n11135 );
or ( n11137 , n11133 , n11136 );
buf ( n11138 , n4829 );
buf ( n11139 , n5853 );
xor ( n11140 , n11138 , n11139 );
or ( n11141 , n11137 , n11140 );
buf ( n11142 , n4830 );
buf ( n11143 , n5854 );
xor ( n11144 , n11142 , n11143 );
or ( n11145 , n11141 , n11144 );
buf ( n11146 , n4831 );
buf ( n11147 , n5855 );
xor ( n11148 , n11146 , n11147 );
or ( n11149 , n11145 , n11148 );
buf ( n11150 , n4832 );
buf ( n11151 , n5856 );
xor ( n11152 , n11150 , n11151 );
or ( n11153 , n11149 , n11152 );
buf ( n11154 , n4833 );
buf ( n11155 , n5857 );
xor ( n11156 , n11154 , n11155 );
or ( n11157 , n11153 , n11156 );
buf ( n11158 , n4834 );
buf ( n11159 , n5858 );
xor ( n11160 , n11158 , n11159 );
or ( n11161 , n11157 , n11160 );
buf ( n11162 , n4835 );
buf ( n11163 , n5859 );
xor ( n11164 , n11162 , n11163 );
or ( n11165 , n11161 , n11164 );
buf ( n11166 , n4836 );
buf ( n11167 , n5860 );
xor ( n11168 , n11166 , n11167 );
or ( n11169 , n11165 , n11168 );
buf ( n11170 , n4837 );
buf ( n11171 , n5861 );
xor ( n11172 , n11170 , n11171 );
or ( n11173 , n11169 , n11172 );
buf ( n11174 , n4838 );
buf ( n11175 , n5862 );
xor ( n11176 , n11174 , n11175 );
or ( n11177 , n11173 , n11176 );
buf ( n11178 , n4839 );
buf ( n11179 , n5863 );
xor ( n11180 , n11178 , n11179 );
or ( n11181 , n11177 , n11180 );
buf ( n11182 , n4840 );
buf ( n11183 , n5864 );
xor ( n11184 , n11182 , n11183 );
or ( n11185 , n11181 , n11184 );
buf ( n11186 , n4841 );
buf ( n11187 , n5865 );
xor ( n11188 , n11186 , n11187 );
or ( n11189 , n11185 , n11188 );
buf ( n11190 , n4842 );
buf ( n11191 , n5866 );
xor ( n11192 , n11190 , n11191 );
or ( n11193 , n11189 , n11192 );
buf ( n11194 , n4843 );
buf ( n11195 , n5867 );
xor ( n11196 , n11194 , n11195 );
or ( n11197 , n11193 , n11196 );
buf ( n11198 , n4844 );
buf ( n11199 , n5868 );
xor ( n11200 , n11198 , n11199 );
or ( n11201 , n11197 , n11200 );
buf ( n11202 , n4845 );
buf ( n11203 , n5869 );
xor ( n11204 , n11202 , n11203 );
or ( n11205 , n11201 , n11204 );
buf ( n11206 , n4846 );
buf ( n11207 , n5870 );
xor ( n11208 , n11206 , n11207 );
or ( n11209 , n11205 , n11208 );
buf ( n11210 , n4847 );
buf ( n11211 , n5871 );
xor ( n11212 , n11210 , n11211 );
or ( n11213 , n11209 , n11212 );
buf ( n11214 , n4848 );
buf ( n11215 , n5872 );
xor ( n11216 , n11214 , n11215 );
or ( n11217 , n11213 , n11216 );
buf ( n11218 , n4849 );
buf ( n11219 , n5873 );
xor ( n11220 , n11218 , n11219 );
or ( n11221 , n11217 , n11220 );
buf ( n11222 , n4850 );
buf ( n11223 , n5874 );
xor ( n11224 , n11222 , n11223 );
or ( n11225 , n11221 , n11224 );
buf ( n11226 , n4851 );
buf ( n11227 , n5875 );
xor ( n11228 , n11226 , n11227 );
or ( n11229 , n11225 , n11228 );
buf ( n11230 , n4852 );
buf ( n11231 , n5876 );
xor ( n11232 , n11230 , n11231 );
or ( n11233 , n11229 , n11232 );
buf ( n11234 , n4853 );
buf ( n11235 , n5877 );
xor ( n11236 , n11234 , n11235 );
or ( n11237 , n11233 , n11236 );
buf ( n11238 , n4854 );
buf ( n11239 , n5878 );
xor ( n11240 , n11238 , n11239 );
or ( n11241 , n11237 , n11240 );
buf ( n11242 , n4855 );
buf ( n11243 , n5879 );
xor ( n11244 , n11242 , n11243 );
or ( n11245 , n11241 , n11244 );
buf ( n11246 , n4856 );
buf ( n11247 , n5880 );
xor ( n11248 , n11246 , n11247 );
or ( n11249 , n11245 , n11248 );
buf ( n11250 , n4857 );
buf ( n11251 , n5881 );
xor ( n11252 , n11250 , n11251 );
or ( n11253 , n11249 , n11252 );
buf ( n11254 , n4858 );
buf ( n11255 , n5882 );
xor ( n11256 , n11254 , n11255 );
or ( n11257 , n11253 , n11256 );
buf ( n11258 , n4859 );
buf ( n11259 , n5883 );
xor ( n11260 , n11258 , n11259 );
or ( n11261 , n11257 , n11260 );
buf ( n11262 , n4860 );
buf ( n11263 , n5884 );
xor ( n11264 , n11262 , n11263 );
or ( n11265 , n11261 , n11264 );
buf ( n11266 , n4861 );
buf ( n11267 , n5885 );
xor ( n11268 , n11266 , n11267 );
or ( n11269 , n11265 , n11268 );
buf ( n11270 , n4862 );
buf ( n11271 , n5886 );
xor ( n11272 , n11270 , n11271 );
or ( n11273 , n11269 , n11272 );
buf ( n11274 , n4863 );
buf ( n11275 , n5887 );
xor ( n11276 , n11274 , n11275 );
or ( n11277 , n11273 , n11276 );
buf ( n11278 , n4864 );
buf ( n11279 , n5888 );
xor ( n11280 , n11278 , n11279 );
or ( n11281 , n11277 , n11280 );
buf ( n11282 , n4865 );
buf ( n11283 , n5889 );
xor ( n11284 , n11282 , n11283 );
or ( n11285 , n11281 , n11284 );
buf ( n11286 , n4866 );
buf ( n11287 , n5890 );
xor ( n11288 , n11286 , n11287 );
or ( n11289 , n11285 , n11288 );
buf ( n11290 , n4867 );
buf ( n11291 , n5891 );
xor ( n11292 , n11290 , n11291 );
or ( n11293 , n11289 , n11292 );
buf ( n11294 , n4868 );
buf ( n11295 , n5892 );
xor ( n11296 , n11294 , n11295 );
or ( n11297 , n11293 , n11296 );
buf ( n11298 , n4869 );
buf ( n11299 , n5893 );
xor ( n11300 , n11298 , n11299 );
or ( n11301 , n11297 , n11300 );
buf ( n11302 , n4870 );
buf ( n11303 , n5894 );
xor ( n11304 , n11302 , n11303 );
or ( n11305 , n11301 , n11304 );
buf ( n11306 , n4871 );
buf ( n11307 , n5895 );
xor ( n11308 , n11306 , n11307 );
or ( n11309 , n11305 , n11308 );
buf ( n11310 , n4872 );
buf ( n11311 , n5896 );
xor ( n11312 , n11310 , n11311 );
or ( n11313 , n11309 , n11312 );
buf ( n11314 , n4873 );
buf ( n11315 , n5897 );
xor ( n11316 , n11314 , n11315 );
or ( n11317 , n11313 , n11316 );
buf ( n11318 , n4874 );
buf ( n11319 , n5898 );
xor ( n11320 , n11318 , n11319 );
or ( n11321 , n11317 , n11320 );
buf ( n11322 , n4875 );
buf ( n11323 , n5899 );
xor ( n11324 , n11322 , n11323 );
or ( n11325 , n11321 , n11324 );
buf ( n11326 , n4876 );
buf ( n11327 , n5900 );
xor ( n11328 , n11326 , n11327 );
or ( n11329 , n11325 , n11328 );
buf ( n11330 , n4877 );
buf ( n11331 , n5901 );
xor ( n11332 , n11330 , n11331 );
or ( n11333 , n11329 , n11332 );
buf ( n11334 , n4878 );
buf ( n11335 , n5902 );
xor ( n11336 , n11334 , n11335 );
or ( n11337 , n11333 , n11336 );
buf ( n11338 , n4879 );
buf ( n11339 , n5903 );
xor ( n11340 , n11338 , n11339 );
or ( n11341 , n11337 , n11340 );
buf ( n11342 , n4880 );
buf ( n11343 , n5904 );
xor ( n11344 , n11342 , n11343 );
or ( n11345 , n11341 , n11344 );
buf ( n11346 , n4881 );
buf ( n11347 , n5905 );
xor ( n11348 , n11346 , n11347 );
or ( n11349 , n11345 , n11348 );
buf ( n11350 , n4882 );
buf ( n11351 , n5906 );
xor ( n11352 , n11350 , n11351 );
or ( n11353 , n11349 , n11352 );
buf ( n11354 , n4883 );
buf ( n11355 , n5907 );
xor ( n11356 , n11354 , n11355 );
or ( n11357 , n11353 , n11356 );
buf ( n11358 , n4884 );
buf ( n11359 , n5908 );
xor ( n11360 , n11358 , n11359 );
or ( n11361 , n11357 , n11360 );
buf ( n11362 , n4885 );
buf ( n11363 , n5909 );
xor ( n11364 , n11362 , n11363 );
or ( n11365 , n11361 , n11364 );
buf ( n11366 , n4886 );
buf ( n11367 , n5910 );
xor ( n11368 , n11366 , n11367 );
or ( n11369 , n11365 , n11368 );
buf ( n11370 , n4887 );
buf ( n11371 , n5911 );
xor ( n11372 , n11370 , n11371 );
or ( n11373 , n11369 , n11372 );
buf ( n11374 , n4888 );
buf ( n11375 , n5912 );
xor ( n11376 , n11374 , n11375 );
or ( n11377 , n11373 , n11376 );
buf ( n11378 , n4889 );
buf ( n11379 , n5913 );
xor ( n11380 , n11378 , n11379 );
or ( n11381 , n11377 , n11380 );
buf ( n11382 , n4890 );
buf ( n11383 , n5914 );
xor ( n11384 , n11382 , n11383 );
or ( n11385 , n11381 , n11384 );
buf ( n11386 , n4891 );
buf ( n11387 , n5915 );
xor ( n11388 , n11386 , n11387 );
or ( n11389 , n11385 , n11388 );
buf ( n11390 , n4892 );
buf ( n11391 , n5916 );
xor ( n11392 , n11390 , n11391 );
or ( n11393 , n11389 , n11392 );
buf ( n11394 , n4893 );
buf ( n11395 , n5917 );
xor ( n11396 , n11394 , n11395 );
or ( n11397 , n11393 , n11396 );
buf ( n11398 , n4894 );
buf ( n11399 , n5918 );
xor ( n11400 , n11398 , n11399 );
or ( n11401 , n11397 , n11400 );
buf ( n11402 , n4895 );
buf ( n11403 , n5919 );
xor ( n11404 , n11402 , n11403 );
or ( n11405 , n11401 , n11404 );
buf ( n11406 , n4896 );
buf ( n11407 , n5920 );
xor ( n11408 , n11406 , n11407 );
or ( n11409 , n11405 , n11408 );
buf ( n11410 , n4897 );
buf ( n11411 , n5921 );
xor ( n11412 , n11410 , n11411 );
or ( n11413 , n11409 , n11412 );
buf ( n11414 , n4898 );
buf ( n11415 , n5922 );
xor ( n11416 , n11414 , n11415 );
or ( n11417 , n11413 , n11416 );
buf ( n11418 , n4899 );
buf ( n11419 , n5923 );
xor ( n11420 , n11418 , n11419 );
or ( n11421 , n11417 , n11420 );
buf ( n11422 , n4900 );
buf ( n11423 , n5924 );
xor ( n11424 , n11422 , n11423 );
or ( n11425 , n11421 , n11424 );
buf ( n11426 , n4901 );
buf ( n11427 , n5925 );
xor ( n11428 , n11426 , n11427 );
or ( n11429 , n11425 , n11428 );
buf ( n11430 , n4902 );
buf ( n11431 , n5926 );
xor ( n11432 , n11430 , n11431 );
or ( n11433 , n11429 , n11432 );
buf ( n11434 , n4903 );
buf ( n11435 , n5927 );
xor ( n11436 , n11434 , n11435 );
or ( n11437 , n11433 , n11436 );
buf ( n11438 , n4904 );
buf ( n11439 , n5928 );
xor ( n11440 , n11438 , n11439 );
or ( n11441 , n11437 , n11440 );
buf ( n11442 , n4905 );
buf ( n11443 , n5929 );
xor ( n11444 , n11442 , n11443 );
or ( n11445 , n11441 , n11444 );
buf ( n11446 , n4906 );
buf ( n11447 , n5930 );
xor ( n11448 , n11446 , n11447 );
or ( n11449 , n11445 , n11448 );
buf ( n11450 , n4907 );
buf ( n11451 , n5931 );
xor ( n11452 , n11450 , n11451 );
or ( n11453 , n11449 , n11452 );
buf ( n11454 , n4908 );
buf ( n11455 , n5932 );
xor ( n11456 , n11454 , n11455 );
or ( n11457 , n11453 , n11456 );
buf ( n11458 , n4909 );
buf ( n11459 , n5933 );
xor ( n11460 , n11458 , n11459 );
or ( n11461 , n11457 , n11460 );
buf ( n11462 , n4910 );
buf ( n11463 , n5934 );
xor ( n11464 , n11462 , n11463 );
or ( n11465 , n11461 , n11464 );
buf ( n11466 , n4911 );
buf ( n11467 , n5935 );
xor ( n11468 , n11466 , n11467 );
or ( n11469 , n11465 , n11468 );
buf ( n11470 , n4912 );
buf ( n11471 , n5936 );
xor ( n11472 , n11470 , n11471 );
or ( n11473 , n11469 , n11472 );
buf ( n11474 , n4913 );
buf ( n11475 , n5937 );
xor ( n11476 , n11474 , n11475 );
or ( n11477 , n11473 , n11476 );
buf ( n11478 , n4914 );
buf ( n11479 , n5938 );
xor ( n11480 , n11478 , n11479 );
or ( n11481 , n11477 , n11480 );
buf ( n11482 , n4915 );
buf ( n11483 , n5939 );
xor ( n11484 , n11482 , n11483 );
or ( n11485 , n11481 , n11484 );
buf ( n11486 , n4916 );
buf ( n11487 , n5940 );
xor ( n11488 , n11486 , n11487 );
or ( n11489 , n11485 , n11488 );
buf ( n11490 , n4917 );
buf ( n11491 , n5941 );
xor ( n11492 , n11490 , n11491 );
or ( n11493 , n11489 , n11492 );
buf ( n11494 , n4918 );
buf ( n11495 , n5942 );
xor ( n11496 , n11494 , n11495 );
or ( n11497 , n11493 , n11496 );
buf ( n11498 , n4919 );
buf ( n11499 , n5943 );
xor ( n11500 , n11498 , n11499 );
or ( n11501 , n11497 , n11500 );
buf ( n11502 , n4920 );
buf ( n11503 , n5944 );
xor ( n11504 , n11502 , n11503 );
or ( n11505 , n11501 , n11504 );
buf ( n11506 , n4921 );
buf ( n11507 , n5945 );
xor ( n11508 , n11506 , n11507 );
or ( n11509 , n11505 , n11508 );
buf ( n11510 , n4922 );
buf ( n11511 , n5946 );
xor ( n11512 , n11510 , n11511 );
or ( n11513 , n11509 , n11512 );
buf ( n11514 , n4923 );
buf ( n11515 , n5947 );
xor ( n11516 , n11514 , n11515 );
or ( n11517 , n11513 , n11516 );
buf ( n11518 , n4924 );
buf ( n11519 , n5948 );
xor ( n11520 , n11518 , n11519 );
or ( n11521 , n11517 , n11520 );
buf ( n11522 , n4925 );
buf ( n11523 , n5949 );
xor ( n11524 , n11522 , n11523 );
or ( n11525 , n11521 , n11524 );
buf ( n11526 , n4926 );
buf ( n11527 , n5950 );
xor ( n11528 , n11526 , n11527 );
or ( n11529 , n11525 , n11528 );
buf ( n11530 , n4927 );
buf ( n11531 , n5951 );
xor ( n11532 , n11530 , n11531 );
or ( n11533 , n11529 , n11532 );
buf ( n11534 , n4928 );
buf ( n11535 , n5952 );
xor ( n11536 , n11534 , n11535 );
or ( n11537 , n11533 , n11536 );
buf ( n11538 , n4929 );
buf ( n11539 , n5953 );
xor ( n11540 , n11538 , n11539 );
or ( n11541 , n11537 , n11540 );
buf ( n11542 , n4930 );
buf ( n11543 , n5954 );
xor ( n11544 , n11542 , n11543 );
or ( n11545 , n11541 , n11544 );
buf ( n11546 , n4931 );
buf ( n11547 , n5955 );
xor ( n11548 , n11546 , n11547 );
or ( n11549 , n11545 , n11548 );
buf ( n11550 , n4932 );
buf ( n11551 , n5956 );
xor ( n11552 , n11550 , n11551 );
or ( n11553 , n11549 , n11552 );
buf ( n11554 , n4933 );
buf ( n11555 , n5957 );
xor ( n11556 , n11554 , n11555 );
or ( n11557 , n11553 , n11556 );
buf ( n11558 , n4934 );
buf ( n11559 , n5958 );
xor ( n11560 , n11558 , n11559 );
or ( n11561 , n11557 , n11560 );
buf ( n11562 , n4935 );
buf ( n11563 , n5959 );
xor ( n11564 , n11562 , n11563 );
or ( n11565 , n11561 , n11564 );
buf ( n11566 , n4936 );
buf ( n11567 , n5960 );
xor ( n11568 , n11566 , n11567 );
or ( n11569 , n11565 , n11568 );
buf ( n11570 , n4937 );
buf ( n11571 , n5961 );
xor ( n11572 , n11570 , n11571 );
or ( n11573 , n11569 , n11572 );
buf ( n11574 , n4938 );
buf ( n11575 , n5962 );
xor ( n11576 , n11574 , n11575 );
or ( n11577 , n11573 , n11576 );
buf ( n11578 , n4939 );
buf ( n11579 , n5963 );
xor ( n11580 , n11578 , n11579 );
or ( n11581 , n11577 , n11580 );
buf ( n11582 , n4940 );
buf ( n11583 , n5964 );
xor ( n11584 , n11582 , n11583 );
or ( n11585 , n11581 , n11584 );
buf ( n11586 , n4941 );
buf ( n11587 , n5965 );
xor ( n11588 , n11586 , n11587 );
or ( n11589 , n11585 , n11588 );
buf ( n11590 , n4942 );
buf ( n11591 , n5966 );
xor ( n11592 , n11590 , n11591 );
or ( n11593 , n11589 , n11592 );
buf ( n11594 , n4943 );
buf ( n11595 , n5967 );
xor ( n11596 , n11594 , n11595 );
or ( n11597 , n11593 , n11596 );
buf ( n11598 , n4944 );
buf ( n11599 , n5968 );
xor ( n11600 , n11598 , n11599 );
or ( n11601 , n11597 , n11600 );
buf ( n11602 , n4945 );
buf ( n11603 , n5969 );
xor ( n11604 , n11602 , n11603 );
or ( n11605 , n11601 , n11604 );
buf ( n11606 , n4946 );
buf ( n11607 , n5970 );
xor ( n11608 , n11606 , n11607 );
or ( n11609 , n11605 , n11608 );
buf ( n11610 , n4947 );
buf ( n11611 , n5971 );
xor ( n11612 , n11610 , n11611 );
or ( n11613 , n11609 , n11612 );
buf ( n11614 , n4948 );
buf ( n11615 , n5972 );
xor ( n11616 , n11614 , n11615 );
or ( n11617 , n11613 , n11616 );
buf ( n11618 , n4949 );
buf ( n11619 , n5973 );
xor ( n11620 , n11618 , n11619 );
or ( n11621 , n11617 , n11620 );
buf ( n11622 , n4950 );
buf ( n11623 , n5974 );
xor ( n11624 , n11622 , n11623 );
or ( n11625 , n11621 , n11624 );
buf ( n11626 , n4951 );
buf ( n11627 , n5975 );
xor ( n11628 , n11626 , n11627 );
or ( n11629 , n11625 , n11628 );
buf ( n11630 , n4952 );
buf ( n11631 , n5976 );
xor ( n11632 , n11630 , n11631 );
or ( n11633 , n11629 , n11632 );
buf ( n11634 , n4953 );
buf ( n11635 , n5977 );
xor ( n11636 , n11634 , n11635 );
or ( n11637 , n11633 , n11636 );
buf ( n11638 , n4954 );
buf ( n11639 , n5978 );
xor ( n11640 , n11638 , n11639 );
or ( n11641 , n11637 , n11640 );
buf ( n11642 , n4955 );
buf ( n11643 , n5979 );
xor ( n11644 , n11642 , n11643 );
or ( n11645 , n11641 , n11644 );
buf ( n11646 , n4956 );
buf ( n11647 , n5980 );
xor ( n11648 , n11646 , n11647 );
or ( n11649 , n11645 , n11648 );
buf ( n11650 , n4957 );
buf ( n11651 , n5981 );
xor ( n11652 , n11650 , n11651 );
or ( n11653 , n11649 , n11652 );
buf ( n11654 , n4958 );
buf ( n11655 , n5982 );
xor ( n11656 , n11654 , n11655 );
or ( n11657 , n11653 , n11656 );
buf ( n11658 , n4959 );
buf ( n11659 , n5983 );
xor ( n11660 , n11658 , n11659 );
or ( n11661 , n11657 , n11660 );
buf ( n11662 , n4960 );
buf ( n11663 , n5984 );
xor ( n11664 , n11662 , n11663 );
or ( n11665 , n11661 , n11664 );
buf ( n11666 , n4961 );
buf ( n11667 , n5985 );
xor ( n11668 , n11666 , n11667 );
or ( n11669 , n11665 , n11668 );
buf ( n11670 , n4962 );
buf ( n11671 , n5986 );
xor ( n11672 , n11670 , n11671 );
or ( n11673 , n11669 , n11672 );
buf ( n11674 , n4963 );
buf ( n11675 , n5987 );
xor ( n11676 , n11674 , n11675 );
or ( n11677 , n11673 , n11676 );
buf ( n11678 , n4964 );
buf ( n11679 , n5988 );
xor ( n11680 , n11678 , n11679 );
or ( n11681 , n11677 , n11680 );
buf ( n11682 , n4965 );
buf ( n11683 , n5989 );
xor ( n11684 , n11682 , n11683 );
or ( n11685 , n11681 , n11684 );
buf ( n11686 , n4966 );
buf ( n11687 , n5990 );
xor ( n11688 , n11686 , n11687 );
or ( n11689 , n11685 , n11688 );
buf ( n11690 , n4967 );
buf ( n11691 , n5991 );
xor ( n11692 , n11690 , n11691 );
or ( n11693 , n11689 , n11692 );
buf ( n11694 , n4968 );
buf ( n11695 , n5992 );
xor ( n11696 , n11694 , n11695 );
or ( n11697 , n11693 , n11696 );
buf ( n11698 , n4969 );
buf ( n11699 , n5993 );
xor ( n11700 , n11698 , n11699 );
or ( n11701 , n11697 , n11700 );
buf ( n11702 , n4970 );
buf ( n11703 , n5994 );
xor ( n11704 , n11702 , n11703 );
or ( n11705 , n11701 , n11704 );
buf ( n11706 , n4971 );
buf ( n11707 , n5995 );
xor ( n11708 , n11706 , n11707 );
or ( n11709 , n11705 , n11708 );
buf ( n11710 , n4972 );
buf ( n11711 , n5996 );
xor ( n11712 , n11710 , n11711 );
or ( n11713 , n11709 , n11712 );
buf ( n11714 , n4973 );
buf ( n11715 , n5997 );
xor ( n11716 , n11714 , n11715 );
or ( n11717 , n11713 , n11716 );
buf ( n11718 , n4974 );
buf ( n11719 , n5998 );
xor ( n11720 , n11718 , n11719 );
or ( n11721 , n11717 , n11720 );
buf ( n11722 , n4975 );
buf ( n11723 , n5999 );
xor ( n11724 , n11722 , n11723 );
or ( n11725 , n11721 , n11724 );
buf ( n11726 , n4976 );
buf ( n11727 , n6000 );
xor ( n11728 , n11726 , n11727 );
or ( n11729 , n11725 , n11728 );
buf ( n11730 , n4977 );
buf ( n11731 , n6001 );
xor ( n11732 , n11730 , n11731 );
or ( n11733 , n11729 , n11732 );
buf ( n11734 , n4978 );
buf ( n11735 , n6002 );
xor ( n11736 , n11734 , n11735 );
or ( n11737 , n11733 , n11736 );
buf ( n11738 , n4979 );
buf ( n11739 , n6003 );
xor ( n11740 , n11738 , n11739 );
or ( n11741 , n11737 , n11740 );
buf ( n11742 , n4980 );
buf ( n11743 , n6004 );
xor ( n11744 , n11742 , n11743 );
or ( n11745 , n11741 , n11744 );
buf ( n11746 , n4981 );
buf ( n11747 , n6005 );
xor ( n11748 , n11746 , n11747 );
or ( n11749 , n11745 , n11748 );
buf ( n11750 , n4982 );
buf ( n11751 , n6006 );
xor ( n11752 , n11750 , n11751 );
or ( n11753 , n11749 , n11752 );
buf ( n11754 , n4983 );
buf ( n11755 , n6007 );
xor ( n11756 , n11754 , n11755 );
or ( n11757 , n11753 , n11756 );
buf ( n11758 , n4984 );
buf ( n11759 , n6008 );
xor ( n11760 , n11758 , n11759 );
or ( n11761 , n11757 , n11760 );
buf ( n11762 , n4985 );
buf ( n11763 , n6009 );
xor ( n11764 , n11762 , n11763 );
or ( n11765 , n11761 , n11764 );
buf ( n11766 , n4986 );
buf ( n11767 , n6010 );
xor ( n11768 , n11766 , n11767 );
or ( n11769 , n11765 , n11768 );
buf ( n11770 , n4987 );
buf ( n11771 , n6011 );
xor ( n11772 , n11770 , n11771 );
or ( n11773 , n11769 , n11772 );
buf ( n11774 , n4988 );
buf ( n11775 , n6012 );
xor ( n11776 , n11774 , n11775 );
or ( n11777 , n11773 , n11776 );
buf ( n11778 , n4989 );
buf ( n11779 , n6013 );
xor ( n11780 , n11778 , n11779 );
or ( n11781 , n11777 , n11780 );
buf ( n11782 , n4990 );
buf ( n11783 , n6014 );
xor ( n11784 , n11782 , n11783 );
or ( n11785 , n11781 , n11784 );
buf ( n11786 , n4991 );
buf ( n11787 , n6015 );
xor ( n11788 , n11786 , n11787 );
or ( n11789 , n11785 , n11788 );
buf ( n11790 , n4992 );
buf ( n11791 , n6016 );
xor ( n11792 , n11790 , n11791 );
or ( n11793 , n11789 , n11792 );
buf ( n11794 , n4993 );
buf ( n11795 , n6017 );
xor ( n11796 , n11794 , n11795 );
or ( n11797 , n11793 , n11796 );
buf ( n11798 , n4994 );
buf ( n11799 , n6018 );
xor ( n11800 , n11798 , n11799 );
or ( n11801 , n11797 , n11800 );
buf ( n11802 , n4995 );
buf ( n11803 , n6019 );
xor ( n11804 , n11802 , n11803 );
or ( n11805 , n11801 , n11804 );
buf ( n11806 , n4996 );
buf ( n11807 , n6020 );
xor ( n11808 , n11806 , n11807 );
or ( n11809 , n11805 , n11808 );
buf ( n11810 , n4997 );
buf ( n11811 , n6021 );
xor ( n11812 , n11810 , n11811 );
or ( n11813 , n11809 , n11812 );
buf ( n11814 , n4998 );
buf ( n11815 , n6022 );
xor ( n11816 , n11814 , n11815 );
or ( n11817 , n11813 , n11816 );
buf ( n11818 , n4999 );
buf ( n11819 , n6023 );
xor ( n11820 , n11818 , n11819 );
or ( n11821 , n11817 , n11820 );
buf ( n11822 , n5000 );
buf ( n11823 , n6024 );
xor ( n11824 , n11822 , n11823 );
or ( n11825 , n11821 , n11824 );
buf ( n11826 , n5001 );
buf ( n11827 , n6025 );
xor ( n11828 , n11826 , n11827 );
or ( n11829 , n11825 , n11828 );
buf ( n11830 , n5002 );
buf ( n11831 , n6026 );
xor ( n11832 , n11830 , n11831 );
or ( n11833 , n11829 , n11832 );
buf ( n11834 , n5003 );
buf ( n11835 , n6027 );
xor ( n11836 , n11834 , n11835 );
or ( n11837 , n11833 , n11836 );
buf ( n11838 , n5004 );
buf ( n11839 , n6028 );
xor ( n11840 , n11838 , n11839 );
or ( n11841 , n11837 , n11840 );
buf ( n11842 , n5005 );
buf ( n11843 , n6029 );
xor ( n11844 , n11842 , n11843 );
or ( n11845 , n11841 , n11844 );
buf ( n11846 , n5006 );
buf ( n11847 , n6030 );
xor ( n11848 , n11846 , n11847 );
or ( n11849 , n11845 , n11848 );
buf ( n11850 , n5007 );
buf ( n11851 , n6031 );
xor ( n11852 , n11850 , n11851 );
or ( n11853 , n11849 , n11852 );
buf ( n11854 , n5008 );
buf ( n11855 , n6032 );
xor ( n11856 , n11854 , n11855 );
or ( n11857 , n11853 , n11856 );
buf ( n11858 , n5009 );
buf ( n11859 , n6033 );
xor ( n11860 , n11858 , n11859 );
or ( n11861 , n11857 , n11860 );
buf ( n11862 , n5010 );
buf ( n11863 , n6034 );
xor ( n11864 , n11862 , n11863 );
or ( n11865 , n11861 , n11864 );
buf ( n11866 , n5011 );
buf ( n11867 , n6035 );
xor ( n11868 , n11866 , n11867 );
or ( n11869 , n11865 , n11868 );
buf ( n11870 , n5012 );
buf ( n11871 , n6036 );
xor ( n11872 , n11870 , n11871 );
or ( n11873 , n11869 , n11872 );
buf ( n11874 , n5013 );
buf ( n11875 , n6037 );
xor ( n11876 , n11874 , n11875 );
or ( n11877 , n11873 , n11876 );
buf ( n11878 , n5014 );
buf ( n11879 , n6038 );
xor ( n11880 , n11878 , n11879 );
or ( n11881 , n11877 , n11880 );
buf ( n11882 , n5015 );
buf ( n11883 , n6039 );
xor ( n11884 , n11882 , n11883 );
or ( n11885 , n11881 , n11884 );
buf ( n11886 , n5016 );
buf ( n11887 , n6040 );
xor ( n11888 , n11886 , n11887 );
or ( n11889 , n11885 , n11888 );
buf ( n11890 , n5017 );
buf ( n11891 , n6041 );
xor ( n11892 , n11890 , n11891 );
or ( n11893 , n11889 , n11892 );
buf ( n11894 , n5018 );
buf ( n11895 , n6042 );
xor ( n11896 , n11894 , n11895 );
or ( n11897 , n11893 , n11896 );
buf ( n11898 , n5019 );
buf ( n11899 , n6043 );
xor ( n11900 , n11898 , n11899 );
or ( n11901 , n11897 , n11900 );
buf ( n11902 , n5020 );
buf ( n11903 , n6044 );
xor ( n11904 , n11902 , n11903 );
or ( n11905 , n11901 , n11904 );
buf ( n11906 , n5021 );
buf ( n11907 , n6045 );
xor ( n11908 , n11906 , n11907 );
or ( n11909 , n11905 , n11908 );
buf ( n11910 , n5022 );
buf ( n11911 , n6046 );
xor ( n11912 , n11910 , n11911 );
or ( n11913 , n11909 , n11912 );
buf ( n11914 , n5023 );
buf ( n11915 , n6047 );
xor ( n11916 , n11914 , n11915 );
or ( n11917 , n11913 , n11916 );
buf ( n11918 , n5024 );
buf ( n11919 , n6048 );
xor ( n11920 , n11918 , n11919 );
or ( n11921 , n11917 , n11920 );
buf ( n11922 , n5025 );
buf ( n11923 , n6049 );
xor ( n11924 , n11922 , n11923 );
or ( n11925 , n11921 , n11924 );
buf ( n11926 , n5026 );
buf ( n11927 , n6050 );
xor ( n11928 , n11926 , n11927 );
or ( n11929 , n11925 , n11928 );
buf ( n11930 , n5027 );
buf ( n11931 , n6051 );
xor ( n11932 , n11930 , n11931 );
or ( n11933 , n11929 , n11932 );
buf ( n11934 , n5028 );
buf ( n11935 , n6052 );
xor ( n11936 , n11934 , n11935 );
or ( n11937 , n11933 , n11936 );
buf ( n11938 , n5029 );
buf ( n11939 , n6053 );
xor ( n11940 , n11938 , n11939 );
or ( n11941 , n11937 , n11940 );
buf ( n11942 , n5030 );
buf ( n11943 , n6054 );
xor ( n11944 , n11942 , n11943 );
or ( n11945 , n11941 , n11944 );
buf ( n11946 , n5031 );
buf ( n11947 , n6055 );
xor ( n11948 , n11946 , n11947 );
or ( n11949 , n11945 , n11948 );
buf ( n11950 , n5032 );
buf ( n11951 , n6056 );
xor ( n11952 , n11950 , n11951 );
or ( n11953 , n11949 , n11952 );
buf ( n11954 , n5033 );
buf ( n11955 , n6057 );
xor ( n11956 , n11954 , n11955 );
or ( n11957 , n11953 , n11956 );
buf ( n11958 , n5034 );
buf ( n11959 , n6058 );
xor ( n11960 , n11958 , n11959 );
or ( n11961 , n11957 , n11960 );
buf ( n11962 , n5035 );
buf ( n11963 , n6059 );
xor ( n11964 , n11962 , n11963 );
or ( n11965 , n11961 , n11964 );
buf ( n11966 , n5036 );
buf ( n11967 , n6060 );
xor ( n11968 , n11966 , n11967 );
or ( n11969 , n11965 , n11968 );
buf ( n11970 , n5037 );
buf ( n11971 , n6061 );
xor ( n11972 , n11970 , n11971 );
or ( n11973 , n11969 , n11972 );
buf ( n11974 , n5038 );
buf ( n11975 , n6062 );
xor ( n11976 , n11974 , n11975 );
or ( n11977 , n11973 , n11976 );
buf ( n11978 , n5039 );
buf ( n11979 , n6063 );
xor ( n11980 , n11978 , n11979 );
or ( n11981 , n11977 , n11980 );
buf ( n11982 , n5040 );
buf ( n11983 , n6064 );
xor ( n11984 , n11982 , n11983 );
or ( n11985 , n11981 , n11984 );
buf ( n11986 , n5041 );
buf ( n11987 , n6065 );
xor ( n11988 , n11986 , n11987 );
or ( n11989 , n11985 , n11988 );
buf ( n11990 , n5042 );
buf ( n11991 , n6066 );
xor ( n11992 , n11990 , n11991 );
or ( n11993 , n11989 , n11992 );
buf ( n11994 , n5043 );
buf ( n11995 , n6067 );
xor ( n11996 , n11994 , n11995 );
or ( n11997 , n11993 , n11996 );
buf ( n11998 , n5044 );
buf ( n11999 , n6068 );
xor ( n12000 , n11998 , n11999 );
or ( n12001 , n11997 , n12000 );
buf ( n12002 , n5045 );
buf ( n12003 , n6069 );
xor ( n12004 , n12002 , n12003 );
or ( n12005 , n12001 , n12004 );
buf ( n12006 , n5046 );
buf ( n12007 , n6070 );
xor ( n12008 , n12006 , n12007 );
or ( n12009 , n12005 , n12008 );
buf ( n12010 , n5047 );
buf ( n12011 , n6071 );
xor ( n12012 , n12010 , n12011 );
or ( n12013 , n12009 , n12012 );
buf ( n12014 , n5048 );
buf ( n12015 , n6072 );
xor ( n12016 , n12014 , n12015 );
or ( n12017 , n12013 , n12016 );
buf ( n12018 , n5049 );
buf ( n12019 , n6073 );
xor ( n12020 , n12018 , n12019 );
or ( n12021 , n12017 , n12020 );
buf ( n12022 , n5050 );
buf ( n12023 , n6074 );
xor ( n12024 , n12022 , n12023 );
or ( n12025 , n12021 , n12024 );
buf ( n12026 , n5051 );
buf ( n12027 , n6075 );
xor ( n12028 , n12026 , n12027 );
or ( n12029 , n12025 , n12028 );
buf ( n12030 , n5052 );
buf ( n12031 , n6076 );
xor ( n12032 , n12030 , n12031 );
or ( n12033 , n12029 , n12032 );
buf ( n12034 , n5053 );
buf ( n12035 , n6077 );
xor ( n12036 , n12034 , n12035 );
or ( n12037 , n12033 , n12036 );
buf ( n12038 , n5054 );
buf ( n12039 , n6078 );
xor ( n12040 , n12038 , n12039 );
or ( n12041 , n12037 , n12040 );
buf ( n12042 , n5055 );
buf ( n12043 , n6079 );
xor ( n12044 , n12042 , n12043 );
or ( n12045 , n12041 , n12044 );
buf ( n12046 , n5056 );
buf ( n12047 , n6080 );
xor ( n12048 , n12046 , n12047 );
or ( n12049 , n12045 , n12048 );
buf ( n12050 , n5057 );
buf ( n12051 , n6081 );
xor ( n12052 , n12050 , n12051 );
or ( n12053 , n12049 , n12052 );
buf ( n12054 , n5058 );
buf ( n12055 , n6082 );
xor ( n12056 , n12054 , n12055 );
or ( n12057 , n12053 , n12056 );
buf ( n12058 , n5059 );
buf ( n12059 , n6083 );
xor ( n12060 , n12058 , n12059 );
or ( n12061 , n12057 , n12060 );
buf ( n12062 , n5060 );
buf ( n12063 , n6084 );
xor ( n12064 , n12062 , n12063 );
or ( n12065 , n12061 , n12064 );
buf ( n12066 , n5061 );
buf ( n12067 , n6085 );
xor ( n12068 , n12066 , n12067 );
or ( n12069 , n12065 , n12068 );
buf ( n12070 , n5062 );
buf ( n12071 , n6086 );
xor ( n12072 , n12070 , n12071 );
or ( n12073 , n12069 , n12072 );
buf ( n12074 , n5063 );
buf ( n12075 , n6087 );
xor ( n12076 , n12074 , n12075 );
or ( n12077 , n12073 , n12076 );
buf ( n12078 , n5064 );
buf ( n12079 , n6088 );
xor ( n12080 , n12078 , n12079 );
or ( n12081 , n12077 , n12080 );
buf ( n12082 , n5065 );
buf ( n12083 , n6089 );
xor ( n12084 , n12082 , n12083 );
or ( n12085 , n12081 , n12084 );
buf ( n12086 , n5066 );
buf ( n12087 , n6090 );
xor ( n12088 , n12086 , n12087 );
or ( n12089 , n12085 , n12088 );
buf ( n12090 , n5067 );
buf ( n12091 , n6091 );
xor ( n12092 , n12090 , n12091 );
or ( n12093 , n12089 , n12092 );
buf ( n12094 , n5068 );
buf ( n12095 , n6092 );
xor ( n12096 , n12094 , n12095 );
or ( n12097 , n12093 , n12096 );
buf ( n12098 , n5069 );
buf ( n12099 , n6093 );
xor ( n12100 , n12098 , n12099 );
or ( n12101 , n12097 , n12100 );
buf ( n12102 , n5070 );
buf ( n12103 , n6094 );
xor ( n12104 , n12102 , n12103 );
or ( n12105 , n12101 , n12104 );
buf ( n12106 , n5071 );
buf ( n12107 , n6095 );
xor ( n12108 , n12106 , n12107 );
or ( n12109 , n12105 , n12108 );
buf ( n12110 , n5072 );
buf ( n12111 , n6096 );
xor ( n12112 , n12110 , n12111 );
or ( n12113 , n12109 , n12112 );
buf ( n12114 , n5073 );
buf ( n12115 , n6097 );
xor ( n12116 , n12114 , n12115 );
or ( n12117 , n12113 , n12116 );
buf ( n12118 , n5074 );
buf ( n12119 , n6098 );
xor ( n12120 , n12118 , n12119 );
or ( n12121 , n12117 , n12120 );
buf ( n12122 , n5075 );
buf ( n12123 , n6099 );
xor ( n12124 , n12122 , n12123 );
or ( n12125 , n12121 , n12124 );
buf ( n12126 , n5076 );
buf ( n12127 , n6100 );
xor ( n12128 , n12126 , n12127 );
or ( n12129 , n12125 , n12128 );
buf ( n12130 , n5077 );
buf ( n12131 , n6101 );
xor ( n12132 , n12130 , n12131 );
or ( n12133 , n12129 , n12132 );
buf ( n12134 , n5078 );
buf ( n12135 , n6102 );
xor ( n12136 , n12134 , n12135 );
or ( n12137 , n12133 , n12136 );
buf ( n12138 , n5079 );
buf ( n12139 , n6103 );
xor ( n12140 , n12138 , n12139 );
or ( n12141 , n12137 , n12140 );
buf ( n12142 , n5080 );
buf ( n12143 , n6104 );
xor ( n12144 , n12142 , n12143 );
or ( n12145 , n12141 , n12144 );
buf ( n12146 , n5081 );
buf ( n12147 , n6105 );
xor ( n12148 , n12146 , n12147 );
or ( n12149 , n12145 , n12148 );
buf ( n12150 , n5082 );
buf ( n12151 , n6106 );
xor ( n12152 , n12150 , n12151 );
or ( n12153 , n12149 , n12152 );
buf ( n12154 , n5083 );
buf ( n12155 , n6107 );
xor ( n12156 , n12154 , n12155 );
or ( n12157 , n12153 , n12156 );
buf ( n12158 , n5084 );
buf ( n12159 , n6108 );
xor ( n12160 , n12158 , n12159 );
or ( n12161 , n12157 , n12160 );
buf ( n12162 , n5085 );
buf ( n12163 , n6109 );
xor ( n12164 , n12162 , n12163 );
or ( n12165 , n12161 , n12164 );
buf ( n12166 , n5086 );
buf ( n12167 , n6110 );
xor ( n12168 , n12166 , n12167 );
or ( n12169 , n12165 , n12168 );
buf ( n12170 , n5087 );
buf ( n12171 , n6111 );
xor ( n12172 , n12170 , n12171 );
or ( n12173 , n12169 , n12172 );
buf ( n12174 , n5088 );
buf ( n12175 , n6112 );
xor ( n12176 , n12174 , n12175 );
or ( n12177 , n12173 , n12176 );
buf ( n12178 , n5089 );
buf ( n12179 , n6113 );
xor ( n12180 , n12178 , n12179 );
or ( n12181 , n12177 , n12180 );
buf ( n12182 , n5090 );
buf ( n12183 , n6114 );
xor ( n12184 , n12182 , n12183 );
or ( n12185 , n12181 , n12184 );
buf ( n12186 , n5091 );
buf ( n12187 , n6115 );
xor ( n12188 , n12186 , n12187 );
or ( n12189 , n12185 , n12188 );
buf ( n12190 , n5092 );
buf ( n12191 , n6116 );
xor ( n12192 , n12190 , n12191 );
or ( n12193 , n12189 , n12192 );
buf ( n12194 , n5093 );
buf ( n12195 , n6117 );
xor ( n12196 , n12194 , n12195 );
or ( n12197 , n12193 , n12196 );
buf ( n12198 , n5094 );
buf ( n12199 , n6118 );
xor ( n12200 , n12198 , n12199 );
or ( n12201 , n12197 , n12200 );
buf ( n12202 , n5095 );
buf ( n12203 , n6119 );
xor ( n12204 , n12202 , n12203 );
or ( n12205 , n12201 , n12204 );
buf ( n12206 , n5096 );
buf ( n12207 , n6120 );
xor ( n12208 , n12206 , n12207 );
or ( n12209 , n12205 , n12208 );
buf ( n12210 , n5097 );
buf ( n12211 , n6121 );
xor ( n12212 , n12210 , n12211 );
or ( n12213 , n12209 , n12212 );
buf ( n12214 , n5098 );
buf ( n12215 , n6122 );
xor ( n12216 , n12214 , n12215 );
or ( n12217 , n12213 , n12216 );
buf ( n12218 , n5099 );
buf ( n12219 , n6123 );
xor ( n12220 , n12218 , n12219 );
or ( n12221 , n12217 , n12220 );
buf ( n12222 , n5100 );
buf ( n12223 , n6124 );
xor ( n12224 , n12222 , n12223 );
or ( n12225 , n12221 , n12224 );
buf ( n12226 , n5101 );
buf ( n12227 , n6125 );
xor ( n12228 , n12226 , n12227 );
or ( n12229 , n12225 , n12228 );
buf ( n12230 , n5102 );
buf ( n12231 , n6126 );
xor ( n12232 , n12230 , n12231 );
or ( n12233 , n12229 , n12232 );
buf ( n12234 , n5103 );
buf ( n12235 , n6127 );
xor ( n12236 , n12234 , n12235 );
or ( n12237 , n12233 , n12236 );
buf ( n12238 , n5104 );
buf ( n12239 , n6128 );
xor ( n12240 , n12238 , n12239 );
or ( n12241 , n12237 , n12240 );
buf ( n12242 , n5105 );
buf ( n12243 , n6129 );
xor ( n12244 , n12242 , n12243 );
or ( n12245 , n12241 , n12244 );
buf ( n12246 , n5106 );
buf ( n12247 , n6130 );
xor ( n12248 , n12246 , n12247 );
or ( n12249 , n12245 , n12248 );
buf ( n12250 , n5107 );
buf ( n12251 , n6131 );
xor ( n12252 , n12250 , n12251 );
or ( n12253 , n12249 , n12252 );
buf ( n12254 , n5108 );
buf ( n12255 , n6132 );
xor ( n12256 , n12254 , n12255 );
or ( n12257 , n12253 , n12256 );
buf ( n12258 , n5109 );
not ( n12259 , n12258 );
or ( n12260 , n12257 , n12259 );
buf ( n12261 , n5110 );
buf ( n12262 , n6134 );
xor ( n12263 , n12261 , n12262 );
or ( n12264 , n12260 , n12263 );
buf ( n12265 , n5111 );
not ( n12266 , n12265 );
or ( n12267 , n12264 , n12266 );
buf ( n12268 , n5112 );
not ( n12269 , n12268 );
or ( n12270 , n12267 , n12269 );
buf ( n12271 , n5113 );
buf ( n12272 , n6137 );
xor ( n12273 , n12271 , n12272 );
or ( n12274 , n12270 , n12273 );
buf ( n12275 , n5114 );
buf ( n12276 , n6138 );
xor ( n12277 , n12275 , n12276 );
or ( n12278 , n12274 , n12277 );
buf ( n12279 , n5115 );
buf ( n12280 , n6139 );
xor ( n12281 , n12279 , n12280 );
or ( n12282 , n12278 , n12281 );
buf ( n12283 , n5116 );
not ( n12284 , n12283 );
or ( n12285 , n12282 , n12284 );
buf ( n12286 , n5117 );
not ( n12287 , n12286 );
or ( n12288 , n12285 , n12287 );
buf ( n12289 , n5118 );
buf ( n12290 , n6142 );
xor ( n12291 , n12289 , n12290 );
or ( n12292 , n12288 , n12291 );
buf ( n12293 , n5119 );
not ( n12294 , n12293 );
or ( n12295 , n12292 , n12294 );
buf ( n12296 , n5120 );
not ( n12297 , n12296 );
or ( n12298 , n12295 , n12297 );
buf ( n12299 , n5121 );
not ( n12300 , n12299 );
or ( n12301 , n12298 , n12300 );
buf ( n12302 , n5122 );
not ( n12303 , n12302 );
or ( n12304 , n12301 , n12303 );
buf ( n12305 , n5123 );
buf ( n12306 , n6147 );
xor ( n12307 , n12305 , n12306 );
or ( n12308 , n12304 , n12307 );
buf ( n12309 , n5124 );
buf ( n12310 , n6148 );
xor ( n12311 , n12309 , n12310 );
or ( n12312 , n12308 , n12311 );
buf ( n12313 , n5125 );
buf ( n12314 , n6149 );
xor ( n12315 , n12313 , n12314 );
or ( n12316 , n12312 , n12315 );
not ( n12317 , n12316 );
buf ( n12318 , n12317 );
buf ( n12319 , n12318 );
endmodule

