//
// Conformal-LEC Version 16.10-d005 ( 21-Apr-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 ;
output n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 ;

wire n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , 
     n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , 
     n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , 
     n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , 
     n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , 
     n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , 
     n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , 
     n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , 
     n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , 
     n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , 
     n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , 
     n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , 
     n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , 
     n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , 
     n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , 
     n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , 
     n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , 
     n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , 
     n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , 
     n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , 
     n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , 
     n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , 
     n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , 
     n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , 
     n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , 
     n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , 
     n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , 
     n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , 
     n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , 
     n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , 
     n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , 
     n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , 
     n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , 
     n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , 
     n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , 
     n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , 
     n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , 
     n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , 
     n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , 
     n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , 
     n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , 
     n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , 
     n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , 
     n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , 
     n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , 
     n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , 
     n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , 
     n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , 
     n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , 
     n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , 
     n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , 
     n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , 
     n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , 
     n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , 
     n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , 
     n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , 
     n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , 
     n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , 
     n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , 
     n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , 
     n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , 
     n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , 
     n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , 
     n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , 
     n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , 
     n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , 
     n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , 
     n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , 
     n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , 
     n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , 
     n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , 
     n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , 
     n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , 
     n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , 
     n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , 
     n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , 
     n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , 
     n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , 
     n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , 
     n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , 
     n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , 
     n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , 
     n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , 
     n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , 
     n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , 
     n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , 
     n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , 
     n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , 
     n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , 
     n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , 
     n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , 
     n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , 
     n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , 
     n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , 
     n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , 
     n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , 
     n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , 
     n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , 
     n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , 
     n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , 
     n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , 
     n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , 
     n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , 
     n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , 
     n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , 
     n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , 
     n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , 
     n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , 
     n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , 
     n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , 
     n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , 
     n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , 
     n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , 
     n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , 
     n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , 
     n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , 
     n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , 
     n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , 
     n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , 
     n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , 
     n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , 
     n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , 
     n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , 
     n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , 
     n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , 
     n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , 
     n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , 
     n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , 
     n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , 
     n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , 
     n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , 
     n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , 
     n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , 
     n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , 
     n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , 
     n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , 
     n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , 
     n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , 
     n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , 
     n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , 
     n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , 
     n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , 
     n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , 
     n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , 
     n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , 
     n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , 
     n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , 
     n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , 
     n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , 
     n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , 
     n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , 
     n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , 
     n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , 
     n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , 
     n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , 
     n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , 
     n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , 
     n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , 
     n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , 
     n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , 
     n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , 
     n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , 
     n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , 
     n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , 
     n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , 
     n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , 
     n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , 
     n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , 
     n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , 
     n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , 
     n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , 
     n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , 
     n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , 
     n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , 
     n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , 
     n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , 
     n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , 
     n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , 
     n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , 
     n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , 
     n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , 
     n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , 
     n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , 
     n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , 
     n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , 
     n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , 
     n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , 
     n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , 
     n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , 
     n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , 
     n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , 
     n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , 
     n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , 
     n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , 
     n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , 
     n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , 
     n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , 
     n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , 
     n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , 
     n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , 
     n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , 
     n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , 
     n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , 
     n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , 
     n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , 
     n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , 
     n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , 
     n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , 
     n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , 
     n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , 
     n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , 
     n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , 
     n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , 
     n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , 
     n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , 
     n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , 
     n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , 
     n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , 
     n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , 
     n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , 
     n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , 
     n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , 
     n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , 
     n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , 
     n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , 
     n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , 
     n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , 
     n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , 
     n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , 
     n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , 
     n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , 
     n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , 
     n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , 
     n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , 
     n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , 
     n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , 
     n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , 
     n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , 
     n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , 
     n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , 
     n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , 
     n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , 
     n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , 
     n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , 
     n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , 
     n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , 
     n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , 
     n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , 
     n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , 
     n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , 
     n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , 
     n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , 
     n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , 
     n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , 
     n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , 
     n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , 
     n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , 
     n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , 
     n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , 
     n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , 
     n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , 
     n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , 
     n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , 
     n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , 
     n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , 
     n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , 
     n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , 
     n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , 
     n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , 
     n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , 
     n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , 
     n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , 
     n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , 
     n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , 
     n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , 
     n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , 
     n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , 
     n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , 
     n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , 
     n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , 
     n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , 
     n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , 
     n3223 , n3224 ;
buf ( n195 , n1861 );
buf ( n194 , n2305 );
buf ( n196 , n2369 );
buf ( n197 , n2427 );
buf ( n199 , n2757 );
buf ( n201 , n2888 );
buf ( n200 , n2976 );
buf ( n192 , n3041 );
buf ( n193 , n3111 );
buf ( n198 , n3224 );
buf ( n406 , n136 );
buf ( n407 , n25 );
buf ( n408 , n94 );
buf ( n409 , n2 );
buf ( n410 , n132 );
buf ( n411 , n156 );
buf ( n412 , n114 );
buf ( n413 , n159 );
buf ( n414 , n67 );
buf ( n415 , n184 );
buf ( n416 , n111 );
buf ( n417 , n130 );
buf ( n418 , n181 );
buf ( n419 , n52 );
buf ( n420 , n166 );
buf ( n421 , n153 );
buf ( n422 , n131 );
buf ( n423 , n141 );
buf ( n424 , n140 );
buf ( n425 , n9 );
buf ( n426 , n71 );
buf ( n427 , n113 );
buf ( n428 , n43 );
buf ( n429 , n126 );
buf ( n430 , n137 );
buf ( n431 , n22 );
buf ( n432 , n150 );
buf ( n433 , n104 );
buf ( n434 , n73 );
buf ( n435 , n100 );
buf ( n436 , n180 );
buf ( n437 , n167 );
buf ( n438 , n135 );
buf ( n439 , n178 );
buf ( n440 , n106 );
buf ( n441 , n57 );
buf ( n442 , n69 );
buf ( n443 , n175 );
buf ( n444 , n15 );
buf ( n445 , n152 );
buf ( n446 , n24 );
buf ( n447 , n70 );
buf ( n448 , n115 );
buf ( n449 , n68 );
buf ( n450 , n50 );
buf ( n451 , n134 );
buf ( n452 , n4 );
buf ( n453 , n31 );
buf ( n454 , n146 );
buf ( n455 , n59 );
buf ( n456 , n38 );
buf ( n457 , n138 );
buf ( n458 , n0 );
buf ( n459 , n95 );
buf ( n460 , n75 );
buf ( n461 , n60 );
buf ( n462 , n168 );
buf ( n463 , n157 );
buf ( n464 , n169 );
buf ( n465 , n21 );
buf ( n466 , n89 );
buf ( n467 , n92 );
buf ( n468 , n26 );
buf ( n469 , n51 );
buf ( n470 , n34 );
buf ( n471 , n124 );
buf ( n472 , n82 );
buf ( n473 , n62 );
buf ( n474 , n40 );
buf ( n475 , n125 );
buf ( n476 , n54 );
buf ( n477 , n107 );
buf ( n478 , n116 );
buf ( n479 , n88 );
buf ( n480 , n117 );
buf ( n481 , n173 );
buf ( n482 , n127 );
buf ( n483 , n63 );
buf ( n484 , n123 );
buf ( n485 , n1 );
buf ( n486 , n84 );
buf ( n487 , n66 );
buf ( n488 , n7 );
buf ( n489 , n165 );
buf ( n490 , n45 );
buf ( n491 , n163 );
buf ( n492 , n172 );
buf ( n493 , n19 );
buf ( n494 , n171 );
buf ( n495 , n182 );
buf ( n496 , n147 );
buf ( n497 , n55 );
buf ( n498 , n154 );
buf ( n499 , n109 );
buf ( n500 , n121 );
buf ( n501 , n10 );
buf ( n502 , n191 );
buf ( n503 , n122 );
buf ( n504 , n41 );
buf ( n505 , n77 );
buf ( n506 , n98 );
buf ( n507 , n118 );
buf ( n508 , n164 );
buf ( n509 , n44 );
buf ( n510 , n78 );
buf ( n511 , n83 );
buf ( n512 , n129 );
buf ( n513 , n161 );
buf ( n514 , n103 );
buf ( n515 , n33 );
buf ( n516 , n188 );
buf ( n517 , n46 );
buf ( n518 , n30 );
buf ( n519 , n86 );
buf ( n520 , n186 );
buf ( n521 , n155 );
buf ( n522 , n56 );
buf ( n523 , n28 );
buf ( n524 , n85 );
buf ( n525 , n93 );
buf ( n526 , n58 );
buf ( n527 , n102 );
buf ( n528 , n128 );
buf ( n529 , n119 );
buf ( n530 , n53 );
buf ( n531 , n142 );
buf ( n532 , n96 );
buf ( n533 , n160 );
buf ( n534 , n174 );
buf ( n535 , n61 );
buf ( n536 , n65 );
buf ( n537 , n13 );
buf ( n538 , n8 );
buf ( n539 , n36 );
buf ( n540 , n11 );
buf ( n541 , n39 );
buf ( n542 , n177 );
buf ( n543 , n105 );
buf ( n544 , n139 );
buf ( n545 , n12 );
buf ( n546 , n99 );
buf ( n547 , n47 );
buf ( n548 , n79 );
buf ( n549 , n16 );
buf ( n550 , n87 );
buf ( n551 , n162 );
buf ( n552 , n110 );
buf ( n553 , n23 );
buf ( n554 , n187 );
buf ( n555 , n120 );
buf ( n556 , n32 );
buf ( n557 , n158 );
buf ( n558 , n176 );
buf ( n559 , n149 );
buf ( n560 , n148 );
buf ( n561 , n29 );
buf ( n562 , n97 );
buf ( n563 , n144 );
buf ( n564 , n27 );
buf ( n565 , n145 );
buf ( n566 , n108 );
buf ( n567 , n72 );
buf ( n568 , n90 );
buf ( n569 , n3 );
buf ( n570 , n133 );
buf ( n571 , n14 );
buf ( n572 , n6 );
buf ( n573 , n183 );
buf ( n574 , n81 );
buf ( n575 , n112 );
buf ( n576 , n5 );
buf ( n577 , n80 );
buf ( n578 , n17 );
buf ( n579 , n74 );
buf ( n580 , n37 );
buf ( n581 , n91 );
buf ( n582 , n151 );
buf ( n583 , n101 );
buf ( n584 , n189 );
buf ( n585 , n185 );
buf ( n586 , n42 );
buf ( n587 , n49 );
buf ( n588 , n18 );
buf ( n589 , n64 );
buf ( n590 , n48 );
buf ( n591 , n143 );
buf ( n592 , n76 );
buf ( n593 , n20 );
buf ( n594 , n190 );
buf ( n595 , n179 );
buf ( n596 , n35 );
buf ( n597 , n170 );
buf ( n598 , n406 );
buf ( n599 , n407 );
not ( n600 , n599 );
buf ( n601 , n408 );
and ( n602 , n600 , n601 );
not ( n603 , n602 );
buf ( n604 , n409 );
not ( n605 , n604 );
buf ( n606 , n410 );
not ( n607 , n606 );
buf ( n608 , n411 );
not ( n609 , n608 );
buf ( n610 , n412 );
not ( n611 , n610 );
buf ( n612 , n413 );
not ( n613 , n612 );
buf ( n614 , n414 );
not ( n615 , n614 );
buf ( n616 , n415 );
not ( n617 , n616 );
and ( n618 , n615 , n617 );
and ( n619 , n613 , n618 );
buf ( n620 , n416 );
not ( n621 , n620 );
buf ( n622 , n417 );
not ( n623 , n622 );
and ( n624 , n621 , n623 );
buf ( n625 , n418 );
not ( n626 , n625 );
buf ( n627 , n419 );
not ( n628 , n627 );
and ( n629 , n626 , n628 );
and ( n630 , n624 , n629 );
and ( n631 , n619 , n630 );
buf ( n632 , n420 );
not ( n633 , n632 );
buf ( n634 , n421 );
not ( n635 , n634 );
and ( n636 , n633 , n635 );
buf ( n637 , n422 );
not ( n638 , n637 );
buf ( n639 , n423 );
not ( n640 , n639 );
and ( n641 , n638 , n640 );
and ( n642 , n636 , n641 );
buf ( n643 , n424 );
not ( n644 , n643 );
buf ( n645 , n425 );
not ( n646 , n645 );
buf ( n647 , n426 );
not ( n648 , n647 );
buf ( n649 , n427 );
not ( n650 , n649 );
and ( n651 , n648 , n650 );
and ( n652 , n646 , n651 );
and ( n653 , n644 , n652 );
and ( n654 , n642 , n653 );
and ( n655 , n631 , n654 );
and ( n656 , n611 , n655 );
and ( n657 , n609 , n656 );
and ( n658 , n607 , n657 );
and ( n659 , n605 , n658 );
xor ( n660 , n601 , n659 );
not ( n661 , n660 );
and ( n662 , n599 , n661 );
not ( n663 , n662 );
and ( n664 , n603 , n663 );
buf ( n665 , n428 );
and ( n666 , n600 , n665 );
not ( n667 , n666 );
not ( n668 , n601 );
and ( n669 , n668 , n659 );
xor ( n670 , n665 , n669 );
not ( n671 , n670 );
and ( n672 , n599 , n671 );
not ( n673 , n672 );
and ( n674 , n667 , n673 );
and ( n675 , n664 , n674 );
not ( n676 , n675 );
not ( n677 , n674 );
buf ( n678 , n429 );
and ( n679 , n600 , n678 );
not ( n680 , n679 );
buf ( n681 , n430 );
not ( n682 , n681 );
not ( n683 , n665 );
and ( n684 , n683 , n669 );
and ( n685 , n682 , n684 );
xor ( n686 , n678 , n685 );
not ( n687 , n686 );
and ( n688 , n599 , n687 );
not ( n689 , n688 );
and ( n690 , n680 , n689 );
and ( n691 , n677 , n690 );
not ( n692 , n691 );
and ( n693 , n600 , n681 );
not ( n694 , n693 );
xor ( n695 , n681 , n684 );
not ( n696 , n695 );
and ( n697 , n599 , n696 );
not ( n698 , n697 );
and ( n699 , n694 , n698 );
not ( n700 , n699 );
not ( n701 , n690 );
and ( n702 , n700 , n701 );
not ( n703 , n702 );
and ( n704 , n699 , n690 );
not ( n705 , n704 );
and ( n706 , n703 , n705 );
not ( n707 , n706 );
and ( n708 , n676 , n692 , n707 );
not ( n709 , n708 );
buf ( n710 , n431 );
and ( n711 , n600 , n710 );
not ( n712 , n711 );
not ( n713 , n678 );
and ( n714 , n713 , n685 );
xor ( n715 , n710 , n714 );
not ( n716 , n715 );
and ( n717 , n599 , n716 );
not ( n718 , n717 );
and ( n719 , n712 , n718 );
buf ( n720 , n432 );
buf ( n721 , n433 );
and ( n722 , n600 , n721 );
not ( n723 , n722 );
buf ( n724 , n434 );
not ( n725 , n724 );
buf ( n726 , n435 );
not ( n727 , n726 );
not ( n728 , n710 );
and ( n729 , n728 , n714 );
and ( n730 , n727 , n729 );
and ( n731 , n725 , n730 );
xor ( n732 , n721 , n731 );
not ( n733 , n732 );
and ( n734 , n599 , n733 );
not ( n735 , n734 );
and ( n736 , n723 , n735 );
not ( n737 , n736 );
and ( n738 , n600 , n726 );
not ( n739 , n738 );
xor ( n740 , n726 , n729 );
not ( n741 , n740 );
and ( n742 , n599 , n741 );
not ( n743 , n742 );
and ( n744 , n739 , n743 );
not ( n745 , n744 );
and ( n746 , n600 , n724 );
not ( n747 , n746 );
xor ( n748 , n724 , n730 );
not ( n749 , n748 );
and ( n750 , n599 , n749 );
not ( n751 , n750 );
and ( n752 , n747 , n751 );
not ( n753 , n752 );
and ( n754 , n745 , n753 );
and ( n755 , n737 , n754 );
not ( n756 , n755 );
and ( n757 , n720 , n756 );
and ( n758 , n719 , n757 );
buf ( n759 , n436 );
not ( n760 , n759 );
buf ( n761 , n437 );
and ( n762 , n761 , n744 );
and ( n763 , n752 , n762 );
not ( n764 , n763 );
and ( n765 , n760 , n764 );
not ( n766 , n765 );
and ( n767 , n737 , n766 );
not ( n768 , n767 );
not ( n769 , n761 );
and ( n770 , n769 , n752 );
not ( n771 , n770 );
and ( n772 , n737 , n771 );
not ( n773 , n772 );
and ( n774 , n745 , n773 );
not ( n775 , n774 );
and ( n776 , n768 , n775 );
not ( n777 , n776 );
and ( n778 , n753 , n736 );
not ( n779 , n778 );
buf ( n780 , n438 );
not ( n781 , n780 );
and ( n782 , n769 , n745 );
not ( n783 , n782 );
not ( n784 , n762 );
and ( n785 , n783 , n784 );
not ( n786 , n785 );
and ( n787 , n752 , n786 );
not ( n788 , n787 );
and ( n789 , n781 , n788 );
not ( n790 , n789 );
and ( n791 , n737 , n790 );
not ( n792 , n791 );
and ( n793 , n779 , n792 );
and ( n794 , n709 , n758 , n777 , n793 );
not ( n795 , n794 );
and ( n796 , n598 , n795 );
not ( n797 , n796 );
buf ( n798 , n439 );
and ( n799 , n600 , n798 );
not ( n800 , n799 );
buf ( n801 , n440 );
not ( n802 , n801 );
not ( n803 , n721 );
and ( n804 , n803 , n731 );
and ( n805 , n802 , n804 );
xor ( n806 , n798 , n805 );
not ( n807 , n806 );
and ( n808 , n599 , n807 );
not ( n809 , n808 );
and ( n810 , n800 , n809 );
not ( n811 , n810 );
buf ( n812 , n441 );
buf ( n813 , n442 );
and ( n814 , n600 , n813 );
not ( n815 , n814 );
not ( n816 , n798 );
and ( n817 , n816 , n805 );
xor ( n818 , n813 , n817 );
not ( n819 , n818 );
and ( n820 , n599 , n819 );
not ( n821 , n820 );
and ( n822 , n815 , n821 );
not ( n823 , n822 );
buf ( n824 , n443 );
and ( n825 , n600 , n824 );
not ( n826 , n825 );
not ( n827 , n813 );
and ( n828 , n827 , n817 );
xor ( n829 , n824 , n828 );
not ( n830 , n829 );
and ( n831 , n599 , n830 );
not ( n832 , n831 );
and ( n833 , n826 , n832 );
and ( n834 , n823 , n833 );
and ( n835 , n812 , n834 );
not ( n836 , n835 );
buf ( n837 , n444 );
and ( n838 , n822 , n833 );
and ( n839 , n837 , n838 );
not ( n840 , n839 );
buf ( n841 , n445 );
not ( n842 , n833 );
and ( n843 , n823 , n842 );
and ( n844 , n841 , n843 );
not ( n845 , n844 );
buf ( n846 , n446 );
and ( n847 , n822 , n842 );
and ( n848 , n846 , n847 );
not ( n849 , n848 );
and ( n850 , n836 , n840 , n845 , n849 );
buf ( n851 , n447 );
and ( n852 , n851 , n834 );
not ( n853 , n852 );
buf ( n854 , n448 );
and ( n855 , n854 , n838 );
not ( n856 , n855 );
buf ( n857 , n449 );
and ( n858 , n857 , n843 );
not ( n859 , n858 );
buf ( n860 , n450 );
and ( n861 , n860 , n847 );
not ( n862 , n861 );
and ( n863 , n853 , n856 , n859 , n862 );
not ( n864 , n863 );
buf ( n865 , n451 );
and ( n866 , n865 , n838 );
not ( n867 , n866 );
buf ( n868 , n452 );
and ( n869 , n868 , n843 );
not ( n870 , n869 );
and ( n871 , n867 , n870 );
buf ( n872 , n453 );
and ( n873 , n872 , n847 );
not ( n874 , n873 );
buf ( n875 , n454 );
and ( n876 , n875 , n834 );
not ( n877 , n876 );
and ( n878 , n874 , n877 );
and ( n879 , n871 , n878 );
not ( n880 , n879 );
and ( n881 , n864 , n880 );
buf ( n882 , n455 );
and ( n883 , n882 , n834 );
not ( n884 , n883 );
buf ( n885 , n456 );
and ( n886 , n885 , n838 );
not ( n887 , n886 );
buf ( n888 , n457 );
and ( n889 , n888 , n843 );
not ( n890 , n889 );
buf ( n891 , n458 );
and ( n892 , n891 , n847 );
not ( n893 , n892 );
and ( n894 , n884 , n887 , n890 , n893 );
not ( n895 , n894 );
buf ( n896 , n459 );
and ( n897 , n896 , n834 );
not ( n898 , n897 );
buf ( n899 , n460 );
and ( n900 , n899 , n838 );
not ( n901 , n900 );
buf ( n902 , n461 );
and ( n903 , n902 , n843 );
not ( n904 , n903 );
buf ( n905 , n462 );
and ( n906 , n905 , n847 );
not ( n907 , n906 );
and ( n908 , n898 , n901 , n904 , n907 );
not ( n909 , n908 );
buf ( n910 , n463 );
and ( n911 , n910 , n834 );
not ( n912 , n911 );
buf ( n913 , n464 );
and ( n914 , n913 , n838 );
not ( n915 , n914 );
buf ( n916 , n465 );
and ( n917 , n916 , n843 );
not ( n918 , n917 );
buf ( n919 , n466 );
and ( n920 , n919 , n847 );
not ( n921 , n920 );
and ( n922 , n912 , n915 , n918 , n921 );
not ( n923 , n922 );
buf ( n924 , n467 );
and ( n925 , n924 , n834 );
not ( n926 , n925 );
buf ( n927 , n468 );
and ( n928 , n927 , n838 );
not ( n929 , n928 );
buf ( n930 , n469 );
and ( n931 , n930 , n843 );
not ( n932 , n931 );
buf ( n933 , n470 );
and ( n934 , n933 , n847 );
not ( n935 , n934 );
and ( n936 , n926 , n929 , n932 , n935 );
not ( n937 , n936 );
and ( n938 , n923 , n937 );
and ( n939 , n895 , n909 , n938 );
buf ( n940 , n471 );
and ( n941 , n940 , n834 );
not ( n942 , n941 );
buf ( n943 , n472 );
and ( n944 , n943 , n838 );
not ( n945 , n944 );
buf ( n946 , n473 );
and ( n947 , n946 , n843 );
not ( n948 , n947 );
buf ( n949 , n474 );
and ( n950 , n949 , n847 );
not ( n951 , n950 );
and ( n952 , n942 , n945 , n948 , n951 );
not ( n953 , n952 );
buf ( n954 , n475 );
and ( n955 , n954 , n834 );
not ( n956 , n955 );
buf ( n957 , n476 );
and ( n958 , n957 , n838 );
not ( n959 , n958 );
buf ( n960 , n477 );
and ( n961 , n960 , n843 );
not ( n962 , n961 );
buf ( n963 , n478 );
and ( n964 , n963 , n847 );
not ( n965 , n964 );
and ( n966 , n956 , n959 , n962 , n965 );
not ( n967 , n966 );
and ( n968 , n953 , n967 );
buf ( n969 , n479 );
and ( n970 , n969 , n834 );
not ( n971 , n970 );
buf ( n972 , n480 );
and ( n973 , n972 , n838 );
not ( n974 , n973 );
buf ( n975 , n481 );
and ( n976 , n975 , n843 );
not ( n977 , n976 );
buf ( n978 , n482 );
and ( n979 , n978 , n847 );
not ( n980 , n979 );
and ( n981 , n971 , n974 , n977 , n980 );
not ( n982 , n981 );
buf ( n983 , n483 );
and ( n984 , n983 , n834 );
not ( n985 , n984 );
buf ( n986 , n484 );
and ( n987 , n986 , n838 );
not ( n988 , n987 );
buf ( n989 , n485 );
and ( n990 , n989 , n843 );
not ( n991 , n990 );
buf ( n992 , n486 );
and ( n993 , n992 , n847 );
not ( n994 , n993 );
and ( n995 , n985 , n988 , n991 , n994 );
not ( n996 , n995 );
buf ( n997 , n487 );
and ( n998 , n997 , n834 );
not ( n999 , n998 );
buf ( n1000 , n488 );
and ( n1001 , n1000 , n838 );
not ( n1002 , n1001 );
buf ( n1003 , n489 );
and ( n1004 , n1003 , n843 );
not ( n1005 , n1004 );
buf ( n1006 , n490 );
and ( n1007 , n1006 , n847 );
not ( n1008 , n1007 );
and ( n1009 , n999 , n1002 , n1005 , n1008 );
not ( n1010 , n1009 );
and ( n1011 , n843 , n982 , n996 , n1010 );
and ( n1012 , n968 , n1011 );
and ( n1013 , n881 , n939 , n1012 );
and ( n1014 , n850 , n1013 );
not ( n1015 , n1014 );
not ( n1016 , n850 );
not ( n1017 , n1013 );
and ( n1018 , n1016 , n1017 );
not ( n1019 , n1018 );
and ( n1020 , n1015 , n1019 );
not ( n1021 , n1020 );
and ( n1022 , n811 , n1021 );
not ( n1023 , n1022 );
buf ( n1024 , n491 );
and ( n1025 , n1024 , n834 );
not ( n1026 , n1025 );
buf ( n1027 , n492 );
and ( n1028 , n1027 , n838 );
not ( n1029 , n1028 );
buf ( n1030 , n493 );
and ( n1031 , n1030 , n843 );
not ( n1032 , n1031 );
buf ( n1033 , n494 );
and ( n1034 , n1033 , n847 );
not ( n1035 , n1034 );
and ( n1036 , n1026 , n1029 , n1032 , n1035 );
and ( n1037 , n895 , n909 );
and ( n1038 , n598 , n834 );
not ( n1039 , n1038 );
buf ( n1040 , n495 );
and ( n1041 , n1040 , n838 );
not ( n1042 , n1041 );
buf ( n1043 , n496 );
and ( n1044 , n1043 , n843 );
not ( n1045 , n1044 );
buf ( n1046 , n497 );
and ( n1047 , n1046 , n847 );
not ( n1048 , n1047 );
and ( n1049 , n1039 , n1042 , n1045 , n1048 );
not ( n1050 , n1049 );
and ( n1051 , n1016 , n1050 );
and ( n1052 , n1037 , n1051 );
and ( n1053 , n923 , n937 , n953 , n967 );
and ( n1054 , n1053 , n881 );
and ( n1055 , n1011 , n1052 , n1054 );
xor ( n1056 , n1036 , n1055 );
buf ( n1057 , n498 );
and ( n1058 , n1057 , n834 );
not ( n1059 , n1058 );
buf ( n1060 , n499 );
and ( n1061 , n1060 , n838 );
not ( n1062 , n1061 );
buf ( n1063 , n500 );
and ( n1064 , n1063 , n847 );
not ( n1065 , n1064 );
and ( n1066 , n1059 , n1062 , n1065 );
not ( n1067 , n1066 );
buf ( n1068 , n501 );
and ( n1069 , n1068 , n838 );
not ( n1070 , n1069 );
buf ( n1071 , n502 );
and ( n1072 , n1071 , n834 );
not ( n1073 , n1072 );
and ( n1074 , n1070 , n1073 );
buf ( n1075 , n503 );
and ( n1076 , n1075 , n843 );
not ( n1077 , n1076 );
buf ( n1078 , n504 );
and ( n1079 , n1078 , n847 );
not ( n1080 , n1079 );
and ( n1081 , n1077 , n1080 );
and ( n1082 , n1074 , n1081 );
not ( n1083 , n1082 );
and ( n1084 , n1067 , n1083 );
and ( n1085 , n1016 , n881 );
and ( n1086 , n939 , n1012 );
and ( n1087 , n1085 , n1086 );
xor ( n1088 , n1049 , n1087 );
not ( n1089 , n1088 );
and ( n1090 , n1021 , n1089 );
and ( n1091 , n864 , n939 , n1012 );
xor ( n1092 , n879 , n1091 );
not ( n1093 , n1092 );
xor ( n1094 , n936 , n1012 );
not ( n1095 , n1094 );
and ( n1096 , n1004 , n996 , n968 );
and ( n1097 , n981 , n1096 );
not ( n1098 , n1097 );
not ( n1099 , n1096 );
and ( n1100 , n982 , n1099 );
not ( n1101 , n1100 );
and ( n1102 , n1098 , n1101 );
not ( n1103 , n1102 );
not ( n1104 , n843 );
and ( n1105 , n1104 , n1009 );
not ( n1106 , n1105 );
and ( n1107 , n1005 , n1106 );
buf ( n1108 , n505 );
and ( n1109 , n1108 , n834 );
not ( n1110 , n1109 );
buf ( n1111 , n506 );
and ( n1112 , n1111 , n838 );
not ( n1113 , n1112 );
buf ( n1114 , n507 );
and ( n1115 , n1114 , n843 );
not ( n1116 , n1115 );
buf ( n1117 , n508 );
and ( n1118 , n1117 , n847 );
not ( n1119 , n1118 );
and ( n1120 , n1110 , n1113 , n1116 , n1119 );
not ( n1121 , n1120 );
buf ( n1122 , n509 );
and ( n1123 , n1122 , n838 );
not ( n1124 , n1123 );
buf ( n1125 , n510 );
and ( n1126 , n1125 , n834 );
not ( n1127 , n1126 );
and ( n1128 , n1124 , n1127 );
buf ( n1129 , n511 );
and ( n1130 , n1129 , n843 );
not ( n1131 , n1130 );
buf ( n1132 , n512 );
and ( n1133 , n1132 , n847 );
not ( n1134 , n1133 );
and ( n1135 , n1131 , n1134 );
and ( n1136 , n1128 , n1135 );
not ( n1137 , n1136 );
and ( n1138 , n1121 , n1137 );
and ( n1139 , n1004 , n966 );
not ( n1140 , n1139 );
and ( n1141 , n1005 , n967 );
not ( n1142 , n1141 );
and ( n1143 , n1140 , n1142 );
not ( n1144 , n1143 );
and ( n1145 , n1107 , n1138 , n1144 );
and ( n1146 , n1004 , n968 );
and ( n1147 , n995 , n1146 );
not ( n1148 , n1147 );
not ( n1149 , n1146 );
and ( n1150 , n996 , n1149 );
not ( n1151 , n1150 );
and ( n1152 , n1148 , n1151 );
not ( n1153 , n1152 );
and ( n1154 , n1004 , n967 );
not ( n1155 , n1154 );
and ( n1156 , n952 , n1155 );
not ( n1157 , n1156 );
and ( n1158 , n1149 , n1157 );
and ( n1159 , n1153 , n1158 );
and ( n1160 , n1145 , n1159 );
and ( n1161 , n1095 , n1103 , n1160 );
and ( n1162 , n909 , n938 , n1012 );
and ( n1163 , n894 , n1162 );
not ( n1164 , n1163 );
not ( n1165 , n1162 );
and ( n1166 , n895 , n1165 );
not ( n1167 , n1166 );
and ( n1168 , n1164 , n1167 );
not ( n1169 , n1168 );
and ( n1170 , n863 , n1086 );
not ( n1171 , n1170 );
not ( n1172 , n1086 );
and ( n1173 , n864 , n1172 );
not ( n1174 , n1173 );
and ( n1175 , n1171 , n1174 );
not ( n1176 , n1175 );
and ( n1177 , n1169 , n1176 );
and ( n1178 , n938 , n1012 );
and ( n1179 , n908 , n1178 );
not ( n1180 , n1179 );
not ( n1181 , n1178 );
and ( n1182 , n909 , n1181 );
not ( n1183 , n1182 );
and ( n1184 , n1180 , n1183 );
not ( n1185 , n1184 );
and ( n1186 , n937 , n1012 );
and ( n1187 , n922 , n1186 );
not ( n1188 , n1187 );
not ( n1189 , n1186 );
and ( n1190 , n923 , n1189 );
not ( n1191 , n1190 );
and ( n1192 , n1188 , n1191 );
not ( n1193 , n1192 );
and ( n1194 , n1185 , n1193 );
and ( n1195 , n1177 , n1194 );
and ( n1196 , n1093 , n1161 , n1195 );
and ( n1197 , n1090 , n1196 );
and ( n1198 , n1084 , n1197 );
and ( n1199 , n1056 , n1198 );
not ( n1200 , n1199 );
not ( n1201 , n1056 );
not ( n1202 , n1198 );
and ( n1203 , n1201 , n1202 );
not ( n1204 , n1203 );
and ( n1205 , n1200 , n1204 );
not ( n1206 , n1205 );
and ( n1207 , n810 , n1206 );
not ( n1208 , n1207 );
and ( n1209 , n1023 , n1208 );
not ( n1210 , n1209 );
and ( n1211 , n702 , n1210 );
not ( n1212 , n1211 );
and ( n1213 , n699 , n691 );
buf ( n1214 , n513 );
and ( n1215 , n600 , n801 );
not ( n1216 , n1215 );
xor ( n1217 , n801 , n804 );
not ( n1218 , n1217 );
and ( n1219 , n599 , n1218 );
not ( n1220 , n1219 );
and ( n1221 , n1216 , n1220 );
not ( n1222 , n1221 );
and ( n1223 , n1222 , n810 );
not ( n1224 , n1223 );
and ( n1225 , n1221 , n811 );
not ( n1226 , n1225 );
and ( n1227 , n1224 , n1226 );
and ( n1228 , n1221 , n1227 );
not ( n1229 , n1228 );
and ( n1230 , n1214 , n1229 );
not ( n1231 , n1230 );
and ( n1232 , n600 , n610 );
not ( n1233 , n1232 );
xor ( n1234 , n610 , n655 );
not ( n1235 , n1234 );
and ( n1236 , n599 , n1235 );
not ( n1237 , n1236 );
and ( n1238 , n1233 , n1237 );
not ( n1239 , n1238 );
and ( n1240 , n1239 , n1228 );
not ( n1241 , n1240 );
and ( n1242 , n1231 , n1241 );
not ( n1243 , n1242 );
and ( n1244 , n1213 , n1243 );
not ( n1245 , n1244 );
and ( n1246 , n664 , n674 , n699 , n690 );
buf ( n1247 , n514 );
and ( n1248 , n1247 , n1229 );
not ( n1249 , n1248 );
and ( n1250 , n600 , n612 );
not ( n1251 , n1250 );
and ( n1252 , n630 , n654 );
and ( n1253 , n617 , n1252 );
and ( n1254 , n615 , n1253 );
xor ( n1255 , n612 , n1254 );
not ( n1256 , n1255 );
and ( n1257 , n599 , n1256 );
not ( n1258 , n1257 );
and ( n1259 , n1251 , n1258 );
not ( n1260 , n1259 );
and ( n1261 , n1260 , n1228 );
not ( n1262 , n1261 );
and ( n1263 , n1249 , n1262 );
buf ( n1264 , n515 );
and ( n1265 , n1264 , n1229 );
not ( n1266 , n1265 );
and ( n1267 , n600 , n620 );
not ( n1268 , n1267 );
and ( n1269 , n623 , n629 );
and ( n1270 , n1269 , n654 );
xor ( n1271 , n620 , n1270 );
not ( n1272 , n1271 );
and ( n1273 , n599 , n1272 );
not ( n1274 , n1273 );
and ( n1275 , n1268 , n1274 );
not ( n1276 , n1275 );
and ( n1277 , n1276 , n1228 );
not ( n1278 , n1277 );
and ( n1279 , n1266 , n1278 );
buf ( n1280 , n516 );
and ( n1281 , n1280 , n1229 );
not ( n1282 , n1281 );
and ( n1283 , n600 , n622 );
not ( n1284 , n1283 );
and ( n1285 , n629 , n654 );
xor ( n1286 , n622 , n1285 );
not ( n1287 , n1286 );
and ( n1288 , n599 , n1287 );
not ( n1289 , n1288 );
and ( n1290 , n1284 , n1289 );
not ( n1291 , n1290 );
and ( n1292 , n1291 , n1228 );
not ( n1293 , n1292 );
and ( n1294 , n1282 , n1293 );
buf ( n1295 , n517 );
and ( n1296 , n1295 , n1229 );
not ( n1297 , n1296 );
and ( n1298 , n600 , n627 );
not ( n1299 , n1298 );
xor ( n1300 , n627 , n654 );
not ( n1301 , n1300 );
and ( n1302 , n599 , n1301 );
not ( n1303 , n1302 );
and ( n1304 , n1299 , n1303 );
not ( n1305 , n1304 );
and ( n1306 , n1305 , n1228 );
not ( n1307 , n1306 );
and ( n1308 , n1297 , n1307 );
buf ( n1309 , n518 );
and ( n1310 , n1309 , n1229 );
not ( n1311 , n1310 );
and ( n1312 , n600 , n625 );
not ( n1313 , n1312 );
and ( n1314 , n628 , n654 );
xor ( n1315 , n625 , n1314 );
not ( n1316 , n1315 );
and ( n1317 , n599 , n1316 );
not ( n1318 , n1317 );
and ( n1319 , n1313 , n1318 );
not ( n1320 , n1319 );
and ( n1321 , n1320 , n1228 );
not ( n1322 , n1321 );
and ( n1323 , n1311 , n1322 );
and ( n1324 , n1308 , n1323 );
and ( n1325 , n1279 , n1294 , n1324 );
buf ( n1326 , n519 );
and ( n1327 , n1326 , n1229 );
not ( n1328 , n1327 );
and ( n1329 , n600 , n616 );
not ( n1330 , n1329 );
xor ( n1331 , n616 , n1252 );
not ( n1332 , n1331 );
and ( n1333 , n599 , n1332 );
not ( n1334 , n1333 );
and ( n1335 , n1330 , n1334 );
not ( n1336 , n1335 );
and ( n1337 , n1336 , n1228 );
not ( n1338 , n1337 );
and ( n1339 , n1328 , n1338 );
buf ( n1340 , n520 );
and ( n1341 , n1340 , n1229 );
not ( n1342 , n1341 );
and ( n1343 , n600 , n614 );
not ( n1344 , n1343 );
xor ( n1345 , n614 , n1253 );
not ( n1346 , n1345 );
and ( n1347 , n599 , n1346 );
not ( n1348 , n1347 );
and ( n1349 , n1344 , n1348 );
not ( n1350 , n1349 );
and ( n1351 , n1350 , n1228 );
not ( n1352 , n1351 );
and ( n1353 , n1342 , n1352 );
and ( n1354 , n1339 , n1353 );
and ( n1355 , n1263 , n1325 , n1354 );
buf ( n1356 , n521 );
and ( n1357 , n1356 , n1229 );
not ( n1358 , n1357 );
and ( n1359 , n600 , n643 );
not ( n1360 , n1359 );
xor ( n1361 , n643 , n652 );
not ( n1362 , n1361 );
and ( n1363 , n599 , n1362 );
not ( n1364 , n1363 );
and ( n1365 , n1360 , n1364 );
not ( n1366 , n1365 );
and ( n1367 , n1366 , n1228 );
not ( n1368 , n1367 );
and ( n1369 , n1358 , n1368 );
buf ( n1370 , n522 );
and ( n1371 , n1370 , n1229 );
not ( n1372 , n1371 );
and ( n1373 , n600 , n645 );
not ( n1374 , n1373 );
xor ( n1375 , n645 , n651 );
not ( n1376 , n1375 );
and ( n1377 , n599 , n1376 );
not ( n1378 , n1377 );
and ( n1379 , n1374 , n1378 );
not ( n1380 , n1379 );
and ( n1381 , n1380 , n1228 );
not ( n1382 , n1381 );
and ( n1383 , n1372 , n1382 );
and ( n1384 , n1369 , n1383 );
buf ( n1385 , n523 );
and ( n1386 , n1385 , n1229 );
not ( n1387 , n1386 );
and ( n1388 , n649 , n1228 );
not ( n1389 , n1388 );
and ( n1390 , n1387 , n1389 );
buf ( n1391 , n524 );
and ( n1392 , n1391 , n1229 );
not ( n1393 , n1392 );
and ( n1394 , n600 , n647 );
not ( n1395 , n1394 );
xor ( n1396 , n647 , n649 );
and ( n1397 , n599 , n1396 );
not ( n1398 , n1397 );
and ( n1399 , n1395 , n1398 );
not ( n1400 , n1399 );
and ( n1401 , n1400 , n1228 );
not ( n1402 , n1401 );
and ( n1403 , n1393 , n1402 );
and ( n1404 , n1390 , n1403 );
and ( n1405 , n1384 , n1404 );
buf ( n1406 , n525 );
and ( n1407 , n1406 , n1229 );
not ( n1408 , n1407 );
and ( n1409 , n600 , n632 );
not ( n1410 , n1409 );
and ( n1411 , n640 , n653 );
and ( n1412 , n638 , n1411 );
and ( n1413 , n635 , n1412 );
xor ( n1414 , n632 , n1413 );
not ( n1415 , n1414 );
and ( n1416 , n599 , n1415 );
not ( n1417 , n1416 );
and ( n1418 , n1410 , n1417 );
not ( n1419 , n1418 );
and ( n1420 , n1419 , n1228 );
not ( n1421 , n1420 );
and ( n1422 , n1408 , n1421 );
buf ( n1423 , n526 );
and ( n1424 , n1423 , n1229 );
not ( n1425 , n1424 );
and ( n1426 , n600 , n637 );
not ( n1427 , n1426 );
xor ( n1428 , n637 , n1411 );
not ( n1429 , n1428 );
and ( n1430 , n599 , n1429 );
not ( n1431 , n1430 );
and ( n1432 , n1427 , n1431 );
not ( n1433 , n1432 );
and ( n1434 , n1433 , n1228 );
not ( n1435 , n1434 );
and ( n1436 , n1425 , n1435 );
and ( n1437 , n1422 , n1436 );
buf ( n1438 , n527 );
and ( n1439 , n1438 , n1229 );
not ( n1440 , n1439 );
and ( n1441 , n600 , n634 );
not ( n1442 , n1441 );
xor ( n1443 , n634 , n1412 );
not ( n1444 , n1443 );
and ( n1445 , n599 , n1444 );
not ( n1446 , n1445 );
and ( n1447 , n1442 , n1446 );
not ( n1448 , n1447 );
and ( n1449 , n1448 , n1228 );
not ( n1450 , n1449 );
and ( n1451 , n1440 , n1450 );
buf ( n1452 , n528 );
and ( n1453 , n1452 , n1229 );
not ( n1454 , n1453 );
and ( n1455 , n600 , n639 );
not ( n1456 , n1455 );
xor ( n1457 , n639 , n653 );
not ( n1458 , n1457 );
and ( n1459 , n599 , n1458 );
not ( n1460 , n1459 );
and ( n1461 , n1456 , n1460 );
not ( n1462 , n1461 );
and ( n1463 , n1462 , n1228 );
not ( n1464 , n1463 );
and ( n1465 , n1454 , n1464 );
and ( n1466 , n1451 , n1465 );
and ( n1467 , n1437 , n1466 );
and ( n1468 , n1405 , n1467 );
and ( n1469 , n1355 , n1468 );
and ( n1470 , n1243 , n1469 );
not ( n1471 , n1470 );
not ( n1472 , n1469 );
and ( n1473 , n1242 , n1472 );
not ( n1474 , n1473 );
and ( n1475 , n1471 , n1474 );
not ( n1476 , n1475 );
and ( n1477 , n1246 , n1476 );
not ( n1478 , n1477 );
and ( n1479 , n1245 , n1478 );
not ( n1480 , n664 );
and ( n1481 , n1480 , n701 );
not ( n1482 , n1481 );
and ( n1483 , n1482 , n692 );
and ( n1484 , n1483 , n706 );
not ( n1485 , n1263 );
and ( n1486 , n1485 , n1016 );
and ( n1487 , n1242 , n1050 );
not ( n1488 , n1487 );
and ( n1489 , n1243 , n1049 );
not ( n1490 , n1489 );
and ( n1491 , n1488 , n1490 );
not ( n1492 , n1491 );
and ( n1493 , n1486 , n1492 );
not ( n1494 , n1493 );
not ( n1495 , n1486 );
and ( n1496 , n1495 , n1491 );
not ( n1497 , n1496 );
and ( n1498 , n1494 , n1497 );
not ( n1499 , n1353 );
and ( n1500 , n1499 , n880 );
not ( n1501 , n1500 );
and ( n1502 , n1263 , n1016 );
not ( n1503 , n1502 );
and ( n1504 , n1485 , n850 );
not ( n1505 , n1504 );
and ( n1506 , n1503 , n1505 );
and ( n1507 , n1501 , n1506 );
not ( n1508 , n1507 );
not ( n1509 , n1279 );
and ( n1510 , n1509 , n895 );
not ( n1511 , n1510 );
not ( n1512 , n1339 );
and ( n1513 , n1512 , n863 );
not ( n1514 , n1513 );
and ( n1515 , n1339 , n864 );
not ( n1516 , n1515 );
and ( n1517 , n1514 , n1516 );
and ( n1518 , n1511 , n1517 );
not ( n1519 , n1518 );
and ( n1520 , n1512 , n864 );
not ( n1521 , n1520 );
and ( n1522 , n1353 , n879 );
not ( n1523 , n1522 );
and ( n1524 , n1501 , n1523 );
not ( n1525 , n1524 );
and ( n1526 , n1521 , n1525 );
not ( n1527 , n1526 );
and ( n1528 , n1519 , n1527 );
and ( n1529 , n1508 , n1528 );
not ( n1530 , n1294 );
and ( n1531 , n1530 , n909 );
and ( n1532 , n1509 , n894 );
not ( n1533 , n1532 );
and ( n1534 , n1279 , n895 );
not ( n1535 , n1534 );
and ( n1536 , n1533 , n1535 );
not ( n1537 , n1536 );
and ( n1538 , n1531 , n1537 );
not ( n1539 , n1538 );
xor ( n1540 , n1294 , n908 );
not ( n1541 , n1540 );
not ( n1542 , n1323 );
and ( n1543 , n1542 , n923 );
not ( n1544 , n1543 );
and ( n1545 , n1541 , n1544 );
not ( n1546 , n1545 );
not ( n1547 , n1531 );
and ( n1548 , n1547 , n1536 );
not ( n1549 , n1548 );
and ( n1550 , n1546 , n1549 );
not ( n1551 , n1550 );
and ( n1552 , n1539 , n1551 );
not ( n1553 , n1552 );
and ( n1554 , n1540 , n1543 );
not ( n1555 , n1554 );
xor ( n1556 , n1323 , n922 );
not ( n1557 , n1308 );
and ( n1558 , n1557 , n937 );
and ( n1559 , n1556 , n1558 );
not ( n1560 , n1559 );
and ( n1561 , n1555 , n1539 , n1560 );
not ( n1562 , n1556 );
not ( n1563 , n1558 );
and ( n1564 , n1562 , n1563 );
not ( n1565 , n1564 );
not ( n1566 , n1422 );
and ( n1567 , n1566 , n982 );
and ( n1568 , n1557 , n936 );
not ( n1569 , n1568 );
and ( n1570 , n1308 , n937 );
not ( n1571 , n1570 );
and ( n1572 , n1569 , n1571 );
not ( n1573 , n1572 );
and ( n1574 , n1567 , n1573 );
and ( n1575 , n1565 , n1574 );
not ( n1576 , n1575 );
and ( n1577 , n1561 , n1576 );
not ( n1578 , n1577 );
and ( n1579 , n1553 , n1578 );
and ( n1580 , n1529 , n1579 );
not ( n1581 , n1580 );
not ( n1582 , n1506 );
and ( n1583 , n1500 , n1582 );
not ( n1584 , n1583 );
and ( n1585 , n1520 , n1524 );
not ( n1586 , n1585 );
not ( n1587 , n1517 );
and ( n1588 , n1510 , n1587 );
and ( n1589 , n1588 , n1527 );
not ( n1590 , n1589 );
and ( n1591 , n1586 , n1590 );
not ( n1592 , n1591 );
and ( n1593 , n1508 , n1592 );
not ( n1594 , n1593 );
and ( n1595 , n1584 , n1594 );
and ( n1596 , n1581 , n1595 );
not ( n1597 , n1567 );
and ( n1598 , n1597 , n1572 );
not ( n1599 , n1598 );
and ( n1600 , n1565 , n1599 );
and ( n1601 , n1550 , n1600 );
and ( n1602 , n1529 , n1601 );
not ( n1603 , n1451 );
and ( n1604 , n1603 , n996 );
and ( n1605 , n1422 , n981 );
not ( n1606 , n1605 );
and ( n1607 , n1597 , n1606 );
and ( n1608 , n1604 , n1607 );
not ( n1609 , n1608 );
not ( n1610 , n1604 );
not ( n1611 , n1607 );
and ( n1612 , n1610 , n1611 );
not ( n1613 , n1612 );
not ( n1614 , n1436 );
and ( n1615 , n1614 , n953 );
and ( n1616 , n1451 , n996 );
not ( n1617 , n1616 );
and ( n1618 , n1603 , n995 );
not ( n1619 , n1618 );
and ( n1620 , n1617 , n1619 );
not ( n1621 , n1620 );
and ( n1622 , n1615 , n1621 );
and ( n1623 , n1613 , n1622 );
not ( n1624 , n1623 );
and ( n1625 , n1609 , n1624 );
not ( n1626 , n1615 );
and ( n1627 , n1626 , n1620 );
not ( n1628 , n1627 );
and ( n1629 , n1613 , n1628 );
not ( n1630 , n1465 );
and ( n1631 , n1630 , n967 );
and ( n1632 , n1614 , n952 );
not ( n1633 , n1632 );
and ( n1634 , n1436 , n953 );
not ( n1635 , n1634 );
and ( n1636 , n1633 , n1635 );
not ( n1637 , n1636 );
and ( n1638 , n1631 , n1637 );
not ( n1639 , n1638 );
not ( n1640 , n1631 );
and ( n1641 , n1640 , n1636 );
not ( n1642 , n1641 );
and ( n1643 , n1465 , n967 );
not ( n1644 , n1643 );
and ( n1645 , n1630 , n966 );
not ( n1646 , n1645 );
and ( n1647 , n1644 , n1646 );
not ( n1648 , n1647 );
not ( n1649 , n1369 );
and ( n1650 , n1649 , n1107 );
not ( n1651 , n1650 );
and ( n1652 , n1005 , n1651 );
not ( n1653 , n1652 );
and ( n1654 , n1648 , n1653 );
and ( n1655 , n1642 , n1654 );
not ( n1656 , n1655 );
and ( n1657 , n1639 , n1656 );
not ( n1658 , n1657 );
and ( n1659 , n1629 , n1658 );
not ( n1660 , n1659 );
and ( n1661 , n1625 , n1660 );
and ( n1662 , n1647 , n1652 );
not ( n1663 , n1662 );
and ( n1664 , n1642 , n1663 );
and ( n1665 , n1629 , n1664 );
not ( n1666 , n1383 );
and ( n1667 , n1666 , n1137 );
xor ( n1668 , n1369 , n1107 );
not ( n1669 , n1668 );
and ( n1670 , n1667 , n1669 );
not ( n1671 , n1670 );
not ( n1672 , n1667 );
and ( n1673 , n1672 , n1668 );
not ( n1674 , n1673 );
not ( n1675 , n1403 );
and ( n1676 , n1675 , n1121 );
xor ( n1677 , n1383 , n1136 );
and ( n1678 , n1676 , n1677 );
and ( n1679 , n1674 , n1678 );
not ( n1680 , n1679 );
xor ( n1681 , n1403 , n1120 );
not ( n1682 , n1390 );
and ( n1683 , n1682 , n1083 );
and ( n1684 , n1681 , n1683 );
not ( n1685 , n1676 );
not ( n1686 , n1677 );
and ( n1687 , n1685 , n1686 );
not ( n1688 , n1687 );
and ( n1689 , n1684 , n1688 );
and ( n1690 , n1674 , n1689 );
not ( n1691 , n1690 );
and ( n1692 , n1671 , n1680 , n1691 );
not ( n1693 , n1692 );
and ( n1694 , n1665 , n1693 );
not ( n1695 , n1694 );
and ( n1696 , n1661 , n1695 );
not ( n1697 , n1696 );
and ( n1698 , n1602 , n1697 );
not ( n1699 , n1698 );
and ( n1700 , n1596 , n1699 );
and ( n1701 , n1498 , n1700 );
not ( n1702 , n1701 );
not ( n1703 , n1498 );
not ( n1704 , n1700 );
and ( n1705 , n1703 , n1704 );
not ( n1706 , n1705 );
and ( n1707 , n1702 , n1706 );
not ( n1708 , n1707 );
and ( n1709 , n1484 , n1708 );
not ( n1710 , n1709 );
and ( n1711 , n1479 , n1710 );
and ( n1712 , n691 , n705 );
not ( n1713 , n1712 );
and ( n1714 , n1482 , n1713 );
not ( n1715 , n1714 );
xor ( n1716 , n1502 , n1491 );
and ( n1717 , n1353 , n880 );
and ( n1718 , n1717 , n1506 );
not ( n1719 , n1718 );
not ( n1720 , n1717 );
and ( n1721 , n1720 , n1582 );
not ( n1722 , n1721 );
and ( n1723 , n1515 , n1525 );
not ( n1724 , n1723 );
and ( n1725 , n1516 , n1524 );
not ( n1726 , n1725 );
and ( n1727 , n1534 , n1517 );
and ( n1728 , n1726 , n1727 );
not ( n1729 , n1728 );
and ( n1730 , n1724 , n1729 );
not ( n1731 , n1730 );
and ( n1732 , n1722 , n1731 );
not ( n1733 , n1732 );
and ( n1734 , n1719 , n1733 );
and ( n1735 , n1535 , n1587 );
not ( n1736 , n1735 );
and ( n1737 , n1726 , n1736 );
and ( n1738 , n1722 , n1737 );
and ( n1739 , n1294 , n909 );
and ( n1740 , n1739 , n1536 );
not ( n1741 , n1740 );
not ( n1742 , n1739 );
and ( n1743 , n1742 , n1537 );
not ( n1744 , n1743 );
and ( n1745 , n1323 , n923 );
and ( n1746 , n1541 , n1745 );
and ( n1747 , n1744 , n1746 );
not ( n1748 , n1747 );
and ( n1749 , n1741 , n1748 );
not ( n1750 , n1745 );
and ( n1751 , n1540 , n1750 );
not ( n1752 , n1751 );
and ( n1753 , n1744 , n1752 );
and ( n1754 , n1562 , n1570 );
not ( n1755 , n1754 );
and ( n1756 , n1556 , n1571 );
not ( n1757 , n1756 );
and ( n1758 , n1422 , n982 );
and ( n1759 , n1758 , n1572 );
and ( n1760 , n1757 , n1759 );
not ( n1761 , n1760 );
and ( n1762 , n1755 , n1761 );
not ( n1763 , n1762 );
and ( n1764 , n1753 , n1763 );
not ( n1765 , n1764 );
and ( n1766 , n1749 , n1765 );
not ( n1767 , n1766 );
and ( n1768 , n1738 , n1767 );
not ( n1769 , n1768 );
and ( n1770 , n1734 , n1769 );
not ( n1771 , n1758 );
and ( n1772 , n1771 , n1573 );
not ( n1773 , n1772 );
and ( n1774 , n1744 , n1752 , n1757 , n1773 );
and ( n1775 , n1738 , n1774 );
and ( n1776 , n1616 , n1611 );
not ( n1777 , n1776 );
and ( n1778 , n1617 , n1607 );
not ( n1779 , n1778 );
and ( n1780 , n1634 , n1620 );
and ( n1781 , n1779 , n1780 );
not ( n1782 , n1781 );
and ( n1783 , n1777 , n1782 );
and ( n1784 , n1635 , n1621 );
not ( n1785 , n1784 );
and ( n1786 , n1779 , n1785 );
and ( n1787 , n1643 , n1636 );
not ( n1788 , n1787 );
and ( n1789 , n1644 , n1637 );
not ( n1790 , n1789 );
and ( n1791 , n1369 , n1106 );
not ( n1792 , n1791 );
and ( n1793 , n1005 , n1792 );
not ( n1794 , n1793 );
and ( n1795 , n1647 , n1794 );
and ( n1796 , n1790 , n1795 );
not ( n1797 , n1796 );
and ( n1798 , n1788 , n1797 );
not ( n1799 , n1798 );
and ( n1800 , n1786 , n1799 );
not ( n1801 , n1800 );
and ( n1802 , n1783 , n1801 );
and ( n1803 , n1648 , n1793 );
not ( n1804 , n1803 );
and ( n1805 , n1790 , n1804 );
and ( n1806 , n1805 , n1786 );
and ( n1807 , n1383 , n1137 );
not ( n1808 , n1807 );
and ( n1809 , n1808 , n1669 );
not ( n1810 , n1809 );
and ( n1811 , n1390 , n1082 );
not ( n1812 , n1811 );
not ( n1813 , n1681 );
and ( n1814 , n1083 , n1813 );
not ( n1815 , n1814 );
and ( n1816 , n1812 , n1815 );
not ( n1817 , n1816 );
and ( n1818 , n1082 , n1681 );
not ( n1819 , n1818 );
and ( n1820 , n1403 , n1121 );
not ( n1821 , n1820 );
and ( n1822 , n1821 , n1677 );
not ( n1823 , n1822 );
and ( n1824 , n1819 , n1823 );
and ( n1825 , n1817 , n1824 );
and ( n1826 , n1810 , n1825 );
not ( n1827 , n1826 );
and ( n1828 , n1807 , n1668 );
not ( n1829 , n1828 );
and ( n1830 , n1820 , n1686 );
and ( n1831 , n1830 , n1810 );
not ( n1832 , n1831 );
and ( n1833 , n1829 , n1832 );
and ( n1834 , n1827 , n1833 );
not ( n1835 , n1834 );
and ( n1836 , n1806 , n1835 );
not ( n1837 , n1836 );
and ( n1838 , n1802 , n1837 );
not ( n1839 , n1838 );
and ( n1840 , n1775 , n1839 );
not ( n1841 , n1840 );
and ( n1842 , n1770 , n1841 );
and ( n1843 , n1716 , n1842 );
not ( n1844 , n1843 );
not ( n1845 , n1716 );
not ( n1846 , n1842 );
and ( n1847 , n1845 , n1846 );
not ( n1848 , n1847 );
and ( n1849 , n1844 , n1848 );
not ( n1850 , n1849 );
and ( n1851 , n1715 , n1850 );
not ( n1852 , n1851 );
and ( n1853 , n1711 , n1852 );
and ( n1854 , n1212 , n1853 );
not ( n1855 , n1854 );
and ( n1856 , n794 , n1855 );
not ( n1857 , n1856 );
and ( n1858 , n797 , n1857 );
not ( n1859 , n1858 );
buf ( n1860 , n1859 );
buf ( n1861 , n1860 );
buf ( n1862 , n529 );
and ( n1863 , n709 , n758 , n776 , n793 );
not ( n1864 , n1863 );
and ( n1865 , n1862 , n1864 );
not ( n1866 , n1865 );
buf ( n1867 , n530 );
and ( n1868 , n1867 , n1229 );
and ( n1869 , n1868 , n1213 );
not ( n1870 , n1869 );
not ( n1871 , n1868 );
buf ( n1872 , n531 );
and ( n1873 , n1872 , n1229 );
not ( n1874 , n1873 );
buf ( n1875 , n532 );
and ( n1876 , n1875 , n1229 );
not ( n1877 , n1876 );
and ( n1878 , n1874 , n1877 );
buf ( n1879 , n533 );
and ( n1880 , n1879 , n1229 );
not ( n1881 , n1880 );
buf ( n1882 , n534 );
and ( n1883 , n1882 , n1229 );
not ( n1884 , n1883 );
and ( n1885 , n1881 , n1884 );
buf ( n1886 , n535 );
and ( n1887 , n1886 , n1229 );
not ( n1888 , n1887 );
buf ( n1889 , n536 );
and ( n1890 , n1889 , n1229 );
not ( n1891 , n1890 );
and ( n1892 , n1888 , n1891 );
and ( n1893 , n1885 , n1892 );
buf ( n1894 , n537 );
and ( n1895 , n1894 , n1229 );
not ( n1896 , n1895 );
buf ( n1897 , n538 );
and ( n1898 , n1897 , n1229 );
not ( n1899 , n1898 );
and ( n1900 , n1896 , n1899 );
buf ( n1901 , n539 );
and ( n1902 , n1901 , n1229 );
not ( n1903 , n1902 );
buf ( n1904 , n540 );
and ( n1905 , n1904 , n1229 );
not ( n1906 , n1905 );
and ( n1907 , n1903 , n1906 );
and ( n1908 , n1900 , n1907 );
buf ( n1909 , n541 );
and ( n1910 , n1909 , n1229 );
not ( n1911 , n1910 );
and ( n1912 , n600 , n606 );
not ( n1913 , n1912 );
xor ( n1914 , n606 , n657 );
not ( n1915 , n1914 );
and ( n1916 , n599 , n1915 );
not ( n1917 , n1916 );
and ( n1918 , n1913 , n1917 );
not ( n1919 , n1918 );
and ( n1920 , n1919 , n1228 );
not ( n1921 , n1920 );
and ( n1922 , n1911 , n1921 );
buf ( n1923 , n542 );
and ( n1924 , n1923 , n1229 );
not ( n1925 , n1924 );
and ( n1926 , n600 , n608 );
not ( n1927 , n1926 );
xor ( n1928 , n608 , n656 );
not ( n1929 , n1928 );
and ( n1930 , n599 , n1929 );
not ( n1931 , n1930 );
and ( n1932 , n1927 , n1931 );
not ( n1933 , n1932 );
and ( n1934 , n1933 , n1228 );
not ( n1935 , n1934 );
and ( n1936 , n1925 , n1935 );
and ( n1937 , n1922 , n1936 );
buf ( n1938 , n543 );
and ( n1939 , n1938 , n1229 );
not ( n1940 , n1939 );
and ( n1941 , n600 , n604 );
not ( n1942 , n1941 );
xor ( n1943 , n604 , n658 );
not ( n1944 , n1943 );
and ( n1945 , n599 , n1944 );
not ( n1946 , n1945 );
and ( n1947 , n1942 , n1946 );
not ( n1948 , n1947 );
and ( n1949 , n1948 , n1228 );
not ( n1950 , n1949 );
and ( n1951 , n1940 , n1950 );
buf ( n1952 , n544 );
and ( n1953 , n1952 , n1229 );
not ( n1954 , n1953 );
and ( n1955 , n1480 , n1228 );
not ( n1956 , n1955 );
and ( n1957 , n1954 , n1956 );
and ( n1958 , n1951 , n1957 );
and ( n1959 , n1937 , n1958 );
and ( n1960 , n1908 , n1959 );
and ( n1961 , n1878 , n1893 , n1960 );
and ( n1962 , n1263 , n1242 );
and ( n1963 , n1437 , n1384 , n1466 , n1962 );
and ( n1964 , n1325 , n1404 , n1354 , n1963 );
and ( n1965 , n1961 , n1964 );
not ( n1966 , n1965 );
and ( n1967 , n1871 , n1966 );
not ( n1968 , n1967 );
and ( n1969 , n1868 , n1965 );
not ( n1970 , n1969 );
and ( n1971 , n1968 , n1970 );
not ( n1972 , n1971 );
and ( n1973 , n1246 , n1972 );
not ( n1974 , n1973 );
and ( n1975 , n1870 , n1974 );
and ( n1976 , n769 , n810 );
not ( n1977 , n1976 );
and ( n1978 , n1229 , n1977 );
not ( n1979 , n1978 );
and ( n1980 , n702 , n1979 );
buf ( n1981 , n545 );
and ( n1982 , n1981 , n834 );
not ( n1983 , n1982 );
and ( n1984 , n1862 , n838 );
not ( n1985 , n1984 );
buf ( n1986 , n546 );
and ( n1987 , n1986 , n847 );
not ( n1988 , n1987 );
and ( n1989 , n1983 , n1985 , n1988 );
not ( n1990 , n1989 );
buf ( n1991 , n547 );
and ( n1992 , n1991 , n834 );
not ( n1993 , n1992 );
buf ( n1994 , n548 );
and ( n1995 , n1994 , n838 );
not ( n1996 , n1995 );
buf ( n1997 , n549 );
and ( n1998 , n1997 , n847 );
not ( n1999 , n1998 );
and ( n2000 , n1993 , n1996 , n1999 );
buf ( n2001 , n550 );
and ( n2002 , n2001 , n838 );
not ( n2003 , n2002 );
buf ( n2004 , n551 );
and ( n2005 , n2004 , n843 );
not ( n2006 , n2005 );
and ( n2007 , n2003 , n2006 );
buf ( n2008 , n552 );
and ( n2009 , n2008 , n847 );
not ( n2010 , n2009 );
buf ( n2011 , n553 );
and ( n2012 , n2011 , n834 );
not ( n2013 , n2012 );
and ( n2014 , n2010 , n2013 );
and ( n2015 , n2007 , n2014 );
not ( n2016 , n2015 );
buf ( n2017 , n554 );
and ( n2018 , n2017 , n834 );
not ( n2019 , n2018 );
buf ( n2020 , n555 );
and ( n2021 , n2020 , n847 );
not ( n2022 , n2021 );
and ( n2023 , n2019 , n2022 );
buf ( n2024 , n556 );
and ( n2025 , n2024 , n838 );
not ( n2026 , n2025 );
buf ( n2027 , n557 );
and ( n2028 , n2027 , n843 );
not ( n2029 , n2028 );
and ( n2030 , n2026 , n2029 );
and ( n2031 , n2023 , n2030 );
not ( n2032 , n2031 );
buf ( n2033 , n558 );
and ( n2034 , n2033 , n838 );
not ( n2035 , n2034 );
buf ( n2036 , n559 );
and ( n2037 , n2036 , n843 );
not ( n2038 , n2037 );
and ( n2039 , n2035 , n2038 );
buf ( n2040 , n560 );
and ( n2041 , n2040 , n847 );
not ( n2042 , n2041 );
buf ( n2043 , n561 );
and ( n2044 , n2043 , n834 );
not ( n2045 , n2044 );
and ( n2046 , n2042 , n2045 );
and ( n2047 , n2039 , n2046 );
not ( n2048 , n2047 );
and ( n2049 , n2032 , n2048 );
buf ( n2050 , n562 );
and ( n2051 , n2050 , n838 );
not ( n2052 , n2051 );
buf ( n2053 , n563 );
and ( n2054 , n2053 , n843 );
not ( n2055 , n2054 );
and ( n2056 , n2052 , n2055 );
buf ( n2057 , n564 );
and ( n2058 , n2057 , n834 );
not ( n2059 , n2058 );
buf ( n2060 , n565 );
and ( n2061 , n2060 , n847 );
not ( n2062 , n2061 );
and ( n2063 , n2059 , n2062 );
and ( n2064 , n2056 , n2063 );
not ( n2065 , n2064 );
buf ( n2066 , n566 );
and ( n2067 , n2066 , n838 );
not ( n2068 , n2067 );
buf ( n2069 , n567 );
and ( n2070 , n2069 , n843 );
not ( n2071 , n2070 );
and ( n2072 , n2068 , n2071 );
buf ( n2073 , n568 );
and ( n2074 , n2073 , n834 );
not ( n2075 , n2074 );
buf ( n2076 , n569 );
and ( n2077 , n2076 , n847 );
not ( n2078 , n2077 );
and ( n2079 , n2075 , n2078 );
and ( n2080 , n2072 , n2079 );
not ( n2081 , n2080 );
and ( n2082 , n2065 , n2081 );
and ( n2083 , n2049 , n2082 );
and ( n2084 , n2016 , n2083 );
buf ( n2085 , n570 );
and ( n2086 , n2085 , n834 );
not ( n2087 , n2086 );
buf ( n2088 , n571 );
and ( n2089 , n2088 , n838 );
not ( n2090 , n2089 );
buf ( n2091 , n572 );
and ( n2092 , n2091 , n843 );
not ( n2093 , n2092 );
buf ( n2094 , n573 );
and ( n2095 , n2094 , n847 );
not ( n2096 , n2095 );
and ( n2097 , n2087 , n2090 , n2093 , n2096 );
not ( n2098 , n2097 );
buf ( n2099 , n574 );
and ( n2100 , n2099 , n838 );
not ( n2101 , n2100 );
buf ( n2102 , n575 );
and ( n2103 , n2102 , n847 );
not ( n2104 , n2103 );
and ( n2105 , n2101 , n2104 );
buf ( n2106 , n576 );
and ( n2107 , n2106 , n843 );
not ( n2108 , n2107 );
buf ( n2109 , n577 );
and ( n2110 , n2109 , n834 );
not ( n2111 , n2110 );
and ( n2112 , n2108 , n2111 );
and ( n2113 , n2105 , n2112 );
not ( n2114 , n2113 );
buf ( n2115 , n578 );
and ( n2116 , n2115 , n838 );
not ( n2117 , n2116 );
buf ( n2118 , n579 );
and ( n2119 , n2118 , n847 );
not ( n2120 , n2119 );
and ( n2121 , n2117 , n2120 );
buf ( n2122 , n580 );
and ( n2123 , n2122 , n843 );
not ( n2124 , n2123 );
buf ( n2125 , n581 );
and ( n2126 , n2125 , n834 );
not ( n2127 , n2126 );
and ( n2128 , n2124 , n2127 );
and ( n2129 , n2121 , n2128 );
not ( n2130 , n2129 );
buf ( n2131 , n582 );
and ( n2132 , n2131 , n838 );
not ( n2133 , n2132 );
buf ( n2134 , n583 );
and ( n2135 , n2134 , n843 );
not ( n2136 , n2135 );
and ( n2137 , n2133 , n2136 );
buf ( n2138 , n584 );
and ( n2139 , n2138 , n834 );
not ( n2140 , n2139 );
buf ( n2141 , n585 );
and ( n2142 , n2141 , n847 );
not ( n2143 , n2142 );
and ( n2144 , n2140 , n2143 );
and ( n2145 , n2137 , n2144 );
not ( n2146 , n2145 );
and ( n2147 , n2098 , n2114 , n2130 , n2146 );
buf ( n2148 , n586 );
and ( n2149 , n2148 , n834 );
not ( n2150 , n2149 );
buf ( n2151 , n587 );
and ( n2152 , n2151 , n838 );
not ( n2153 , n2152 );
buf ( n2154 , n588 );
and ( n2155 , n2154 , n843 );
not ( n2156 , n2155 );
buf ( n2157 , n589 );
and ( n2158 , n2157 , n847 );
not ( n2159 , n2158 );
and ( n2160 , n2150 , n2153 , n2156 , n2159 );
not ( n2161 , n2160 );
not ( n2162 , n1036 );
and ( n2163 , n2161 , n2162 );
buf ( n2164 , n590 );
and ( n2165 , n2164 , n838 );
not ( n2166 , n2165 );
buf ( n2167 , n591 );
and ( n2168 , n2167 , n843 );
not ( n2169 , n2168 );
and ( n2170 , n2166 , n2169 );
buf ( n2171 , n592 );
and ( n2172 , n2171 , n834 );
not ( n2173 , n2172 );
buf ( n2174 , n593 );
and ( n2175 , n2174 , n847 );
not ( n2176 , n2175 );
and ( n2177 , n2173 , n2176 );
and ( n2178 , n2170 , n2177 );
not ( n2179 , n2178 );
buf ( n2180 , n594 );
and ( n2181 , n2180 , n838 );
not ( n2182 , n2181 );
buf ( n2183 , n595 );
and ( n2184 , n2183 , n843 );
not ( n2185 , n2184 );
and ( n2186 , n2182 , n2185 );
buf ( n2187 , n596 );
and ( n2188 , n2187 , n834 );
not ( n2189 , n2188 );
buf ( n2190 , n597 );
and ( n2191 , n2190 , n847 );
not ( n2192 , n2191 );
and ( n2193 , n2189 , n2192 );
and ( n2194 , n2186 , n2193 );
not ( n2195 , n2194 );
and ( n2196 , n2179 , n2195 );
and ( n2197 , n2163 , n2196 );
and ( n2198 , n2147 , n2197 );
and ( n2199 , n2084 , n2198 );
and ( n2200 , n1055 , n2199 );
not ( n2201 , n2200 );
and ( n2202 , n2000 , n2201 );
not ( n2203 , n2202 );
and ( n2204 , n2083 , n2198 );
and ( n2205 , n1055 , n2204 );
xor ( n2206 , n2015 , n2205 );
not ( n2207 , n2206 );
not ( n2208 , n2205 );
and ( n2209 , n2032 , n2082 );
and ( n2210 , n2209 , n2198 );
and ( n2211 , n1055 , n2210 );
not ( n2212 , n2211 );
and ( n2213 , n2047 , n2212 );
not ( n2214 , n2213 );
and ( n2215 , n2208 , n2214 );
and ( n2216 , n2082 , n2198 );
and ( n2217 , n1055 , n2216 );
not ( n2218 , n2217 );
and ( n2219 , n2065 , n2198 );
and ( n2220 , n1055 , n2219 );
not ( n2221 , n2220 );
and ( n2222 , n2080 , n2221 );
not ( n2223 , n2222 );
and ( n2224 , n2218 , n2223 );
and ( n2225 , n2031 , n2218 );
not ( n2226 , n2225 );
and ( n2227 , n2212 , n2226 );
and ( n2228 , n2224 , n2227 );
and ( n2229 , n2215 , n2228 );
and ( n2230 , n1055 , n2198 );
not ( n2231 , n2230 );
and ( n2232 , n2064 , n2231 );
not ( n2233 , n2232 );
and ( n2234 , n2221 , n2233 );
and ( n2235 , n2098 , n2146 );
and ( n2236 , n2163 , n2235 );
and ( n2237 , n2130 , n2195 );
and ( n2238 , n2114 , n2237 );
and ( n2239 , n2236 , n2238 );
and ( n2240 , n1055 , n2239 );
not ( n2241 , n2240 );
and ( n2242 , n2178 , n2241 );
not ( n2243 , n2242 );
and ( n2244 , n2231 , n2243 );
and ( n2245 , n2237 , n2236 );
and ( n2246 , n1055 , n2245 );
not ( n2247 , n2246 );
and ( n2248 , n2113 , n2247 );
not ( n2249 , n2248 );
and ( n2250 , n2241 , n2249 );
and ( n2251 , n2244 , n2250 );
and ( n2252 , n2234 , n2251 );
and ( n2253 , n1161 , n1194 );
and ( n2254 , n1177 , n2252 , n2253 );
and ( n2255 , n2146 , n2163 );
and ( n2256 , n2255 , n1055 );
not ( n2257 , n2256 );
and ( n2258 , n2163 , n1055 );
not ( n2259 , n2258 );
and ( n2260 , n2145 , n2259 );
not ( n2261 , n2260 );
and ( n2262 , n2257 , n2261 );
xor ( n2263 , n2097 , n2256 );
not ( n2264 , n2263 );
and ( n2265 , n2162 , n1055 );
not ( n2266 , n2265 );
and ( n2267 , n2160 , n2266 );
not ( n2268 , n2267 );
and ( n2269 , n2259 , n2268 );
and ( n2270 , n2264 , n2269 );
and ( n2271 , n2130 , n2236 );
and ( n2272 , n1055 , n2271 );
not ( n2273 , n2272 );
and ( n2274 , n2236 , n1055 );
not ( n2275 , n2274 );
and ( n2276 , n2129 , n2275 );
not ( n2277 , n2276 );
and ( n2278 , n2273 , n2277 );
and ( n2279 , n2194 , n2272 );
not ( n2280 , n2279 );
and ( n2281 , n2195 , n2273 );
not ( n2282 , n2281 );
and ( n2283 , n2280 , n2282 );
not ( n2284 , n2283 );
and ( n2285 , n2278 , n2284 );
and ( n2286 , n1093 , n1201 );
and ( n2287 , n1090 , n2286 );
and ( n2288 , n2262 , n2270 , n2285 , n2287 );
and ( n2289 , n1084 , n2288 );
and ( n2290 , n2229 , n2254 , n2289 );
and ( n2291 , n2207 , n2290 );
and ( n2292 , n2203 , n2291 );
and ( n2293 , n1990 , n2292 );
not ( n2294 , n2293 );
and ( n2295 , n1067 , n2294 );
and ( n2296 , n1980 , n2295 );
not ( n2297 , n2296 );
and ( n2298 , n1975 , n2297 );
not ( n2299 , n2298 );
and ( n2300 , n1863 , n2299 );
not ( n2301 , n2300 );
and ( n2302 , n1866 , n2301 );
not ( n2303 , n2302 );
buf ( n2304 , n2303 );
buf ( n2305 , n2304 );
and ( n2306 , n997 , n795 );
not ( n2307 , n2306 );
not ( n2308 , n1830 );
not ( n2309 , n1825 );
and ( n2310 , n2308 , n2309 );
and ( n2311 , n1829 , n1810 );
xor ( n2312 , n2310 , n2311 );
not ( n2313 , n2312 );
and ( n2314 , n1715 , n2313 );
not ( n2315 , n2314 );
and ( n2316 , n1649 , n1213 );
not ( n2317 , n2316 );
and ( n2318 , n1383 , n1404 );
not ( n2319 , n2318 );
and ( n2320 , n1369 , n2319 );
not ( n2321 , n2320 );
and ( n2322 , n1649 , n2318 );
not ( n2323 , n2322 );
and ( n2324 , n2321 , n2323 );
not ( n2325 , n2324 );
and ( n2326 , n1246 , n2325 );
not ( n2327 , n2326 );
and ( n2328 , n2317 , n2327 );
and ( n2329 , n1671 , n1674 );
not ( n2330 , n1678 );
not ( n2331 , n1689 );
and ( n2332 , n2330 , n2331 );
and ( n2333 , n2329 , n2332 );
not ( n2334 , n2333 );
not ( n2335 , n2329 );
not ( n2336 , n2332 );
and ( n2337 , n2335 , n2336 );
not ( n2338 , n2337 );
and ( n2339 , n2334 , n2338 );
not ( n2340 , n2339 );
and ( n2341 , n1484 , n2340 );
not ( n2342 , n2341 );
and ( n2343 , n2328 , n2342 );
and ( n2344 , n2315 , n2343 );
and ( n2345 , n811 , n1137 );
not ( n2346 , n2345 );
and ( n2347 , n1145 , n1084 );
not ( n2348 , n2347 );
and ( n2349 , n1121 , n1084 );
and ( n2350 , n1137 , n2349 );
and ( n2351 , n1107 , n2350 );
not ( n2352 , n2351 );
and ( n2353 , n1143 , n2352 );
not ( n2354 , n2353 );
and ( n2355 , n2348 , n2354 );
and ( n2356 , n810 , n2355 );
not ( n2357 , n2356 );
and ( n2358 , n2346 , n2357 );
not ( n2359 , n2358 );
and ( n2360 , n702 , n2359 );
not ( n2361 , n2360 );
and ( n2362 , n2344 , n2361 );
not ( n2363 , n2362 );
and ( n2364 , n794 , n2363 );
not ( n2365 , n2364 );
and ( n2366 , n2307 , n2365 );
not ( n2367 , n2366 );
buf ( n2368 , n2367 );
buf ( n2369 , n2368 );
and ( n2370 , n1122 , n1864 );
not ( n2371 , n2370 );
and ( n2372 , n1811 , n1819 );
not ( n2373 , n2372 );
and ( n2374 , n1815 , n2373 );
and ( n2375 , n2308 , n1823 );
and ( n2376 , n2374 , n2375 );
not ( n2377 , n2376 );
not ( n2378 , n2374 );
not ( n2379 , n2375 );
and ( n2380 , n2378 , n2379 );
not ( n2381 , n2380 );
and ( n2382 , n2377 , n2381 );
not ( n2383 , n2382 );
and ( n2384 , n1715 , n2383 );
not ( n2385 , n2384 );
and ( n2386 , n1213 , n1666 );
not ( n2387 , n2386 );
not ( n2388 , n1404 );
and ( n2389 , n1383 , n2388 );
not ( n2390 , n2389 );
and ( n2391 , n1666 , n1404 );
not ( n2392 , n2391 );
and ( n2393 , n2390 , n2392 );
not ( n2394 , n2393 );
and ( n2395 , n1246 , n2394 );
not ( n2396 , n2395 );
and ( n2397 , n2387 , n2396 );
not ( n2398 , n1684 );
and ( n2399 , n2330 , n1688 );
and ( n2400 , n2398 , n2399 );
not ( n2401 , n2400 );
not ( n2402 , n2399 );
and ( n2403 , n1684 , n2402 );
not ( n2404 , n2403 );
and ( n2405 , n2401 , n2404 );
not ( n2406 , n2405 );
and ( n2407 , n1484 , n2406 );
not ( n2408 , n2407 );
and ( n2409 , n2397 , n2408 );
and ( n2410 , n2385 , n2409 );
and ( n2411 , n811 , n1121 );
not ( n2412 , n2411 );
xor ( n2413 , n1107 , n2350 );
and ( n2414 , n810 , n2413 );
not ( n2415 , n2414 );
and ( n2416 , n2412 , n2415 );
not ( n2417 , n2416 );
and ( n2418 , n702 , n2417 );
not ( n2419 , n2418 );
and ( n2420 , n2410 , n2419 );
not ( n2421 , n2420 );
and ( n2422 , n1863 , n2421 );
not ( n2423 , n2422 );
and ( n2424 , n2371 , n2423 );
not ( n2425 , n2424 );
buf ( n2426 , n2425 );
buf ( n2427 , n2426 );
and ( n2428 , n720 , n675 );
and ( n2429 , n2428 , n702 , n756 );
not ( n2430 , n793 );
and ( n2431 , n719 , n777 , n2430 );
and ( n2432 , n2429 , n2431 );
and ( n2433 , n811 , n2284 );
not ( n2434 , n2433 );
not ( n2435 , n2244 );
and ( n2436 , n1161 , n1177 , n1194 );
and ( n2437 , n1084 , n2436 );
and ( n2438 , n2288 , n2437 );
and ( n2439 , n2250 , n2438 );
not ( n2440 , n2439 );
and ( n2441 , n2435 , n2440 );
not ( n2442 , n2441 );
and ( n2443 , n2244 , n2439 );
not ( n2444 , n2443 );
and ( n2445 , n2442 , n2444 );
and ( n2446 , n810 , n2445 );
not ( n2447 , n2446 );
and ( n2448 , n2434 , n2447 );
not ( n2449 , n2448 );
and ( n2450 , n2432 , n2449 );
not ( n2451 , n2450 );
not ( n2452 , n1483 );
and ( n2453 , n2452 , n706 );
and ( n2454 , n757 , n2431 );
and ( n2455 , n2453 , n2454 );
and ( n2456 , n1899 , n2195 );
and ( n2457 , n1902 , n2113 );
not ( n2458 , n2457 );
and ( n2459 , n1903 , n2114 );
not ( n2460 , n2459 );
and ( n2461 , n2458 , n2460 );
xor ( n2462 , n2456 , n2461 );
and ( n2463 , n1896 , n2130 );
and ( n2464 , n1898 , n2195 );
not ( n2465 , n2464 );
and ( n2466 , n1899 , n2194 );
not ( n2467 , n2466 );
and ( n2468 , n2465 , n2467 );
not ( n2469 , n2468 );
and ( n2470 , n2463 , n2469 );
not ( n2471 , n2470 );
not ( n2472 , n2463 );
and ( n2473 , n2472 , n2468 );
not ( n2474 , n2473 );
and ( n2475 , n1957 , n2098 );
and ( n2476 , n1895 , n2129 );
not ( n2477 , n2476 );
and ( n2478 , n2477 , n2472 );
and ( n2479 , n2475 , n2478 );
and ( n2480 , n2474 , n2479 );
not ( n2481 , n2480 );
and ( n2482 , n2471 , n2481 );
not ( n2483 , n2475 );
not ( n2484 , n2478 );
and ( n2485 , n2483 , n2484 );
not ( n2486 , n2485 );
and ( n2487 , n2474 , n2486 );
not ( n2488 , n1957 );
and ( n2489 , n2488 , n2097 );
not ( n2490 , n2489 );
and ( n2491 , n2483 , n2490 );
and ( n2492 , n1951 , n2146 );
and ( n2493 , n2491 , n2492 );
not ( n2494 , n2493 );
not ( n2495 , n2491 );
not ( n2496 , n2492 );
and ( n2497 , n2495 , n2496 );
not ( n2498 , n2497 );
and ( n2499 , n1922 , n2161 );
not ( n2500 , n1951 );
and ( n2501 , n2500 , n2145 );
not ( n2502 , n2501 );
and ( n2503 , n2502 , n2496 );
and ( n2504 , n2499 , n2503 );
and ( n2505 , n2498 , n2504 );
not ( n2506 , n2505 );
and ( n2507 , n2494 , n2506 );
not ( n2508 , n2499 );
not ( n2509 , n2503 );
and ( n2510 , n2508 , n2509 );
not ( n2511 , n2510 );
and ( n2512 , n2498 , n2511 );
and ( n2513 , n1936 , n2162 );
not ( n2514 , n1922 );
and ( n2515 , n2514 , n2161 );
not ( n2516 , n2515 );
and ( n2517 , n1922 , n2160 );
not ( n2518 , n2517 );
and ( n2519 , n2516 , n2518 );
not ( n2520 , n2519 );
and ( n2521 , n2513 , n2520 );
not ( n2522 , n2521 );
not ( n2523 , n2513 );
and ( n2524 , n2523 , n2519 );
not ( n2525 , n2524 );
not ( n2526 , n1936 );
and ( n2527 , n2526 , n1036 );
not ( n2528 , n2527 );
and ( n2529 , n2528 , n2523 );
and ( n2530 , n1487 , n2529 );
and ( n2531 , n2525 , n2530 );
not ( n2532 , n2531 );
and ( n2533 , n2522 , n2532 );
not ( n2534 , n2533 );
and ( n2535 , n2512 , n2534 );
not ( n2536 , n2535 );
and ( n2537 , n2507 , n2536 );
not ( n2538 , n2537 );
and ( n2539 , n2487 , n2538 );
not ( n2540 , n2539 );
and ( n2541 , n2482 , n2540 );
not ( n2542 , n2529 );
and ( n2543 , n1488 , n2542 );
not ( n2544 , n2543 );
and ( n2545 , n2525 , n2544 );
and ( n2546 , n2545 , n2512 );
and ( n2547 , n2487 , n2546 );
and ( n2548 , n1503 , n1492 );
not ( n2549 , n2548 );
and ( n2550 , n1722 , n2549 );
and ( n2551 , n1737 , n2550 );
not ( n2552 , n1786 );
and ( n2553 , n1783 , n2552 );
not ( n2554 , n2553 );
and ( n2555 , n1777 , n1788 , n1782 , n1797 );
not ( n2556 , n2555 );
and ( n2557 , n1774 , n2551 , n2554 , n2556 );
not ( n2558 , n2557 );
and ( n2559 , n2551 , n1764 );
not ( n2560 , n2559 );
and ( n2561 , n2308 , n1829 );
and ( n2562 , n2309 , n2561 );
not ( n2563 , n2562 );
and ( n2564 , n1757 , n1773 );
and ( n2565 , n1753 , n1805 , n2564 , n1810 );
and ( n2566 , n2551 , n2554 , n2563 , n2565 );
not ( n2567 , n2566 );
and ( n2568 , n1502 , n1491 );
not ( n2569 , n2568 );
and ( n2570 , n1718 , n2549 );
not ( n2571 , n2570 );
and ( n2572 , n2569 , n2571 );
and ( n2573 , n2550 , n1731 );
not ( n2574 , n2573 );
and ( n2575 , n2572 , n2574 );
not ( n2576 , n1749 );
and ( n2577 , n2551 , n2576 );
not ( n2578 , n2577 );
and ( n2579 , n2575 , n2578 );
and ( n2580 , n2558 , n2560 , n2567 , n2579 );
not ( n2581 , n2580 );
and ( n2582 , n2547 , n2581 );
not ( n2583 , n2582 );
and ( n2584 , n2541 , n2583 );
not ( n2585 , n2584 );
and ( n2586 , n2462 , n2585 );
not ( n2587 , n2586 );
not ( n2588 , n2462 );
and ( n2589 , n2588 , n2584 );
not ( n2590 , n2589 );
and ( n2591 , n2587 , n2590 );
and ( n2592 , n2455 , n2591 );
not ( n2593 , n2592 );
not ( n2594 , n720 );
and ( n2595 , n2594 , n2106 );
not ( n2596 , n2595 );
and ( n2597 , n2428 , n704 , n756 );
and ( n2598 , n2597 , n2431 );
and ( n2599 , n1900 , n1959 );
and ( n2600 , n2599 , n1964 );
not ( n2601 , n2600 );
and ( n2602 , n1903 , n2601 );
not ( n2603 , n2602 );
and ( n2604 , n1902 , n2600 );
not ( n2605 , n2604 );
and ( n2606 , n2603 , n2605 );
not ( n2607 , n2606 );
and ( n2608 , n2598 , n2607 );
not ( n2609 , n2608 );
and ( n2610 , n2596 , n2609 );
and ( n2611 , n1480 , n674 );
and ( n2612 , n720 , n2611 );
and ( n2613 , n719 , n2612 , n704 , n756 );
not ( n2614 , n2613 );
and ( n2615 , n1213 , n2454 );
not ( n2616 , n2615 );
and ( n2617 , n2614 , n2616 );
not ( n2618 , n2617 );
and ( n2619 , n1902 , n2618 );
not ( n2620 , n2619 );
and ( n2621 , n1003 , n960 );
and ( n2622 , n946 , n2621 );
and ( n2623 , n989 , n2622 );
and ( n2624 , n975 , n2623 );
and ( n2625 , n930 , n2624 );
and ( n2626 , n916 , n2625 );
and ( n2627 , n902 , n2626 );
and ( n2628 , n888 , n2627 );
and ( n2629 , n857 , n2628 );
and ( n2630 , n868 , n2629 );
and ( n2631 , n841 , n2630 );
and ( n2632 , n1043 , n2631 );
and ( n2633 , n1030 , n2632 );
and ( n2634 , n2154 , n2633 );
and ( n2635 , n2134 , n2634 );
and ( n2636 , n2091 , n2635 );
and ( n2637 , n2122 , n2636 );
and ( n2638 , n2183 , n2637 );
xor ( n2639 , n2106 , n2638 );
not ( n2640 , n2455 );
and ( n2641 , n1484 , n2454 );
not ( n2642 , n2641 );
not ( n2643 , n2432 );
and ( n2644 , n720 , n2643 );
and ( n2645 , n2640 , n2642 , n2644 );
not ( n2646 , n2598 );
and ( n2647 , n2646 , n2617 );
and ( n2648 , n2645 , n2647 );
and ( n2649 , n2639 , n2648 );
not ( n2650 , n2649 );
and ( n2651 , n2610 , n2620 , n2650 );
not ( n2652 , n2461 );
and ( n2653 , n2464 , n2652 );
not ( n2654 , n2653 );
and ( n2655 , n2465 , n2461 );
not ( n2656 , n2655 );
and ( n2657 , n2654 , n2656 );
and ( n2658 , n1895 , n2130 );
and ( n2659 , n2658 , n2468 );
not ( n2660 , n2659 );
and ( n2661 , n2488 , n2098 );
and ( n2662 , n2661 , n2484 );
not ( n2663 , n2658 );
and ( n2664 , n2663 , n2469 );
not ( n2665 , n2664 );
and ( n2666 , n2662 , n2665 );
not ( n2667 , n2666 );
and ( n2668 , n2660 , n2667 );
not ( n2669 , n2661 );
and ( n2670 , n2669 , n2478 );
not ( n2671 , n2670 );
and ( n2672 , n2665 , n2671 );
and ( n2673 , n2500 , n2146 );
not ( n2674 , n2673 );
and ( n2675 , n2491 , n2674 );
not ( n2676 , n2675 );
and ( n2677 , n2516 , n2503 );
not ( n2678 , n2677 );
and ( n2679 , n2676 , n2678 );
and ( n2680 , n2526 , n2162 );
and ( n2681 , n2680 , n2519 );
not ( n2682 , n2681 );
and ( n2683 , n1243 , n1050 );
and ( n2684 , n2683 , n2542 );
not ( n2685 , n2680 );
and ( n2686 , n2685 , n2520 );
not ( n2687 , n2686 );
and ( n2688 , n2684 , n2687 );
not ( n2689 , n2688 );
and ( n2690 , n2682 , n2689 );
not ( n2691 , n2690 );
and ( n2692 , n2679 , n2691 );
not ( n2693 , n2692 );
and ( n2694 , n2495 , n2673 );
not ( n2695 , n2694 );
and ( n2696 , n2515 , n2509 );
and ( n2697 , n2676 , n2696 );
not ( n2698 , n2697 );
and ( n2699 , n2695 , n2698 );
and ( n2700 , n2693 , n2699 );
not ( n2701 , n2700 );
and ( n2702 , n2672 , n2701 );
not ( n2703 , n2702 );
and ( n2704 , n2668 , n2703 );
not ( n2705 , n2683 );
and ( n2706 , n2705 , n2529 );
not ( n2707 , n2706 );
and ( n2708 , n2687 , n2707 );
and ( n2709 , n2679 , n2708 );
and ( n2710 , n2672 , n2709 );
and ( n2711 , n1508 , n1497 );
not ( n2712 , n2711 );
and ( n2713 , n1583 , n1497 );
not ( n2714 , n2713 );
and ( n2715 , n1494 , n2714 );
and ( n2716 , n2712 , n2715 );
not ( n2717 , n2716 );
and ( n2718 , n1528 , n1553 , n1578 );
not ( n2719 , n2718 );
and ( n2720 , n1591 , n2715 );
and ( n2721 , n2719 , n2720 );
not ( n2722 , n2721 );
and ( n2723 , n2717 , n2722 );
not ( n2724 , n2723 );
not ( n2725 , n1629 );
and ( n2726 , n2725 , n1625 );
not ( n2727 , n2726 );
and ( n2728 , n2711 , n1528 , n1601 , n2727 );
and ( n2729 , n1671 , n2330 , n2331 );
not ( n2730 , n2729 );
and ( n2731 , n1674 , n1664 , n2730 );
not ( n2732 , n2731 );
and ( n2733 , n1625 , n1657 );
and ( n2734 , n2732 , n2733 );
not ( n2735 , n2734 );
and ( n2736 , n2728 , n2735 );
not ( n2737 , n2736 );
and ( n2738 , n2724 , n2737 );
not ( n2739 , n2738 );
and ( n2740 , n2710 , n2739 );
not ( n2741 , n2740 );
and ( n2742 , n2704 , n2741 );
not ( n2743 , n2742 );
and ( n2744 , n2657 , n2743 );
not ( n2745 , n2744 );
not ( n2746 , n2657 );
and ( n2747 , n2746 , n2742 );
not ( n2748 , n2747 );
and ( n2749 , n2745 , n2748 );
and ( n2750 , n2641 , n2749 );
not ( n2751 , n2750 );
and ( n2752 , n2651 , n2751 );
and ( n2753 , n2593 , n2752 );
and ( n2754 , n2451 , n2753 );
not ( n2755 , n2754 );
buf ( n2756 , n2755 );
buf ( n2757 , n2756 );
and ( n2758 , n2050 , n1864 );
not ( n2759 , n2758 );
and ( n2760 , n811 , n2244 );
not ( n2761 , n2760 );
and ( n2762 , n2288 , n2254 );
and ( n2763 , n1084 , n2762 );
and ( n2764 , n2224 , n2763 );
not ( n2765 , n2764 );
not ( n2766 , n2224 );
not ( n2767 , n2763 );
and ( n2768 , n2766 , n2767 );
not ( n2769 , n2768 );
and ( n2770 , n2765 , n2769 );
and ( n2771 , n810 , n2770 );
not ( n2772 , n2771 );
and ( n2773 , n2761 , n2772 );
not ( n2774 , n2773 );
and ( n2775 , n702 , n2774 );
not ( n2776 , n2775 );
and ( n2777 , n1906 , n2179 );
not ( n2778 , n2777 );
and ( n2779 , n1883 , n2065 );
not ( n2780 , n2779 );
and ( n2781 , n1884 , n2064 );
not ( n2782 , n2781 );
and ( n2783 , n2780 , n2782 );
xor ( n2784 , n2778 , n2783 );
and ( n2785 , n1905 , n2179 );
not ( n2786 , n2785 );
and ( n2787 , n1906 , n2178 );
not ( n2788 , n2787 );
and ( n2789 , n2786 , n2788 );
not ( n2790 , n2789 );
and ( n2791 , n2459 , n2790 );
not ( n2792 , n2791 );
and ( n2793 , n2456 , n2461 );
and ( n2794 , n2460 , n2789 );
not ( n2795 , n2794 );
and ( n2796 , n2793 , n2795 );
not ( n2797 , n2796 );
and ( n2798 , n2792 , n2797 );
not ( n2799 , n2456 );
and ( n2800 , n2799 , n2652 );
not ( n2801 , n2800 );
and ( n2802 , n2801 , n2795 );
not ( n2803 , n2482 );
and ( n2804 , n2802 , n2803 );
not ( n2805 , n2804 );
and ( n2806 , n2798 , n2805 );
and ( n2807 , n2487 , n2802 );
and ( n2808 , n2807 , n2538 );
not ( n2809 , n2808 );
and ( n2810 , n2806 , n2809 );
and ( n2811 , n2807 , n2546 );
and ( n2812 , n2811 , n2581 );
not ( n2813 , n2812 );
and ( n2814 , n2810 , n2813 );
not ( n2815 , n2814 );
and ( n2816 , n2784 , n2815 );
not ( n2817 , n2816 );
not ( n2818 , n2784 );
and ( n2819 , n2818 , n2814 );
not ( n2820 , n2819 );
and ( n2821 , n2817 , n2820 );
and ( n2822 , n1715 , n2821 );
not ( n2823 , n2822 );
and ( n2824 , n1883 , n1213 );
not ( n2825 , n2824 );
and ( n2826 , n1960 , n1964 );
not ( n2827 , n2826 );
and ( n2828 , n1884 , n2827 );
not ( n2829 , n2828 );
and ( n2830 , n1883 , n2826 );
not ( n2831 , n2830 );
and ( n2832 , n2829 , n2831 );
not ( n2833 , n2832 );
and ( n2834 , n1246 , n2833 );
not ( n2835 , n2834 );
and ( n2836 , n2825 , n2835 );
not ( n2837 , n2783 );
and ( n2838 , n2786 , n2837 );
not ( n2839 , n2838 );
and ( n2840 , n2785 , n2783 );
not ( n2841 , n2840 );
and ( n2842 , n2839 , n2841 );
and ( n2843 , n1902 , n2114 );
and ( n2844 , n2843 , n2789 );
not ( n2845 , n2844 );
not ( n2846 , n2843 );
and ( n2847 , n2846 , n2790 );
not ( n2848 , n2847 );
and ( n2849 , n2653 , n2848 );
not ( n2850 , n2849 );
and ( n2851 , n2845 , n2850 );
and ( n2852 , n2668 , n2851 );
and ( n2853 , n2693 , n2852 , n2699 );
not ( n2854 , n2853 );
not ( n2855 , n2672 );
and ( n2856 , n2855 , n2852 );
not ( n2857 , n2856 );
and ( n2858 , n2656 , n2848 );
not ( n2859 , n2858 );
and ( n2860 , n2859 , n2851 );
not ( n2861 , n2860 );
and ( n2862 , n2857 , n2861 );
and ( n2863 , n2854 , n2862 );
not ( n2864 , n2863 );
and ( n2865 , n2858 , n2672 );
and ( n2866 , n2865 , n2709 );
and ( n2867 , n2866 , n2739 );
not ( n2868 , n2867 );
and ( n2869 , n2864 , n2868 );
not ( n2870 , n2869 );
and ( n2871 , n2842 , n2870 );
not ( n2872 , n2871 );
not ( n2873 , n2842 );
and ( n2874 , n2873 , n2869 );
not ( n2875 , n2874 );
and ( n2876 , n2872 , n2875 );
and ( n2877 , n1484 , n2876 );
not ( n2878 , n2877 );
and ( n2879 , n2836 , n2878 );
and ( n2880 , n2823 , n2879 );
and ( n2881 , n2776 , n2880 );
not ( n2882 , n2881 );
and ( n2883 , n1863 , n2882 );
not ( n2884 , n2883 );
and ( n2885 , n2759 , n2884 );
not ( n2886 , n2885 );
buf ( n2887 , n2886 );
buf ( n2888 , n2887 );
and ( n2889 , n776 , n2430 );
and ( n2890 , n758 , n2889 );
and ( n2891 , n2453 , n2890 );
and ( n2892 , n2522 , n2525 );
not ( n2893 , n2530 );
and ( n2894 , n2544 , n2581 );
not ( n2895 , n2894 );
and ( n2896 , n2893 , n2895 );
xor ( n2897 , n2892 , n2896 );
not ( n2898 , n2897 );
and ( n2899 , n2891 , n2898 );
not ( n2900 , n2899 );
and ( n2901 , n675 , n702 );
and ( n2902 , n2901 , n2890 );
and ( n2903 , n811 , n1201 );
not ( n2904 , n2903 );
not ( n2905 , n2262 );
and ( n2906 , n1201 , n1090 );
and ( n2907 , n2269 , n2906 );
and ( n2908 , n2907 , n1196 );
and ( n2909 , n1084 , n2908 );
and ( n2910 , n2905 , n2909 );
not ( n2911 , n2910 );
not ( n2912 , n2909 );
and ( n2913 , n2262 , n2912 );
not ( n2914 , n2913 );
and ( n2915 , n2911 , n2914 );
not ( n2916 , n2915 );
and ( n2917 , n810 , n2916 );
not ( n2918 , n2917 );
and ( n2919 , n2904 , n2918 );
not ( n2920 , n2919 );
and ( n2921 , n2902 , n2920 );
not ( n2922 , n2921 );
and ( n2923 , n709 , n777 );
not ( n2924 , n2923 );
and ( n2925 , n676 , n702 );
not ( n2926 , n2925 );
and ( n2927 , n719 , n2926 , n757 );
and ( n2928 , n2611 , n704 );
not ( n2929 , n2928 );
and ( n2930 , n2929 , n793 );
not ( n2931 , n2930 );
and ( n2932 , n2927 , n2931 );
and ( n2933 , n2924 , n2932 );
not ( n2934 , n2933 );
and ( n2935 , n2157 , n2934 );
not ( n2936 , n2935 );
and ( n2937 , n1936 , n1964 );
not ( n2938 , n2937 );
and ( n2939 , n1922 , n2938 );
not ( n2940 , n2939 );
and ( n2941 , n2514 , n2937 );
not ( n2942 , n2941 );
and ( n2943 , n2940 , n2942 );
not ( n2944 , n2943 );
and ( n2945 , n1246 , n2890 );
and ( n2946 , n2944 , n2945 );
not ( n2947 , n2946 );
xor ( n2948 , n2154 , n2633 );
and ( n2949 , n2948 , n2613 );
not ( n2950 , n2949 );
and ( n2951 , n1213 , n2890 );
and ( n2952 , n2514 , n2951 );
not ( n2953 , n2952 );
and ( n2954 , n2950 , n2953 );
and ( n2955 , n2936 , n2947 , n2954 );
and ( n2956 , n1484 , n2890 );
and ( n2957 , n2682 , n2687 );
not ( n2958 , n2684 );
and ( n2959 , n2707 , n2739 );
not ( n2960 , n2959 );
and ( n2961 , n2958 , n2960 );
and ( n2962 , n2957 , n2961 );
not ( n2963 , n2962 );
not ( n2964 , n2957 );
not ( n2965 , n2961 );
and ( n2966 , n2964 , n2965 );
not ( n2967 , n2966 );
and ( n2968 , n2963 , n2967 );
not ( n2969 , n2968 );
and ( n2970 , n2956 , n2969 );
not ( n2971 , n2970 );
and ( n2972 , n2955 , n2971 );
and ( n2973 , n2900 , n2922 , n2972 );
not ( n2974 , n2973 );
buf ( n2975 , n2974 );
buf ( n2976 , n2975 );
not ( n2977 , n2504 );
and ( n2978 , n2511 , n2977 );
and ( n2979 , n2545 , n2581 );
not ( n2980 , n2979 );
and ( n2981 , n2533 , n2980 );
xor ( n2982 , n2978 , n2981 );
not ( n2983 , n2982 );
and ( n2984 , n2891 , n2983 );
not ( n2985 , n2984 );
and ( n2986 , n2141 , n2934 );
not ( n2987 , n2986 );
and ( n2988 , n1937 , n1964 );
not ( n2989 , n2988 );
and ( n2990 , n1951 , n2989 );
not ( n2991 , n2990 );
and ( n2992 , n2500 , n2988 );
not ( n2993 , n2992 );
and ( n2994 , n2991 , n2993 );
not ( n2995 , n2994 );
and ( n2996 , n2995 , n2945 );
not ( n2997 , n2996 );
xor ( n2998 , n2134 , n2634 );
and ( n2999 , n2998 , n2613 );
not ( n3000 , n2999 );
and ( n3001 , n2500 , n2951 );
not ( n3002 , n3001 );
and ( n3003 , n3000 , n3002 );
and ( n3004 , n2987 , n2997 , n3003 );
not ( n3005 , n2696 );
and ( n3006 , n3005 , n2678 );
and ( n3007 , n2708 , n2739 );
not ( n3008 , n3007 );
and ( n3009 , n2690 , n3008 );
and ( n3010 , n3006 , n3009 );
not ( n3011 , n3010 );
not ( n3012 , n3006 );
not ( n3013 , n3009 );
and ( n3014 , n3012 , n3013 );
not ( n3015 , n3014 );
and ( n3016 , n3011 , n3015 );
not ( n3017 , n3016 );
and ( n3018 , n2956 , n3017 );
not ( n3019 , n3018 );
and ( n3020 , n3004 , n3019 );
and ( n3021 , n2985 , n3020 );
and ( n3022 , n811 , n2269 );
not ( n3023 , n3022 );
and ( n3024 , n2262 , n2909 );
not ( n3025 , n3024 );
and ( n3026 , n2264 , n3025 );
not ( n3027 , n3026 );
and ( n3028 , n2263 , n3024 );
not ( n3029 , n3028 );
and ( n3030 , n3027 , n3029 );
not ( n3031 , n3030 );
and ( n3032 , n810 , n3031 );
not ( n3033 , n3032 );
and ( n3034 , n3023 , n3033 );
not ( n3035 , n3034 );
and ( n3036 , n2902 , n3035 );
not ( n3037 , n3036 );
and ( n3038 , n3021 , n3037 );
not ( n3039 , n3038 );
buf ( n3040 , n3039 );
buf ( n3041 , n3040 );
and ( n3042 , n2594 , n946 );
not ( n3043 , n3042 );
and ( n3044 , n1465 , n1405 );
not ( n3045 , n3044 );
and ( n3046 , n1436 , n3045 );
not ( n3047 , n3046 );
and ( n3048 , n1614 , n3044 );
not ( n3049 , n3048 );
and ( n3050 , n3047 , n3049 );
not ( n3051 , n3050 );
and ( n3052 , n3051 , n2598 );
not ( n3053 , n3052 );
and ( n3054 , n3043 , n3053 );
and ( n3055 , n1614 , n2618 );
not ( n3056 , n3055 );
and ( n3057 , n3054 , n3056 );
xor ( n3058 , n946 , n2621 );
and ( n3059 , n3058 , n2648 );
not ( n3060 , n3059 );
and ( n3061 , n1639 , n1642 );
not ( n3062 , n1654 );
and ( n3063 , n1663 , n1693 );
not ( n3064 , n3063 );
and ( n3065 , n3062 , n3064 );
and ( n3066 , n3061 , n3065 );
not ( n3067 , n3066 );
not ( n3068 , n3061 );
not ( n3069 , n3065 );
and ( n3070 , n3068 , n3069 );
not ( n3071 , n3070 );
and ( n3072 , n3067 , n3071 );
not ( n3073 , n3072 );
and ( n3074 , n2641 , n3073 );
not ( n3075 , n3074 );
and ( n3076 , n1790 , n1788 );
not ( n3077 , n1795 );
and ( n3078 , n1804 , n1835 );
not ( n3079 , n3078 );
and ( n3080 , n3077 , n3079 );
and ( n3081 , n3076 , n3080 );
not ( n3082 , n3081 );
not ( n3083 , n3076 );
not ( n3084 , n3080 );
and ( n3085 , n3083 , n3084 );
not ( n3086 , n3085 );
and ( n3087 , n3082 , n3086 );
not ( n3088 , n3087 );
and ( n3089 , n2455 , n3088 );
not ( n3090 , n3089 );
and ( n3091 , n3057 , n3060 , n3075 , n3090 );
and ( n3092 , n811 , n1144 );
not ( n3093 , n3092 );
and ( n3094 , n1158 , n2347 );
and ( n3095 , n1152 , n3094 );
not ( n3096 , n3095 );
not ( n3097 , n3094 );
and ( n3098 , n1153 , n3097 );
not ( n3099 , n3098 );
and ( n3100 , n3096 , n3099 );
not ( n3101 , n3100 );
and ( n3102 , n810 , n3101 );
not ( n3103 , n3102 );
and ( n3104 , n3093 , n3103 );
not ( n3105 , n3104 );
and ( n3106 , n2432 , n3105 );
not ( n3107 , n3106 );
and ( n3108 , n3091 , n3107 );
not ( n3109 , n3108 );
buf ( n3110 , n3109 );
buf ( n3111 , n3110 );
and ( n3112 , n2017 , n795 );
not ( n3113 , n3112 );
and ( n3114 , n811 , n2224 );
not ( n3115 , n3114 );
not ( n3116 , n2290 );
not ( n3117 , n2215 );
and ( n3118 , n1084 , n2228 , n2762 );
not ( n3119 , n3118 );
and ( n3120 , n3117 , n3119 );
not ( n3121 , n3120 );
and ( n3122 , n3116 , n3121 );
and ( n3123 , n810 , n3122 );
not ( n3124 , n3123 );
and ( n3125 , n3115 , n3124 );
not ( n3126 , n3125 );
and ( n3127 , n702 , n3126 );
not ( n3128 , n3127 );
and ( n3129 , n1887 , n1213 );
not ( n3130 , n3129 );
and ( n3131 , n1885 , n1937 , n1908 , n1958 );
and ( n3132 , n3131 , n1964 );
not ( n3133 , n3132 );
and ( n3134 , n1888 , n3133 );
not ( n3135 , n3134 );
and ( n3136 , n1887 , n3132 );
not ( n3137 , n3136 );
and ( n3138 , n3135 , n3137 );
not ( n3139 , n3138 );
and ( n3140 , n1246 , n3139 );
not ( n3141 , n3140 );
and ( n3142 , n3130 , n3141 );
and ( n3143 , n1880 , n2081 );
and ( n3144 , n1887 , n2032 );
not ( n3145 , n3144 );
and ( n3146 , n1888 , n2031 );
not ( n3147 , n3146 );
and ( n3148 , n3145 , n3147 );
and ( n3149 , n3143 , n3148 );
not ( n3150 , n3149 );
not ( n3151 , n3143 );
not ( n3152 , n3148 );
and ( n3153 , n3151 , n3152 );
not ( n3154 , n3153 );
and ( n3155 , n3150 , n3154 );
xor ( n3156 , n1880 , n2080 );
not ( n3157 , n3156 );
and ( n3158 , n2779 , n3157 );
not ( n3159 , n3158 );
and ( n3160 , n2780 , n3156 );
not ( n3161 , n3160 );
and ( n3162 , n3161 , n2840 );
not ( n3163 , n3162 );
and ( n3164 , n3159 , n3163 );
and ( n3165 , n3161 , n2839 );
and ( n3166 , n3165 , n2863 );
not ( n3167 , n3166 );
and ( n3168 , n3164 , n3167 );
and ( n3169 , n3165 , n2866 );
and ( n3170 , n3169 , n2739 );
not ( n3171 , n3170 );
and ( n3172 , n3168 , n3171 );
not ( n3173 , n3172 );
and ( n3174 , n3155 , n3173 );
not ( n3175 , n3174 );
not ( n3176 , n3155 );
and ( n3177 , n3176 , n3172 );
not ( n3178 , n3177 );
and ( n3179 , n3175 , n3178 );
and ( n3180 , n1484 , n3179 );
not ( n3181 , n3180 );
and ( n3182 , n3142 , n3181 );
and ( n3183 , n1881 , n2081 );
not ( n3184 , n3183 );
xor ( n3185 , n3184 , n3148 );
and ( n3186 , n2778 , n2783 );
not ( n3187 , n3186 );
and ( n3188 , n1884 , n2065 );
not ( n3189 , n3188 );
and ( n3190 , n3189 , n3157 );
not ( n3191 , n3190 );
and ( n3192 , n3187 , n3191 );
and ( n3193 , n3192 , n2811 );
and ( n3194 , n3193 , n2581 );
not ( n3195 , n3194 );
and ( n3196 , n3188 , n3156 );
not ( n3197 , n3196 );
and ( n3198 , n2777 , n2837 );
and ( n3199 , n3198 , n3191 );
not ( n3200 , n3199 );
and ( n3201 , n3197 , n3200 );
not ( n3202 , n2810 );
and ( n3203 , n3192 , n3202 );
not ( n3204 , n3203 );
and ( n3205 , n3201 , n3204 );
and ( n3206 , n3195 , n3205 );
not ( n3207 , n3206 );
and ( n3208 , n3185 , n3207 );
not ( n3209 , n3208 );
not ( n3210 , n3185 );
and ( n3211 , n3210 , n3206 );
not ( n3212 , n3211 );
and ( n3213 , n3209 , n3212 );
and ( n3214 , n1715 , n3213 );
not ( n3215 , n3214 );
and ( n3216 , n3182 , n3215 );
and ( n3217 , n3128 , n3216 );
not ( n3218 , n3217 );
and ( n3219 , n794 , n3218 );
not ( n3220 , n3219 );
and ( n3221 , n3113 , n3220 );
not ( n3222 , n3221 );
buf ( n3223 , n3222 );
buf ( n3224 , n3223 );
endmodule

