//
// Conformal-LEC Version 16.10-d005 ( 21-Apr-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 ;
output n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 ;

wire n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
     n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
     n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
     n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
     n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
     n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
     n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
     n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
     n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
     n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
     n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
     n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
     n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
     n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
     n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
     n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
     n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
     n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
     n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
     n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
     n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
     n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
     n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
     n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
     n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , 
     n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , 
     n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
     n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , 
     n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
     n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , 
     n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
     n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
     n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
     n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , 
     n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
     n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
     n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
     n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
     n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
     n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
     n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
     n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
     n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
     n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
     n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
     n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
     n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , 
     n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , 
     n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , 
     n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , 
     n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , 
     n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , 
     n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , 
     n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
     n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , 
     n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , 
     n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , 
     n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , 
     n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , 
     n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , 
     n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , 
     n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , 
     n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , 
     n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , 
     n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , 
     n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , 
     n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , 
     n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , 
     n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
     n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
     n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
     n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
     n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
     n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
     n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
     n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
     n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
     n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
     n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
     n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
     n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
     n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
     n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , 
     n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , 
     n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
     n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , 
     n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , 
     n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , 
     n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , 
     n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , 
     n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , 
     n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , 
     n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , 
     n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
     n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , 
     n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , 
     n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , 
     n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
     n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , 
     n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , 
     n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
     n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , 
     n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , 
     n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , 
     n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , 
     n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , 
     n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , 
     n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , 
     n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , 
     n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , 
     n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , 
     n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , 
     n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , 
     n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , 
     n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , 
     n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , 
     n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , 
     n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , 
     n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , 
     n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
     n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , 
     n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , 
     n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , 
     n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , 
     n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , 
     n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , 
     n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , 
     n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , 
     n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , 
     n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , 
     n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , 
     n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , 
     n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , 
     n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , 
     n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , 
     n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , 
     n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , 
     n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , 
     n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , 
     n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , 
     n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , 
     n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , 
     n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , 
     n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , 
     n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , 
     n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , 
     n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , 
     n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , 
     n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , 
     n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , 
     n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , 
     n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , 
     n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , 
     n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , 
     n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , 
     n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , 
     n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , 
     n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , 
     n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , 
     n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , 
     n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , 
     n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , 
     n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , 
     n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , 
     n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , 
     n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , 
     n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , 
     n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , 
     n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , 
     n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , 
     n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , 
     n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , 
     n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , 
     n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , 
     n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , 
     n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , 
     n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , 
     n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , 
     n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , 
     n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , 
     n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , 
     n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , 
     n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , 
     n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , 
     n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , 
     n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , 
     n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , 
     n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , 
     n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , 
     n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , 
     n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , 
     n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , 
     n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , 
     n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , 
     n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , 
     n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , 
     n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , 
     n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , 
     n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , 
     n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , 
     n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , 
     n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , 
     n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , 
     n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , 
     n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , 
     n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , 
     n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , 
     n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , 
     n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , 
     n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , 
     n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , 
     n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , 
     n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , 
     n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , 
     n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , 
     n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , 
     n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , 
     n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , 
     n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , 
     n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , 
     n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , 
     n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , 
     n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , 
     n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , 
     n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , 
     n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , 
     n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , 
     n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , 
     n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , 
     n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , 
     n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , 
     n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , 
     n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , 
     n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , 
     n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , 
     n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , 
     n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , 
     n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , 
     n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , 
     n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , 
     n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , 
     n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , 
     n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , 
     n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , 
     n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , 
     n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , 
     n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , 
     n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , 
     n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , 
     n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , 
     n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , 
     n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , 
     n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , 
     n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , 
     n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , 
     n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , 
     n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , 
     n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , 
     n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , 
     n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , 
     n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , 
     n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , 
     n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , 
     n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , 
     n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , 
     n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , 
     n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , 
     n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , 
     n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , 
     n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , 
     n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , 
     n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , 
     n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , 
     n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , 
     n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , 
     n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , 
     n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , 
     n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , 
     n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , 
     n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , 
     n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , 
     n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , 
     n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , 
     n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , 
     n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , 
     n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , 
     n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , 
     n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , 
     n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , 
     n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , 
     n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , 
     n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , 
     n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , 
     n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , 
     n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , 
     n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , 
     n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , 
     n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , 
     n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , 
     n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , 
     n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , 
     n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , 
     n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , 
     n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , 
     n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , 
     n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , 
     n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , 
     n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , 
     n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , 
     n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , 
     n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , 
     n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , 
     n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , 
     n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , 
     n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , 
     n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , 
     n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , 
     n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , 
     n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , 
     n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , 
     n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , 
     n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , 
     n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , 
     n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , 
     n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , 
     n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , 
     n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , 
     n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , 
     n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , 
     n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , 
     n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , 
     n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , 
     n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , 
     n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , 
     n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , 
     n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , 
     n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , 
     n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , 
     n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , 
     n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , 
     n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , 
     n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , 
     n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , 
     n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , 
     n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , 
     n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , 
     n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , 
     n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , 
     n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , 
     n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , 
     n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , 
     n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , 
     n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , 
     n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , 
     n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , 
     n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , 
     n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , 
     n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , 
     n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , 
     n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , 
     n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , 
     n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , 
     n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , 
     n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , 
     n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , 
     n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , 
     n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , 
     n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , 
     n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , 
     n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , 
     n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , 
     n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , 
     n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , 
     n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , 
     n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , 
     n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , 
     n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , 
     n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , 
     n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , 
     n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , 
     n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , 
     n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , 
     n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , 
     n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , 
     n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , 
     n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , 
     n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , 
     n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , 
     n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , 
     n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , 
     n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , 
     n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , 
     n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , 
     n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , 
     n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , 
     n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , 
     n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , 
     n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , 
     n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , 
     n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , 
     n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , 
     n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , 
     n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , 
     n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , 
     n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , 
     n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , 
     n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , 
     n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , 
     n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , 
     n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , 
     n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , 
     n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , 
     n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , 
     n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , 
     n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , 
     n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , 
     n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , 
     n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , 
     n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , 
     n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , 
     n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , 
     n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , 
     n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , 
     n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , 
     n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , 
     n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , 
     n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , 
     n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , 
     n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , 
     n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , 
     n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , 
     n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , 
     n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , 
     n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , 
     n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , 
     n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , 
     n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , 
     n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , 
     n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , 
     n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , 
     n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , 
     n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , 
     n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , 
     n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , 
     n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , 
     n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , 
     n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , 
     n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , 
     n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , 
     n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , 
     n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , 
     n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , 
     n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , 
     n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , 
     n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , 
     n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , 
     n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , 
     n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , 
     n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , 
     n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , 
     n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , 
     n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , 
     n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , 
     n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , 
     n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , 
     n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , 
     n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , 
     n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , 
     n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , 
     n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , 
     n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , 
     n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , 
     n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , 
     n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , 
     n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , 
     n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , 
     n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , 
     n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , 
     n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , 
     n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , 
     n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , 
     n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , 
     n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , 
     n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , 
     n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , 
     n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , 
     n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , 
     n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , 
     n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , 
     n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , 
     n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , 
     n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , 
     n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , 
     n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , 
     n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , 
     n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , 
     n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , 
     n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , 
     n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , 
     n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , 
     n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , 
     n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , 
     n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , 
     n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , 
     n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , 
     n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , 
     n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , 
     n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , 
     n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , 
     n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , 
     n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , 
     n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , 
     n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , 
     n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , 
     n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , 
     n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , 
     n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , 
     n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , 
     n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , 
     n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , 
     n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , 
     n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , 
     n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , 
     n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , 
     n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , 
     n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , 
     n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , 
     n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , 
     n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , 
     n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , 
     n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , 
     n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , 
     n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , 
     n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , 
     n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , 
     n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , 
     n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , 
     n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , 
     n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , 
     n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , 
     n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , 
     n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , 
     n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , 
     n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , 
     n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , 
     n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , 
     n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , 
     n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , 
     n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , 
     n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , 
     n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , 
     n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , 
     n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , 
     n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , 
     n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , 
     n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , 
     n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , 
     n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , 
     n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , 
     n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , 
     n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , 
     n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , 
     n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , 
     n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , 
     n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , 
     n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , 
     n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , 
     n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , 
     n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , 
     n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , 
     n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , 
     n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , 
     n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , 
     n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , 
     n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , 
     n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , 
     n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , 
     n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , 
     n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , 
     n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , 
     n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , 
     n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , 
     n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , 
     n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , 
     n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , 
     n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , 
     n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , 
     n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , 
     n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , 
     n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , 
     n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , 
     n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , 
     n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , 
     n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , 
     n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , 
     n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , 
     n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , 
     n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , 
     n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , 
     n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , 
     n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , 
     n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , 
     n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , 
     n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , 
     n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , 
     n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , 
     n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , 
     n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , 
     n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , 
     n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , 
     n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , 
     n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , 
     n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , 
     n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , 
     n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , 
     n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , 
     n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , 
     n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , 
     n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , 
     n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , 
     n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , 
     n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , 
     n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , 
     n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , 
     n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , 
     n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , 
     n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , 
     n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , 
     n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , 
     n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , 
     n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , 
     n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , 
     n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , 
     n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , 
     n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , 
     n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , 
     n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , 
     n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , 
     n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , 
     n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , 
     n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , 
     n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , 
     n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , 
     n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , 
     n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , 
     n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , 
     n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , 
     n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , 
     n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , 
     n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , 
     n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , 
     n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , 
     n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , 
     n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , 
     n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , 
     n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , 
     n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , 
     n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , 
     n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , 
     n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , 
     n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , 
     n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , 
     n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , 
     n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , 
     n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , 
     n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , 
     n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , 
     n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , 
     n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , 
     n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , 
     n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , 
     n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , 
     n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , 
     n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , 
     n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , 
     n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , 
     n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , 
     n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , 
     n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , 
     n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , 
     n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , 
     n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , 
     n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , 
     n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , 
     n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , 
     n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , 
     n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , 
     n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , 
     n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , 
     n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , 
     n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , 
     n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , 
     n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , 
     n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , 
     n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , 
     n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , 
     n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , 
     n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , 
     n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , 
     n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , 
     n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , 
     n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , 
     n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , 
     n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , 
     n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , 
     n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , 
     n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , 
     n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , 
     n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , 
     n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , 
     n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , 
     n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , 
     n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , 
     n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , 
     n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , 
     n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , 
     n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , 
     n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , 
     n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , 
     n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , 
     n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , 
     n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , 
     n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , 
     n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , 
     n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , 
     n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , 
     n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , 
     n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , 
     n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , 
     n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , 
     n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , 
     n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , 
     n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , 
     n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , 
     n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , 
     n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , 
     n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , 
     n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , 
     n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , 
     n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , 
     n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , 
     n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , 
     n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , 
     n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , 
     n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , 
     n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , 
     n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , 
     n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , 
     n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , 
     n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , 
     n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , 
     n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , 
     n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , 
     n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , 
     n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , 
     n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , 
     n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , 
     n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , 
     n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , 
     n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , 
     n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , 
     n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , 
     n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , 
     n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , 
     n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , 
     n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , 
     n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , 
     n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , 
     n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , 
     n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , 
     n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , 
     n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , 
     n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , 
     n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , 
     n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , 
     n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , 
     n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , 
     n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , 
     n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , 
     n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , 
     n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , 
     n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , 
     n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , 
     n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , 
     n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , 
     n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , 
     n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , 
     n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , 
     n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , 
     n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , 
     n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , 
     n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , 
     n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , 
     n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , 
     n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , 
     n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , 
     n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , 
     n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , 
     n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , 
     n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , 
     n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , 
     n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , 
     n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , 
     n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , 
     n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , 
     n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , 
     n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , 
     n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , 
     n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , 
     n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , 
     n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , 
     n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , 
     n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , 
     n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , 
     n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , 
     n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , 
     n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , 
     n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , 
     n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , 
     n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , 
     n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , 
     n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , 
     n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , 
     n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , 
     n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , 
     n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , 
     n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , 
     n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , 
     n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , 
     n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , 
     n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , 
     n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , 
     n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , 
     n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , 
     n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , 
     n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , 
     n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , 
     n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , 
     n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , 
     n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , 
     n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , 
     n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , 
     n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , 
     n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , 
     n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , 
     n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , 
     n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , 
     n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , 
     n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , 
     n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , 
     n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , 
     n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , 
     n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , 
     n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , 
     n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , 
     n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , 
     n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , 
     n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , 
     n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , 
     n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , 
     n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , 
     n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , 
     n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , 
     n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , 
     n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , 
     n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , 
     n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , 
     n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , 
     n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , 
     n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , 
     n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , 
     n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , 
     n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , 
     n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , 
     n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , 
     n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , 
     n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , 
     n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , 
     n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , 
     n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , 
     n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , 
     n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , 
     n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , 
     n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , 
     n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , 
     n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , 
     n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , 
     n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , 
     n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , 
     n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , 
     n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , 
     n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , 
     n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , 
     n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , 
     n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , 
     n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , 
     n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , 
     n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , 
     n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , 
     n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , 
     n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , 
     n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , 
     n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , 
     n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , 
     n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , 
     n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , 
     n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , 
     n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , 
     n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , 
     n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , 
     n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , 
     n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , 
     n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , 
     n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , 
     n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , 
     n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , 
     n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , 
     n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , 
     n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , 
     n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , 
     n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , 
     n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , 
     n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , 
     n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , 
     n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , 
     n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , 
     n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , 
     n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , 
     n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , 
     n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , 
     n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , 
     n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , 
     n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , 
     n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , 
     n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , 
     n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , 
     n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , 
     n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , 
     n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , 
     n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , 
     n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , 
     n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , 
     n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , 
     n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , 
     n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , 
     n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , 
     n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , 
     n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , 
     n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , 
     n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , 
     n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , 
     n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , 
     n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , 
     n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , 
     n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , 
     n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , 
     n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , 
     n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , 
     n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , 
     n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , 
     n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , 
     n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , 
     n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , 
     n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , 
     n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , 
     n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , 
     n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , 
     n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , 
     n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , 
     n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , 
     n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , 
     n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , 
     n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , 
     n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , 
     n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , 
     n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , 
     n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , 
     n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , 
     n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , 
     n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , 
     n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , 
     n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , 
     n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , 
     n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , 
     n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , 
     n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , 
     n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , 
     n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , 
     n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , 
     n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , 
     n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , 
     n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , 
     n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , 
     n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , 
     n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , 
     n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , 
     n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , 
     n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , 
     n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , 
     n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , 
     n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , 
     n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , 
     n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , 
     n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , 
     n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , 
     n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , 
     n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , 
     n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , 
     n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , 
     n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , 
     n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , 
     n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , 
     n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , 
     n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , 
     n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , 
     n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , 
     n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , 
     n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , 
     n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , 
     n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , 
     n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , 
     n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , 
     n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , 
     n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , 
     n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , 
     n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , 
     n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , 
     n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , 
     n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , 
     n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , 
     n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , 
     n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , 
     n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , 
     n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , 
     n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , 
     n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , 
     n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , 
     n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , 
     n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , 
     n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , 
     n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , 
     n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , 
     n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , 
     n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , 
     n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , 
     n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , 
     n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , 
     n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , 
     n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , 
     n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , 
     n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , 
     n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , 
     n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , 
     n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , 
     n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , 
     n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , 
     n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , 
     n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , 
     n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , 
     n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , 
     n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , 
     n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , 
     n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , 
     n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , 
     n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , 
     n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , 
     n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , 
     n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , 
     n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , 
     n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , 
     n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , 
     n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , 
     n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , 
     n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , 
     n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , 
     n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , 
     n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , 
     n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , 
     n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , 
     n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , 
     n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , 
     n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , 
     n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , 
     n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , 
     n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , 
     n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , 
     n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , 
     n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , 
     n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , 
     n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , 
     n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , 
     n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , 
     n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , 
     n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , 
     n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , 
     n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , 
     n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , 
     n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , 
     n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , 
     n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , 
     n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , 
     n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , 
     n15411 , n15412 ;
buf ( n2187 , n9985 );
buf ( n2195 , n10744 );
buf ( n2192 , n12250 );
buf ( n2188 , n13433 );
buf ( n2190 , n13909 );
buf ( n2186 , n14368 );
buf ( n2191 , n14705 );
buf ( n2194 , n14946 );
buf ( n2193 , n15224 );
buf ( n2189 , n15412 );
buf ( n4394 , n1825 );
buf ( n4395 , n1584 );
buf ( n4396 , n1052 );
buf ( n4397 , n1350 );
buf ( n4398 , n746 );
buf ( n4399 , n1213 );
buf ( n4400 , n1132 );
buf ( n4401 , n420 );
buf ( n4402 , n85 );
buf ( n4403 , n1176 );
buf ( n4404 , n962 );
buf ( n4405 , n542 );
buf ( n4406 , n68 );
buf ( n4407 , n313 );
buf ( n4408 , n1070 );
buf ( n4409 , n719 );
buf ( n4410 , n980 );
buf ( n4411 , n251 );
buf ( n4412 , n295 );
buf ( n4413 , n1998 );
buf ( n4414 , n2091 );
buf ( n4415 , n733 );
buf ( n4416 , n678 );
buf ( n4417 , n13 );
buf ( n4418 , n2176 );
buf ( n4419 , n1534 );
buf ( n4420 , n1378 );
buf ( n4421 , n728 );
buf ( n4422 , n1100 );
buf ( n4423 , n1880 );
buf ( n4424 , n2152 );
buf ( n4425 , n1432 );
buf ( n4426 , n1708 );
buf ( n4427 , n135 );
buf ( n4428 , n2029 );
buf ( n4429 , n1431 );
buf ( n4430 , n1777 );
buf ( n4431 , n1757 );
buf ( n4432 , n1075 );
buf ( n4433 , n1450 );
buf ( n4434 , n455 );
buf ( n4435 , n266 );
buf ( n4436 , n1666 );
buf ( n4437 , n1412 );
buf ( n4438 , n859 );
buf ( n4439 , n548 );
buf ( n4440 , n1812 );
buf ( n4441 , n1937 );
buf ( n4442 , n1877 );
buf ( n4443 , n205 );
buf ( n4444 , n93 );
buf ( n4445 , n1460 );
buf ( n4446 , n370 );
buf ( n4447 , n1591 );
buf ( n4448 , n876 );
buf ( n4449 , n616 );
buf ( n4450 , n1603 );
buf ( n4451 , n682 );
buf ( n4452 , n288 );
buf ( n4453 , n2054 );
buf ( n4454 , n1376 );
buf ( n4455 , n1572 );
buf ( n4456 , n1047 );
buf ( n4457 , n139 );
buf ( n4458 , n901 );
buf ( n4459 , n764 );
buf ( n4460 , n1821 );
buf ( n4461 , n2130 );
buf ( n4462 , n908 );
buf ( n4463 , n587 );
buf ( n4464 , n187 );
buf ( n4465 , n75 );
buf ( n4466 , n924 );
buf ( n4467 , n2094 );
buf ( n4468 , n439 );
buf ( n4469 , n970 );
buf ( n4470 , n1272 );
buf ( n4471 , n1745 );
buf ( n4472 , n844 );
buf ( n4473 , n1719 );
buf ( n4474 , n430 );
buf ( n4475 , n1965 );
buf ( n4476 , n644 );
buf ( n4477 , n21 );
buf ( n4478 , n869 );
buf ( n4479 , n1927 );
buf ( n4480 , n1478 );
buf ( n4481 , n175 );
buf ( n4482 , n1867 );
buf ( n4483 , n1425 );
buf ( n4484 , n322 );
buf ( n4485 , n2083 );
buf ( n4486 , n1306 );
buf ( n4487 , n235 );
buf ( n4488 , n1638 );
buf ( n4489 , n1140 );
buf ( n4490 , n1333 );
buf ( n4491 , n1893 );
buf ( n4492 , n327 );
buf ( n4493 , n37 );
buf ( n4494 , n1182 );
buf ( n4495 , n1489 );
buf ( n4496 , n218 );
buf ( n4497 , n1314 );
buf ( n4498 , n372 );
buf ( n4499 , n656 );
buf ( n4500 , n1039 );
buf ( n4501 , n1889 );
buf ( n4502 , n1630 );
buf ( n4503 , n742 );
buf ( n4504 , n1096 );
buf ( n4505 , n181 );
buf ( n4506 , n1852 );
buf ( n4507 , n1801 );
buf ( n4508 , n811 );
buf ( n4509 , n2024 );
buf ( n4510 , n1293 );
buf ( n4511 , n243 );
buf ( n4512 , n630 );
buf ( n4513 , n515 );
buf ( n4514 , n131 );
buf ( n4515 , n735 );
buf ( n4516 , n423 );
buf ( n4517 , n2040 );
buf ( n4518 , n710 );
buf ( n4519 , n240 );
buf ( n4520 , n1267 );
buf ( n4521 , n592 );
buf ( n4522 , n2075 );
buf ( n4523 , n1384 );
buf ( n4524 , n722 );
buf ( n4525 , n1678 );
buf ( n4526 , n2071 );
buf ( n4527 , n957 );
buf ( n4528 , n76 );
buf ( n4529 , n1305 );
buf ( n4530 , n1410 );
buf ( n4531 , n1466 );
buf ( n4532 , n675 );
buf ( n4533 , n1448 );
buf ( n4534 , n98 );
buf ( n4535 , n1495 );
buf ( n4536 , n1086 );
buf ( n4537 , n1838 );
buf ( n4538 , n1308 );
buf ( n4539 , n407 );
buf ( n4540 , n711 );
buf ( n4541 , n726 );
buf ( n4542 , n2137 );
buf ( n4543 , n473 );
buf ( n4544 , n681 );
buf ( n4545 , n195 );
buf ( n4546 , n1637 );
buf ( n4547 , n427 );
buf ( n4548 , n1320 );
buf ( n4549 , n659 );
buf ( n4550 , n1659 );
buf ( n4551 , n263 );
buf ( n4552 , n586 );
buf ( n4553 , n43 );
buf ( n4554 , n461 );
buf ( n4555 , n2185 );
buf ( n4556 , n1715 );
buf ( n4557 , n2115 );
buf ( n4558 , n2148 );
buf ( n4559 , n1628 );
buf ( n4560 , n867 );
buf ( n4561 , n1179 );
buf ( n4562 , n578 );
buf ( n4563 , n1728 );
buf ( n4564 , n835 );
buf ( n4565 , n781 );
buf ( n4566 , n995 );
buf ( n4567 , n1536 );
buf ( n4568 , n484 );
buf ( n4569 , n1598 );
buf ( n4570 , n921 );
buf ( n4571 , n1918 );
buf ( n4572 , n519 );
buf ( n4573 , n415 );
buf ( n4574 , n1555 );
buf ( n4575 , n824 );
buf ( n4576 , n1463 );
buf ( n4577 , n1142 );
buf ( n4578 , n1675 );
buf ( n4579 , n1321 );
buf ( n4580 , n851 );
buf ( n4581 , n854 );
buf ( n4582 , n1740 );
buf ( n4583 , n1667 );
buf ( n4584 , n1133 );
buf ( n4585 , n1241 );
buf ( n4586 , n1519 );
buf ( n4587 , n2132 );
buf ( n4588 , n1170 );
buf ( n4589 , n353 );
buf ( n4590 , n1670 );
buf ( n4591 , n527 );
buf ( n4592 , n514 );
buf ( n4593 , n1967 );
buf ( n4594 , n513 );
buf ( n4595 , n1787 );
buf ( n4596 , n808 );
buf ( n4597 , n1741 );
buf ( n4598 , n716 );
buf ( n4599 , n2061 );
buf ( n4600 , n1917 );
buf ( n4601 , n308 );
buf ( n4602 , n123 );
buf ( n4603 , n17 );
buf ( n4604 , n1188 );
buf ( n4605 , n1767 );
buf ( n4606 , n137 );
buf ( n4607 , n701 );
buf ( n4608 , n1610 );
buf ( n4609 , n541 );
buf ( n4610 , n299 );
buf ( n4611 , n409 );
buf ( n4612 , n1077 );
buf ( n4613 , n516 );
buf ( n4614 , n1831 );
buf ( n4615 , n418 );
buf ( n4616 , n121 );
buf ( n4617 , n291 );
buf ( n4618 , n1749 );
buf ( n4619 , n2144 );
buf ( n4620 , n790 );
buf ( n4621 , n294 );
buf ( n4622 , n618 );
buf ( n4623 , n470 );
buf ( n4624 , n1229 );
buf ( n4625 , n853 );
buf ( n4626 , n2087 );
buf ( n4627 , n2039 );
buf ( n4628 , n890 );
buf ( n4629 , n1703 );
buf ( n4630 , n2033 );
buf ( n4631 , n1768 );
buf ( n4632 , n1313 );
buf ( n4633 , n302 );
buf ( n4634 , n1023 );
buf ( n4635 , n387 );
buf ( n4636 , n668 );
buf ( n4637 , n1428 );
buf ( n4638 , n1298 );
buf ( n4639 , n1566 );
buf ( n4640 , n483 );
buf ( n4641 , n2022 );
buf ( n4642 , n366 );
buf ( n4643 , n151 );
buf ( n4644 , n1562 );
buf ( n4645 , n1085 );
buf ( n4646 , n936 );
buf ( n4647 , n884 );
buf ( n4648 , n530 );
buf ( n4649 , n720 );
buf ( n4650 , n686 );
buf ( n4651 , n1351 );
buf ( n4652 , n2107 );
buf ( n4653 , n862 );
buf ( n4654 , n687 );
buf ( n4655 , n1597 );
buf ( n4656 , n42 );
buf ( n4657 , n1000 );
buf ( n4658 , n1158 );
buf ( n4659 , n1806 );
buf ( n4660 , n1149 );
buf ( n4661 , n989 );
buf ( n4662 , n1494 );
buf ( n4663 , n1307 );
buf ( n4664 , n2105 );
buf ( n4665 , n1058 );
buf ( n4666 , n839 );
buf ( n4667 , n310 );
buf ( n4668 , n1316 );
buf ( n4669 , n451 );
buf ( n4670 , n1884 );
buf ( n4671 , n880 );
buf ( n4672 , n1533 );
buf ( n4673 , n1003 );
buf ( n4674 , n1586 );
buf ( n4675 , n1035 );
buf ( n4676 , n1726 );
buf ( n4677 , n1711 );
buf ( n4678 , n624 );
buf ( n4679 , n805 );
buf ( n4680 , n569 );
buf ( n4681 , n1447 );
buf ( n4682 , n1166 );
buf ( n4683 , n614 );
buf ( n4684 , n55 );
buf ( n4685 , n1205 );
buf ( n4686 , n1248 );
buf ( n4687 , n1765 );
buf ( n4688 , n1512 );
buf ( n4689 , n1021 );
buf ( n4690 , n1727 );
buf ( n4691 , n1932 );
buf ( n4692 , n1007 );
buf ( n4693 , n1287 );
buf ( n4694 , n1413 );
buf ( n4695 , n1357 );
buf ( n4696 , n236 );
buf ( n4697 , n622 );
buf ( n4698 , n1582 );
buf ( n4699 , n1712 );
buf ( n4700 , n130 );
buf ( n4701 , n1243 );
buf ( n4702 , n1976 );
buf ( n4703 , n1090 );
buf ( n4704 , n388 );
buf ( n4705 , n964 );
buf ( n4706 , n1049 );
buf ( n4707 , n1850 );
buf ( n4708 , n1291 );
buf ( n4709 , n413 );
buf ( n4710 , n1441 );
buf ( n4711 , n1265 );
buf ( n4712 , n296 );
buf ( n4713 , n2066 );
buf ( n4714 , n1702 );
buf ( n4715 , n2182 );
buf ( n4716 , n1315 );
buf ( n4717 , n1554 );
buf ( n4718 , n341 );
buf ( n4719 , n1330 );
buf ( n4720 , n143 );
buf ( n4721 , n600 );
buf ( n4722 , n505 );
buf ( n4723 , n2150 );
buf ( n4724 , n1988 );
buf ( n4725 , n206 );
buf ( n4726 , n1289 );
buf ( n4727 , n1285 );
buf ( n4728 , n1589 );
buf ( n4729 , n1558 );
buf ( n4730 , n18 );
buf ( n4731 , n1946 );
buf ( n4732 , n1508 );
buf ( n4733 , n2073 );
buf ( n4734 , n1421 );
buf ( n4735 , n1110 );
buf ( n4736 , n1464 );
buf ( n4737 , n1046 );
buf ( n4738 , n99 );
buf ( n4739 , n1762 );
buf ( n4740 , n749 );
buf ( n4741 , n1802 );
buf ( n4742 , n1846 );
buf ( n4743 , n197 );
buf ( n4744 , n621 );
buf ( n4745 , n1922 );
buf ( n4746 , n159 );
buf ( n4747 , n1340 );
buf ( n4748 , n765 );
buf ( n4749 , n792 );
buf ( n4750 , n813 );
buf ( n4751 , n1861 );
buf ( n4752 , n886 );
buf ( n4753 , n1290 );
buf ( n4754 , n1575 );
buf ( n4755 , n499 );
buf ( n4756 , n545 );
buf ( n4757 , n665 );
buf ( n4758 , n1177 );
buf ( n4759 , n2168 );
buf ( n4760 , n1405 );
buf ( n4761 , n167 );
buf ( n4762 , n1948 );
buf ( n4763 , n1153 );
buf ( n4764 , n359 );
buf ( n4765 , n494 );
buf ( n4766 , n1300 );
buf ( n4767 , n628 );
buf ( n4768 , n1989 );
buf ( n4769 , n1012 );
buf ( n4770 , n588 );
buf ( n4771 , n1963 );
buf ( n4772 , n1004 );
buf ( n4773 , n1528 );
buf ( n4774 , n761 );
buf ( n4775 , n1337 );
buf ( n4776 , n31 );
buf ( n4777 , n250 );
buf ( n4778 , n1362 );
buf ( n4779 , n597 );
buf ( n4780 , n1420 );
buf ( n4781 , n814 );
buf ( n4782 , n1226 );
buf ( n4783 , n1548 );
buf ( n4784 , n392 );
buf ( n4785 , n400 );
buf ( n4786 , n504 );
buf ( n4787 , n2012 );
buf ( n4788 , n1601 );
buf ( n4789 , n657 );
buf ( n4790 , n399 );
buf ( n4791 , n1203 );
buf ( n4792 , n1266 );
buf ( n4793 , n1430 );
buf ( n4794 , n2076 );
buf ( n4795 , n1953 );
buf ( n4796 , n1234 );
buf ( n4797 , n257 );
buf ( n4798 , n2085 );
buf ( n4799 , n510 );
buf ( n4800 , n1923 );
buf ( n4801 , n2155 );
buf ( n4802 , n1629 );
buf ( n4803 , n39 );
buf ( n4804 , n830 );
buf ( n4805 , n1576 );
buf ( n4806 , n625 );
buf ( n4807 , n1418 );
buf ( n4808 , n1634 );
buf ( n4809 , n1855 );
buf ( n4810 , n1982 );
buf ( n4811 , n271 );
buf ( n4812 , n1286 );
buf ( n4813 , n396 );
buf ( n4814 , n405 );
buf ( n4815 , n1113 );
buf ( n4816 , n1843 );
buf ( n4817 , n672 );
buf ( n4818 , n2003 );
buf ( n4819 , n2088 );
buf ( n4820 , n317 );
buf ( n4821 , n727 );
buf ( n4822 , n603 );
buf ( n4823 , n1786 );
buf ( n4824 , n1688 );
buf ( n4825 , n67 );
buf ( n4826 , n2099 );
buf ( n4827 , n339 );
buf ( n4828 , n1553 );
buf ( n4829 , n180 );
buf ( n4830 , n1736 );
buf ( n4831 , n691 );
buf ( n4832 , n1792 );
buf ( n4833 , n1274 );
buf ( n4834 , n436 );
buf ( n4835 , n715 );
buf ( n4836 , n154 );
buf ( n4837 , n705 );
buf ( n4838 , n2042 );
buf ( n4839 , n1909 );
buf ( n4840 , n191 );
buf ( n4841 , n2001 );
buf ( n4842 , n1108 );
buf ( n4843 , n1006 );
buf ( n4844 , n589 );
buf ( n4845 , n1244 );
buf ( n4846 , n2013 );
buf ( n4847 , n369 );
buf ( n4848 , n2124 );
buf ( n4849 , n1636 );
buf ( n4850 , n1525 );
buf ( n4851 , n1198 );
buf ( n4852 , n4 );
buf ( n4853 , n1820 );
buf ( n4854 , n1644 );
buf ( n4855 , n583 );
buf ( n4856 , n356 );
buf ( n4857 , n1978 );
buf ( n4858 , n949 );
buf ( n4859 , n1024 );
buf ( n4860 , n1201 );
buf ( n4861 , n562 );
buf ( n4862 , n633 );
buf ( n4863 , n350 );
buf ( n4864 , n1643 );
buf ( n4865 , n651 );
buf ( n4866 , n882 );
buf ( n4867 , n2036 );
buf ( n4868 , n397 );
buf ( n4869 , n2175 );
buf ( n4870 , n15 );
buf ( n4871 , n390 );
buf ( n4872 , n897 );
buf ( n4873 , n1277 );
buf ( n4874 , n971 );
buf ( n4875 , n3 );
buf ( n4876 , n1185 );
buf ( n4877 , n1853 );
buf ( n4878 , n2134 );
buf ( n4879 , n1841 );
buf ( n4880 , n54 );
buf ( n4881 , n769 );
buf ( n4882 , n1474 );
buf ( n4883 , n1327 );
buf ( n4884 , n332 );
buf ( n4885 , n690 );
buf ( n4886 , n1453 );
buf ( n4887 , n2139 );
buf ( n4888 , n368 );
buf ( n4889 , n2110 );
buf ( n4890 , n2121 );
buf ( n4891 , n645 );
buf ( n4892 , n1294 );
buf ( n4893 , n1936 );
buf ( n4894 , n211 );
buf ( n4895 , n1099 );
buf ( n4896 , n1763 );
buf ( n4897 , n785 );
buf ( n4898 , n108 );
buf ( n4899 , n703 );
buf ( n4900 , n1310 );
buf ( n4901 , n1399 );
buf ( n4902 , n1184 );
buf ( n4903 , n609 );
buf ( n4904 , n275 );
buf ( n4905 , n1619 );
buf ( n4906 , n1117 );
buf ( n4907 , n903 );
buf ( n4908 , n1839 );
buf ( n4909 , n907 );
buf ( n4910 , n1128 );
buf ( n4911 , n926 );
buf ( n4912 , n1623 );
buf ( n4913 , n1939 );
buf ( n4914 , n1661 );
buf ( n4915 , n10 );
buf ( n4916 , n462 );
buf ( n4917 , n1393 );
buf ( n4918 , n1774 );
buf ( n4919 , n2177 );
buf ( n4920 , n525 );
buf ( n4921 , n756 );
buf ( n4922 , n343 );
buf ( n4923 , n28 );
buf ( n4924 , n1124 );
buf ( n4925 , n1523 );
buf ( n4926 , n1772 );
buf ( n4927 , n2170 );
buf ( n4928 , n1750 );
buf ( n4929 , n1050 );
buf ( n4930 , n596 );
buf ( n4931 , n741 );
buf ( n4932 , n344 );
buf ( n4933 , n1960 );
buf ( n4934 , n1088 );
buf ( n4935 , n1183 );
buf ( n4936 , n1511 );
buf ( n4937 , n1779 );
buf ( n4938 , n1089 );
buf ( n4939 , n655 );
buf ( n4940 , n2045 );
buf ( n4941 , n573 );
buf ( n4942 , n1473 );
buf ( n4943 , n736 );
buf ( n4944 , n1349 );
buf ( n4945 , n2055 );
buf ( n4946 , n977 );
buf ( n4947 , n1613 );
buf ( n4948 , n920 );
buf ( n4949 , n311 );
buf ( n4950 , n414 );
buf ( n4951 , n1235 );
buf ( n4952 , n1156 );
buf ( n4953 , n1367 );
buf ( n4954 , n684 );
buf ( n4955 , n1181 );
buf ( n4956 , n33 );
buf ( n4957 , n2147 );
buf ( n4958 , n885 );
buf ( n4959 , n112 );
buf ( n4960 , n658 );
buf ( n4961 , n721 );
buf ( n4962 , n918 );
buf ( n4963 , n373 );
buf ( n4964 , n1284 );
buf ( n4965 , n531 );
buf ( n4966 , n2097 );
buf ( n4967 , n283 );
buf ( n4968 , n739 );
buf ( n4969 , n1723 );
buf ( n4970 , n1172 );
buf ( n4971 , n1627 );
buf ( n4972 , n1251 );
buf ( n4973 , n2031 );
buf ( n4974 , n1196 );
buf ( n4975 , n606 );
buf ( n4976 , n836 );
buf ( n4977 , n988 );
buf ( n4978 , n2002 );
buf ( n4979 , n996 );
buf ( n4980 , n393 );
buf ( n4981 , n2164 );
buf ( n4982 , n2172 );
buf ( n4983 , n491 );
buf ( n4984 , n745 );
buf ( n4985 , n1498 );
buf ( n4986 , n928 );
buf ( n4987 , n1390 );
buf ( n4988 , n1514 );
buf ( n4989 , n265 );
buf ( n4990 , n454 );
buf ( n4991 , n1220 );
buf ( n4992 , n899 );
buf ( n4993 , n300 );
buf ( n4994 , n227 );
buf ( n4995 , n2092 );
buf ( n4996 , n1633 );
buf ( n4997 , n750 );
buf ( n4998 , n245 );
buf ( n4999 , n1782 );
buf ( n5000 , n930 );
buf ( n5001 , n2116 );
buf ( n5002 , n1747 );
buf ( n5003 , n772 );
buf ( n5004 , n538 );
buf ( n5005 , n1987 );
buf ( n5006 , n26 );
buf ( n5007 , n917 );
buf ( n5008 , n1479 );
buf ( n5009 , n643 );
buf ( n5010 , n789 );
buf ( n5011 , n1858 );
buf ( n5012 , n1370 );
buf ( n5013 , n1535 );
buf ( n5014 , n87 );
buf ( n5015 , n156 );
buf ( n5016 , n1397 );
buf ( n5017 , n1790 );
buf ( n5018 , n342 );
buf ( n5019 , n837 );
buf ( n5020 , n446 );
buf ( n5021 , n1914 );
buf ( n5022 , n1452 );
buf ( n5023 , n1232 );
buf ( n5024 , n161 );
buf ( n5025 , n1053 );
buf ( n5026 , n186 );
buf ( n5027 , n304 );
buf ( n5028 , n779 );
buf ( n5029 , n2023 );
buf ( n5030 , n239 );
buf ( n5031 , n258 );
buf ( n5032 , n1257 );
buf ( n5033 , n2010 );
buf ( n5034 , n340 );
buf ( n5035 , n432 );
buf ( n5036 , n693 );
buf ( n5037 , n1130 );
buf ( n5038 , n558 );
buf ( n5039 , n636 );
buf ( n5040 , n2006 );
buf ( n5041 , n1022 );
buf ( n5042 , n1301 );
buf ( n5043 , n1374 );
buf ( n5044 , n1904 );
buf ( n5045 , n1549 );
buf ( n5046 , n226 );
buf ( n5047 , n5 );
buf ( n5048 , n489 );
buf ( n5049 , n685 );
buf ( n5050 , n394 );
buf ( n5051 , n1326 );
buf ( n5052 , n249 );
buf ( n5053 , n916 );
buf ( n5054 , n65 );
buf ( n5055 , n1694 );
buf ( n5056 , n314 );
buf ( n5057 , n1335 );
buf ( n5058 , n1336 );
buf ( n5059 , n1258 );
buf ( n5060 , n1093 );
buf ( n5061 , n570 );
buf ( n5062 , n1766 );
buf ( n5063 , n1458 );
buf ( n5064 , n1137 );
buf ( n5065 , n817 );
buf ( n5066 , n581 );
buf ( n5067 , n911 );
buf ( n5068 , n2070 );
buf ( n5069 , n563 );
buf ( n5070 , n820 );
buf ( n5071 , n941 );
buf ( n5072 , n1202 );
buf ( n5073 , n80 );
buf ( n5074 , n708 );
buf ( n5075 , n1513 );
buf ( n5076 , n367 );
buf ( n5077 , n416 );
buf ( n5078 , n162 );
buf ( n5079 , n1119 );
buf ( n5080 , n555 );
buf ( n5081 , n648 );
buf ( n5082 , n860 );
buf ( n5083 , n334 );
buf ( n5084 , n165 );
buf ( n5085 , n838 );
buf ( n5086 , n1173 );
buf ( n5087 , n1187 );
buf ( n5088 , n1488 );
buf ( n5089 , n307 );
buf ( n5090 , n1552 );
buf ( n5091 , n1828 );
buf ( n5092 , n892 );
buf ( n5093 , n1868 );
buf ( n5094 , n1219 );
buf ( n5095 , n2142 );
buf ( n5096 , n8 );
buf ( n5097 , n371 );
buf ( n5098 , n153 );
buf ( n5099 , n1123 );
buf ( n5100 , n1343 );
buf ( n5101 , n1994 );
buf ( n5102 , n1738 );
buf ( n5103 , n0 );
buf ( n5104 , n1255 );
buf ( n5105 , n463 );
buf ( n5106 , n612 );
buf ( n5107 , n1118 );
buf ( n5108 , n200 );
buf ( n5109 , n301 );
buf ( n5110 , n476 );
buf ( n5111 , n1168 );
buf ( n5112 , n244 );
buf ( n5113 , n1876 );
buf ( n5114 , n138 );
buf ( n5115 , n1700 );
buf ( n5116 , n1484 );
buf ( n5117 , n1217 );
buf ( n5118 , n883 );
buf ( n5119 , n401 );
buf ( n5120 , n1863 );
buf ( n5121 , n896 );
buf ( n5122 , n149 );
buf ( n5123 , n1596 );
buf ( n5124 , n1592 );
buf ( n5125 , n652 );
buf ( n5126 , n352 );
buf ( n5127 , n203 );
buf ( n5128 , n744 );
buf ( n5129 , n986 );
buf ( n5130 , n1121 );
buf ( n5131 , n1773 );
buf ( n5132 , n966 );
buf ( n5133 , n386 );
buf ( n5134 , n2145 );
buf ( n5135 , n582 );
buf ( n5136 , n1721 );
buf ( n5137 , n1455 );
buf ( n5138 , n1561 );
buf ( n5139 , n747 );
buf ( n5140 , n475 );
buf ( n5141 , n142 );
buf ( n5142 , n1568 );
buf ( n5143 , n1073 );
buf ( n5144 , n2112 );
buf ( n5145 , n2044 );
buf ( n5146 , n2181 );
buf ( n5147 , n176 );
buf ( n5148 , n1483 );
buf ( n5149 , n492 );
buf ( n5150 , n83 );
buf ( n5151 , n1268 );
buf ( n5152 , n472 );
buf ( n5153 , n723 );
buf ( n5154 , n613 );
buf ( n5155 , n101 );
buf ( n5156 , n1769 );
buf ( n5157 , n1363 );
buf ( n5158 , n554 );
buf ( n5159 , n1192 );
buf ( n5160 , n1709 );
buf ( n5161 , n1152 );
buf ( n5162 , n450 );
buf ( n5163 , n1583 );
buf ( n5164 , n1364 );
buf ( n5165 , n1911 );
buf ( n5166 , n459 );
buf ( n5167 , n2106 );
buf ( n5168 , n242 );
buf ( n5169 , n1887 );
buf ( n5170 , n169 );
buf ( n5171 , n1794 );
buf ( n5172 , n654 );
buf ( n5173 , n469 );
buf ( n5174 , n823 );
buf ( n5175 , n1710 );
buf ( n5176 , n788 );
buf ( n5177 , n1467 );
buf ( n5178 , n889 );
buf ( n5179 , n1279 );
buf ( n5180 , n1873 );
buf ( n5181 , n782 );
buf ( n5182 , n1764 );
buf ( n5183 , n1866 );
buf ( n5184 , n1197 );
buf ( n5185 , n1107 );
buf ( n5186 , n1574 );
buf ( n5187 , n1459 );
buf ( n5188 , n848 );
buf ( n5189 , n1322 );
buf ( n5190 , n841 );
buf ( n5191 , n768 );
buf ( n5192 , n1296 );
buf ( n5193 , n365 );
buf ( n5194 , n653 );
buf ( n5195 , n428 );
buf ( n5196 , n1865 );
buf ( n5197 , n1369 );
buf ( n5198 , n2032 );
buf ( n5199 , n133 );
buf ( n5200 , n1814 );
buf ( n5201 , n1817 );
buf ( n5202 , n2133 );
buf ( n5203 , n972 );
buf ( n5204 , n1943 );
buf ( n5205 , n1888 );
buf ( n5206 , n1423 );
buf ( n5207 , n757 );
buf ( n5208 , n480 );
buf ( n5209 , n937 );
buf ( n5210 , n1354 );
buf ( n5211 , n1446 );
buf ( n5212 , n1 );
buf ( n5213 , n919 );
buf ( n5214 , n679 );
buf ( n5215 , n113 );
buf ( n5216 , n1395 );
buf ( n5217 , n1391 );
buf ( n5218 , n2065 );
buf ( n5219 , n1078 );
buf ( n5220 , n1245 );
buf ( n5221 , n117 );
buf ( n5222 , n1571 );
buf ( n5223 , n1684 );
buf ( n5224 , n424 );
buf ( n5225 , n1016 );
buf ( n5226 , n1730 );
buf ( n5227 , n1465 );
buf ( n5228 , n2005 );
buf ( n5229 , n791 );
buf ( n5230 , n994 );
buf ( n5231 , n417 );
buf ( n5232 , n1557 );
buf ( n5233 , n536 );
buf ( n5234 , n947 );
buf ( n5235 , n696 );
buf ( n5236 , n755 );
buf ( n5237 , n1499 );
buf ( n5238 , n1756 );
buf ( n5239 , n1328 );
buf ( n5240 , n1338 );
buf ( n5241 , n496 );
buf ( n5242 , n282 );
buf ( n5243 , n1486 );
buf ( n5244 , n1503 );
buf ( n5245 , n2162 );
buf ( n5246 , n1869 );
buf ( n5247 , n1444 );
buf ( n5248 , n1303 );
buf ( n5249 , n700 );
buf ( n5250 , n992 );
buf ( n5251 , n1160 );
buf ( n5252 , n1585 );
buf ( n5253 , n238 );
buf ( n5254 , n11 );
buf ( n5255 , n1951 );
buf ( n5256 , n2016 );
buf ( n5257 , n349 );
buf ( n5258 , n1950 );
buf ( n5259 , n895 );
buf ( n5260 , n1577 );
buf ( n5261 , n1416 );
buf ( n5262 , n1388 );
buf ( n5263 , n929 );
buf ( n5264 , n1018 );
buf ( n5265 , n106 );
buf ( n5266 , n1346 );
buf ( n5267 , n1231 );
buf ( n5268 , n758 );
buf ( n5269 , n448 );
buf ( n5270 , n1510 );
buf ( n5271 , n213 );
buf ( n5272 , n443 );
buf ( n5273 , n1655 );
buf ( n5274 , n1036 );
buf ( n5275 , n751 );
buf ( n5276 , n1674 );
buf ( n5277 , n1811 );
buf ( n5278 , n1208 );
buf ( n5279 , n1230 );
buf ( n5280 , n601 );
buf ( n5281 , n697 );
buf ( n5282 , n1045 );
buf ( n5283 , n1332 );
buf ( n5284 , n29 );
buf ( n5285 , n997 );
buf ( n5286 , n1797 );
buf ( n5287 , n1031 );
buf ( n5288 , n1681 );
buf ( n5289 , n171 );
buf ( n5290 , n2146 );
buf ( n5291 , n894 );
buf ( n5292 , n207 );
buf ( n5293 , n223 );
buf ( n5294 , n1539 );
buf ( n5295 , n840 );
buf ( n5296 , n1968 );
buf ( n5297 , n224 );
buf ( n5298 , n978 );
buf ( n5299 , n1938 );
buf ( n5300 , n1680 );
buf ( n5301 , n1966 );
buf ( n5302 , n210 );
buf ( n5303 , n498 );
buf ( n5304 , n351 );
buf ( n5305 , n676 );
buf ( n5306 , n406 );
buf ( n5307 , n194 );
buf ( n5308 , n1347 );
buf ( n5309 , n1457 );
buf ( n5310 , n437 );
buf ( n5311 , n855 );
buf ( n5312 , n752 );
buf ( n5313 , n1622 );
buf ( n5314 , n19 );
buf ( n5315 , n1614 );
buf ( n5316 , n961 );
buf ( n5317 , n260 );
buf ( n5318 , n1072 );
buf ( n5319 , n1040 );
buf ( n5320 , n1141 );
buf ( n5321 , n1426 );
buf ( n5322 , n1057 );
buf ( n5323 , n2159 );
buf ( n5324 , n95 );
buf ( n5325 , n114 );
buf ( n5326 , n1477 );
buf ( n5327 , n1106 );
buf ( n5328 , n466 );
buf ( n5329 , n783 );
buf ( n5330 , n1263 );
buf ( n5331 , n255 );
buf ( n5332 , n46 );
buf ( n5333 , n1945 );
buf ( n5334 , n1706 );
buf ( n5335 , n20 );
buf ( n5336 , n585 );
buf ( n5337 , n259 );
buf ( n5338 , n477 );
buf ( n5339 , n64 );
buf ( n5340 , n269 );
buf ( n5341 , n1329 );
buf ( n5342 , n1081 );
buf ( n5343 , n1944 );
buf ( n5344 , n1605 );
buf ( n5345 , n1309 );
buf ( n5346 , n2038 );
buf ( n5347 , n1974 );
buf ( n5348 , n1758 );
buf ( n5349 , n1908 );
buf ( n5350 , n1456 );
buf ( n5351 , n1295 );
buf ( n5352 , n1240 );
buf ( n5353 , n1720 );
buf ( n5354 , n1990 );
buf ( n5355 , n464 );
buf ( n5356 , n2120 );
buf ( n5357 , n1207 );
buf ( n5358 , n599 );
buf ( n5359 , n533 );
buf ( n5360 , n802 );
buf ( n5361 , n1092 );
buf ( n5362 , n1879 );
buf ( n5363 , n584 );
buf ( n5364 , n780 );
buf ( n5365 , n1299 );
buf ( n5366 , n1631 );
buf ( n5367 , n952 );
buf ( n5368 , n1564 );
buf ( n5369 , n1414 );
buf ( n5370 , n361 );
buf ( n5371 , n1729 );
buf ( n5372 , n1451 );
buf ( n5373 , n831 );
buf ( n5374 , n660 );
buf ( n5375 , n826 );
buf ( n5376 , n2020 );
buf ( n5377 , n922 );
buf ( n5378 , n1754 );
buf ( n5379 , n1515 );
buf ( n5380 , n1317 );
buf ( n5381 , n2127 );
buf ( n5382 , n118 );
buf ( n5383 , n1030 );
buf ( n5384 , n440 );
buf ( n5385 , n1250 );
buf ( n5386 , n979 );
buf ( n5387 , n1001 );
buf ( n5388 , n640 );
buf ( n5389 , n1135 );
buf ( n5390 , n821 );
buf ( n5391 , n550 );
buf ( n5392 , n189 );
buf ( n5393 , n1237 );
buf ( n5394 , n453 );
buf ( n5395 , n1928 );
buf ( n5396 , n873 );
buf ( n5397 , n1606 );
buf ( n5398 , n794 );
buf ( n5399 , n888 );
buf ( n5400 , n1621 );
buf ( n5401 , n385 );
buf ( n5402 , n1983 );
buf ( n5403 , n1902 );
buf ( n5404 , n1212 );
buf ( n5405 , n184 );
buf ( n5406 , n102 );
buf ( n5407 , n422 );
buf ( n5408 , n1407 );
buf ( n5409 , n285 );
buf ( n5410 , n1952 );
buf ( n5411 , n1429 );
buf ( n5412 , n1827 );
buf ( n5413 , n712 );
buf ( n5414 , n674 );
buf ( n5415 , n912 );
buf ( n5416 , n875 );
buf ( n5417 , n887 );
buf ( n5418 , n1929 );
buf ( n5419 , n278 );
buf ( n5420 , n1408 );
buf ( n5421 , n1481 );
buf ( n5422 , n1496 );
buf ( n5423 , n246 );
buf ( n5424 , n2119 );
buf ( n5425 , n1999 );
buf ( n5426 , n2117 );
buf ( n5427 , n338 );
buf ( n5428 , n1699 );
buf ( n5429 , n2135 );
buf ( n5430 , n1755 );
buf ( n5431 , n1358 );
buf ( n5432 , n287 );
buf ( n5433 , n2050 );
buf ( n5434 , n1312 );
buf ( n5435 , n1716 );
buf ( n5436 , n1587 );
buf ( n5437 , n1246 );
buf ( n5438 , n1249 );
buf ( n5439 , n384 );
buf ( n5440 , n1262 );
buf ( n5441 , n408 );
buf ( n5442 , n680 );
buf ( n5443 , n2174 );
buf ( n5444 , n1051 );
buf ( n5445 , n2118 );
buf ( n5446 , n1803 );
buf ( n5447 , n560 );
buf ( n5448 , n1278 );
buf ( n5449 , n1344 );
buf ( n5450 , n1996 );
buf ( n5451 , n2053 );
buf ( n5452 , n1878 );
buf ( n5453 , n999 );
buf ( n5454 , n1651 );
buf ( n5455 , n374 );
buf ( n5456 , n1903 );
buf ( n5457 , n946 );
buf ( n5458 , n395 );
buf ( n5459 , n1013 );
buf ( n5460 , n286 );
buf ( n5461 , n872 );
buf ( n5462 , n1043 );
buf ( n5463 , n1546 );
buf ( n5464 , n1506 );
buf ( n5465 , n934 );
buf ( n5466 , n2101 );
buf ( n5467 , n1403 );
buf ( n5468 , n1912 );
buf ( n5469 , n730 );
buf ( n5470 , n567 );
buf ( n5471 , n1832 );
buf ( n5472 , n150 );
buf ( n5473 , n702 );
buf ( n5474 , n1609 );
buf ( n5475 , n276 );
buf ( n5476 , n1462 );
buf ( n5477 , n232 );
buf ( n5478 , n62 );
buf ( n5479 , n1657 );
buf ( n5480 , n215 );
buf ( n5481 , n1521 );
buf ( n5482 , n48 );
buf ( n5483 , n798 );
buf ( n5484 , n71 );
buf ( n5485 , n1771 );
buf ( n5486 , n1044 );
buf ( n5487 , n965 );
buf ( n5488 , n1224 );
buf ( n5489 , n1886 );
buf ( n5490 , n1526 );
buf ( n5491 , n1835 );
buf ( n5492 , n553 );
buf ( n5493 , n650 );
buf ( n5494 , n1162 );
buf ( n5495 , n2184 );
buf ( n5496 , n160 );
buf ( n5497 , n1848 );
buf ( n5498 , n991 );
buf ( n5499 , n1784 );
buf ( n5500 , n360 );
buf ( n5501 , n281 );
buf ( n5502 , n1981 );
buf ( n5503 , n1063 );
buf ( n5504 , n1804 );
buf ( n5505 , n1897 );
buf ( n5506 , n219 );
buf ( n5507 , n1696 );
buf ( n5508 , n1150 );
buf ( n5509 , n140 );
buf ( n5510 , n506 );
buf ( n5511 , n1002 );
buf ( n5512 , n481 );
buf ( n5513 , n445 );
buf ( n5514 , n319 );
buf ( n5515 , n974 );
buf ( n5516 , n92 );
buf ( n5517 , n635 );
buf ( n5518 , n1037 );
buf ( n5519 , n1578 );
buf ( n5520 , n1180 );
buf ( n5521 , n1143 );
buf ( n5522 , n482 );
buf ( n5523 , n900 );
buf ( n5524 , n767 );
buf ( n5525 , n1664 );
buf ( n5526 , n144 );
buf ( n5527 , n60 );
buf ( n5528 , n69 );
buf ( n5529 , n2096 );
buf ( n5530 , n1611 );
buf ( n5531 , n677 );
buf ( n5532 , n1079 );
buf ( n5533 , n1288 );
buf ( n5534 , n345 );
buf ( n5535 , n40 );
buf ( n5536 , n2156 );
buf ( n5537 , n228 );
buf ( n5538 , n833 );
buf ( n5539 , n1163 );
buf ( n5540 , n297 );
buf ( n5541 , n664 );
buf ( n5542 , n192 );
buf ( n5543 , n50 );
buf ( n5544 , n1147 );
buf ( n5545 , n2047 );
buf ( n5546 , n254 );
buf ( n5547 , n923 );
buf ( n5548 , n1958 );
buf ( n5549 , n623 );
buf ( n5550 , n27 );
buf ( n5551 , n104 );
buf ( n5552 , n523 );
buf ( n5553 , n927 );
buf ( n5554 , n1672 );
buf ( n5555 , n438 );
buf ( n5556 , n718 );
buf ( n5557 , n500 );
buf ( n5558 , n766 );
buf ( n5559 , n1104 );
buf ( n5560 , n552 );
buf ( n5561 , n1472 );
buf ( n5562 , n1746 );
buf ( n5563 , n1642 );
buf ( n5564 , n1435 );
buf ( n5565 , n1253 );
buf ( n5566 , n2161 );
buf ( n5567 , n1824 );
buf ( n5568 , n1926 );
buf ( n5569 , n1891 );
buf ( n5570 , n905 );
buf ( n5571 , n1901 );
buf ( n5572 , n2122 );
buf ( n5573 , n1516 );
buf ( n5574 , n2166 );
buf ( n5575 , n1870 );
buf ( n5576 , n429 );
buf ( n5577 , n379 );
buf ( n5578 , n465 );
buf ( n5579 , n933 );
buf ( n5580 , n1693 );
buf ( n5581 , n1930 );
buf ( n5582 , n1146 );
buf ( n5583 , n1341 );
buf ( n5584 , n1404 );
buf ( n5585 , n2058 );
buf ( n5586 , n1134 );
buf ( n5587 , n274 );
buf ( n5588 , n898 );
buf ( n5589 , n1658 );
buf ( n5590 , n1084 );
buf ( n5591 , n25 );
buf ( n5592 , n717 );
buf ( n5593 , n1076 );
buf ( n5594 , n816 );
buf ( n5595 , n732 );
buf ( n5596 , n1256 );
buf ( n5597 , n669 );
buf ( n5598 , n471 );
buf ( n5599 , n595 );
buf ( n5600 , n1669 );
buf ( n5601 , n1713 );
buf ( n5602 , n1190 );
buf ( n5603 , n212 );
buf ( n5604 , n1618 );
buf ( n5605 , n576 );
buf ( n5606 , n1480 );
buf ( n5607 , n1214 );
buf ( n5608 , n1984 );
buf ( n5609 , n753 );
buf ( n5610 , n1379 );
buf ( n5611 , n1238 );
buf ( n5612 , n1437 );
buf ( n5613 , n174 );
buf ( n5614 , n1890 );
buf ( n5615 , n535 );
buf ( n5616 , n136 );
buf ( n5617 , n2163 );
buf ( n5618 , n177 );
buf ( n5619 , n1579 );
buf ( n5620 , n1973 );
buf ( n5621 , n709 );
buf ( n5622 , n1417 );
buf ( n5623 , n1394 );
buf ( n5624 , n692 );
buf ( n5625 , n1154 );
buf ( n5626 , n1373 );
buf ( n5627 , n479 );
buf ( n5628 , n1676 );
buf ( n5629 , n1954 );
buf ( n5630 , n202 );
buf ( n5631 , n1471 );
buf ( n5632 , n1685 );
buf ( n5633 , n842 );
buf ( n5634 , n1590 );
buf ( n5635 , n1748 );
buf ( n5636 , n1259 );
buf ( n5637 , n458 );
buf ( n5638 , n981 );
buf ( n5639 , n1461 );
buf ( n5640 , n2151 );
buf ( n5641 , n557 );
buf ( n5642 , n843 );
buf ( n5643 , n893 );
buf ( n5644 , n748 );
buf ( n5645 , n431 );
buf ( n5646 , n145 );
buf ( n5647 , n1550 );
buf ( n5648 , n2100 );
buf ( n5649 , n88 );
buf ( n5650 , n1324 );
buf ( n5651 , n2046 );
buf ( n5652 , n2077 );
buf ( n5653 , n1325 );
buf ( n5654 , n293 );
buf ( n5655 , n1705 );
buf ( n5656 , n1476 );
buf ( n5657 , n2138 );
buf ( n5658 , n2141 );
buf ( n5659 , n488 );
buf ( n5660 , n1485 );
buf ( n5661 , n1737 );
buf ( n5662 , n2149 );
buf ( n5663 , n615 );
buf ( n5664 , n1080 );
buf ( n5665 , n1872 );
buf ( n5666 , n925 );
buf ( n5667 , n762 );
buf ( n5668 , n631 );
buf ( n5669 , n2179 );
buf ( n5670 , n1805 );
buf ( n5671 , n626 );
buf ( n5672 , n51 );
buf ( n5673 , n1385 );
buf ( n5674 , n738 );
buf ( n5675 , n1221 );
buf ( n5676 , n1302 );
buf ( n5677 , n115 );
buf ( n5678 , n2143 );
buf ( n5679 , n412 );
buf ( n5680 , n507 );
buf ( n5681 , n1164 );
buf ( n5682 , n1282 );
buf ( n5683 , n94 );
buf ( n5684 , n1862 );
buf ( n5685 , n607 );
buf ( n5686 , n521 );
buf ( n5687 , n1541 );
buf ( n5688 , n1647 );
buf ( n5689 , n1438 );
buf ( n5690 , n1895 );
buf ( n5691 , n641 );
buf ( n5692 , n604 );
buf ( n5693 , n673 );
buf ( n5694 , n1334 );
buf ( n5695 , n1735 );
buf ( n5696 , n1751 );
buf ( n5697 , n629 );
buf ( n5698 , n1034 );
buf ( n5699 , n1439 );
buf ( n5700 , n1522 );
buf ( n5701 , n273 );
buf ( n5702 , n1167 );
buf ( n5703 , n1972 );
buf ( n5704 , n444 );
buf ( n5705 , n1011 );
buf ( n5706 , n280 );
buf ( n5707 , n323 );
buf ( n5708 , n59 );
buf ( n5709 , n2111 );
buf ( n5710 , n1283 );
buf ( n5711 , n256 );
buf ( n5712 , n326 );
buf ( n5713 , n829 );
buf ( n5714 , n1789 );
buf ( n5715 , n1353 );
buf ( n5716 , n857 );
buf ( n5717 , n1816 );
buf ( n5718 , n2049 );
buf ( n5719 , n610 );
buf ( n5720 , n1701 );
buf ( n5721 , n847 );
buf ( n5722 , n1612 );
buf ( n5723 , n493 );
buf ( n5724 , n1645 );
buf ( n5725 , n1991 );
buf ( n5726 , n1704 );
buf ( n5727 , n1743 );
buf ( n5728 , n2067 );
buf ( n5729 , n619 );
buf ( n5730 , n874 );
buf ( n5731 , n976 );
buf ( n5732 , n1906 );
buf ( n5733 , n2014 );
buf ( n5734 , n328 );
buf ( n5735 , n1355 );
buf ( n5736 , n942 );
buf ( n5737 , n1993 );
buf ( n5738 , n1010 );
buf ( n5739 , n540 );
buf ( n5740 , n23 );
buf ( n5741 , n948 );
buf ( n5742 , n1380 );
buf ( n5743 , n1776 );
buf ( n5744 , n1372 );
buf ( n5745 , n148 );
buf ( n5746 , n819 );
buf ( n5747 , n511 );
buf ( n5748 , n6 );
buf ( n5749 , n526 );
buf ( n5750 , n1433 );
buf ( n5751 , n803 );
buf ( n5752 , n1697 );
buf ( n5753 , n773 );
buf ( n5754 , n503 );
buf ( n5755 , n1781 );
buf ( n5756 , n1098 );
buf ( n5757 , n1112 );
buf ( n5758 , n1138 );
buf ( n5759 , n1199 );
buf ( n5760 , n1157 );
buf ( n5761 , n456 );
buf ( n5762 , n944 );
buf ( n5763 , n754 );
buf ( n5764 , n247 );
buf ( n5765 , n985 );
buf ( n5766 , n982 );
buf ( n5767 , n666 );
buf ( n5768 , n1588 );
buf ( n5769 , n760 );
buf ( n5770 , n574 );
buf ( n5771 , n58 );
buf ( n5772 , n534 );
buf ( n5773 , n2034 );
buf ( n5774 , n2008 );
buf ( n5775 , n529 );
buf ( n5776 , n1992 );
buf ( n5777 , n163 );
buf ( n5778 , n134 );
buf ( n5779 , n868 );
buf ( n5780 , n1915 );
buf ( n5781 , n2028 );
buf ( n5782 , n594 );
buf ( n5783 , n694 );
buf ( n5784 , n1942 );
buf ( n5785 , n671 );
buf ( n5786 , n1560 );
buf ( n5787 , n1348 );
buf ( n5788 , n1103 );
buf ( n5789 , n667 );
buf ( n5790 , n1071 );
buf ( n5791 , n447 );
buf ( n5792 , n1191 );
buf ( n5793 , n1371 );
buf ( n5794 , n279 );
buf ( n5795 , n1707 );
buf ( n5796 , n1844 );
buf ( n5797 , n1544 );
buf ( n5798 , n1345 );
buf ( n5799 , n1066 );
buf ( n5800 , n591 );
buf ( n5801 , n363 );
buf ( n5802 , n335 );
buf ( n5803 , n787 );
buf ( n5804 , n2079 );
buf ( n5805 , n1065 );
buf ( n5806 , n891 );
buf ( n5807 , n1650 );
buf ( n5808 , n45 );
buf ( n5809 , n1823 );
buf ( n5810 , n1881 );
buf ( n5811 , n797 );
buf ( n5812 , n1626 );
buf ( n5813 , n402 );
buf ( n5814 , n1833 );
buf ( n5815 , n2000 );
buf ( n5816 , n955 );
buf ( n5817 , n714 );
buf ( n5818 , n30 );
buf ( n5819 , n1091 );
buf ( n5820 , n954 );
buf ( n5821 , n1599 );
buf ( n5822 , n960 );
buf ( n5823 , n1542 );
buf ( n5824 , n774 );
buf ( n5825 , n795 );
buf ( n5826 , n1518 );
buf ( n5827 , n1527 );
buf ( n5828 , n1087 );
buf ( n5829 , n193 );
buf ( n5830 , n141 );
buf ( n5831 , n1594 );
buf ( n5832 , n1500 );
buf ( n5833 , n1826 );
buf ( n5834 , n1041 );
buf ( n5835 , n1925 );
buf ( n5836 , n2030 );
buf ( n5837 , n1493 );
buf ( n5838 , n1005 );
buf ( n5839 , n225 );
buf ( n5840 , n77 );
buf ( n5841 , n2109 );
buf ( n5842 , n1482 );
buf ( n5843 , n14 );
buf ( n5844 , n434 );
buf ( n5845 , n1662 );
buf ( n5846 , n1311 );
buf ( n5847 , n376 );
buf ( n5848 , n1261 );
buf ( n5849 , n1019 );
buf ( n5850 , n2015 );
buf ( n5851 , n78 );
buf ( n5852 , n637 );
buf ( n5853 , n1964 );
buf ( n5854 , n1174 );
buf ( n5855 , n442 );
buf ( n5856 , n1434 );
buf ( n5857 , n1061 );
buf ( n5858 , n1490 );
buf ( n5859 , n329 );
buf ( n5860 , n810 );
buf ( n5861 , n850 );
buf ( n5862 , n1377 );
buf ( n5863 , n2167 );
buf ( n5864 , n846 );
buf ( n5865 , n315 );
buf ( n5866 , n1687 );
buf ( n5867 , n1864 );
buf ( n5868 , n1122 );
buf ( n5869 , n2108 );
buf ( n5870 , n956 );
buf ( n5871 , n1829 );
buf ( n5872 , n1671 );
buf ( n5873 , n852 );
buf ( n5874 , n1686 );
buf ( n5875 , n544 );
buf ( n5876 , n35 );
buf ( n5877 , n2078 );
buf ( n5878 , n7 );
buf ( n5879 , n357 );
buf ( n5880 , n1215 );
buf ( n5881 , n2169 );
buf ( n5882 , n1025 );
buf ( n5883 , n1856 );
buf ( n5884 , n1607 );
buf ( n5885 , n321 );
buf ( n5886 , n166 );
buf ( n5887 , n939 );
buf ( n5888 , n602 );
buf ( n5889 , n914 );
buf ( n5890 , n2104 );
buf ( n5891 , n1048 );
buf ( n5892 , n849 );
buf ( n5893 , n1360 );
buf ( n5894 , n1356 );
buf ( n5895 , n66 );
buf ( n5896 , n1885 );
buf ( n5897 , n1724 );
buf ( n5898 , n1392 );
buf ( n5899 , n1949 );
buf ( n5900 , n1673 );
buf ( n5901 , n1770 );
buf ( n5902 , n1725 );
buf ( n5903 , n879 );
buf ( n5904 , n1114 );
buf ( n5905 , n1148 );
buf ( n5906 , n270 );
buf ( n5907 , n2154 );
buf ( n5908 , n870 );
buf ( n5909 , n1193 );
buf ( n5910 , n1175 );
buf ( n5911 , n575 );
buf ( n5912 , n125 );
buf ( n5913 , n398 );
buf ( n5914 , n1778 );
buf ( n5915 , n871 );
buf ( n5916 , n1656 );
buf ( n5917 , n449 );
buf ( n5918 , n1382 );
buf ( n5919 , n950 );
buf ( n5920 , n264 );
buf ( n5921 , n1808 );
buf ( n5922 , n1731 );
buf ( n5923 , n347 );
buf ( n5924 , n559 );
buf ( n5925 , n1401 );
buf ( n5926 , n1898 );
buf ( n5927 , n1859 );
buf ( n5928 , n1038 );
buf ( n5929 , n1529 );
buf ( n5930 , n337 );
buf ( n5931 , n565 );
buf ( n5932 , n1910 );
buf ( n5933 , n120 );
buf ( n5934 , n801 );
buf ( n5935 , n1186 );
buf ( n5936 , n1331 );
buf ( n5937 , n1632 );
buf ( n5938 , n318 );
buf ( n5939 , n277 );
buf ( n5940 , n953 );
buf ( n5941 , n147 );
buf ( n5942 , n96 );
buf ( n5943 , n512 );
buf ( n5944 , n580 );
buf ( n5945 , n1242 );
buf ( n5946 , n1342 );
buf ( n5947 , n959 );
buf ( n5948 , n173 );
buf ( n5949 , n1264 );
buf ( n5950 , n1900 );
buf ( n5951 , n2069 );
buf ( n5952 , n983 );
buf ( n5953 , n22 );
buf ( n5954 , n1620 );
buf ( n5955 , n943 );
buf ( n5956 , n910 );
buf ( n5957 , n1292 );
buf ( n5958 , n627 );
buf ( n5959 , n1366 );
buf ( n5960 , n1892 );
buf ( n5961 , n1559 );
buf ( n5962 , n1698 );
buf ( n5963 , n1419 );
buf ( n5964 , n2171 );
buf ( n5965 , n190 );
buf ( n5966 , n122 );
buf ( n5967 , n1236 );
buf ( n5968 , n1468 );
buf ( n5969 , n222 );
buf ( n5970 , n1753 );
buf ( n5971 , n132 );
buf ( n5972 , n1874 );
buf ( n5973 , n647 );
buf ( n5974 , n725 );
buf ( n5975 , n182 );
buf ( n5976 , n877 );
buf ( n5977 , n348 );
buf ( n5978 , n63 );
buf ( n5979 , n289 );
buf ( n5980 , n1055 );
buf ( n5981 , n1540 );
buf ( n5982 , n1744 );
buf ( n5983 , n2113 );
buf ( n5984 , n1837 );
buf ( n5985 , n198 );
buf ( n5986 , n214 );
buf ( n5987 , n1815 );
buf ( n5988 , n1491 );
buf ( n5989 , n818 );
buf ( n5990 , n1204 );
buf ( n5991 , n551 );
buf ( n5992 , n320 );
buf ( n5993 , n2048 );
buf ( n5994 , n825 );
buf ( n5995 , n501 );
buf ( n5996 , n1691 );
buf ( n5997 , n1275 );
buf ( n5998 , n1008 );
buf ( n5999 , n968 );
buf ( n6000 , n1959 );
buf ( n6001 , n178 );
buf ( n6002 , n1986 );
buf ( n6003 , n382 );
buf ( n6004 , n129 );
buf ( n6005 , n1977 );
buf ( n6006 , n1504 );
buf ( n6007 , n649 );
buf ( n6008 , n800 );
buf ( n6009 , n639 );
buf ( n6010 , n1127 );
buf ( n6011 , n303 );
buf ( n6012 , n1424 );
buf ( n6013 , n1155 );
buf ( n6014 , n425 );
buf ( n6015 , n346 );
buf ( n6016 , n1505 );
buf ( n6017 , n642 );
buf ( n6018 , n82 );
buf ( n6019 , n2103 );
buf ( n6020 , n572 );
buf ( n6021 , n743 );
buf ( n6022 , n2026 );
buf ( n6023 , n771 );
buf ( n6024 , n2153 );
buf ( n6025 , n1082 );
buf ( n6026 , n41 );
buf ( n6027 , n1126 );
buf ( n6028 , n298 );
buf ( n6029 , n1151 );
buf ( n6030 , n79 );
buf ( n6031 , n1975 );
buf ( n6032 , n605 );
buf ( n6033 , n1159 );
buf ( n6034 , n248 );
buf ( n6035 , n1570 );
buf ( n6036 , n1969 );
buf ( n6037 , n906 );
buf ( n6038 , n2062 );
buf ( n6039 , n549 );
buf ( n6040 , n1365 );
buf ( n6041 , n441 );
buf ( n6042 , n306 );
buf ( n6043 , n158 );
buf ( n6044 , n1304 );
buf ( n6045 , n617 );
buf ( n6046 , n1116 );
buf ( n6047 , n2025 );
buf ( n6048 , n740 );
buf ( n6049 , n1062 );
buf ( n6050 , n699 );
buf ( n6051 , n1222 );
buf ( n6052 , n706 );
buf ( n6053 , n1136 );
buf ( n6054 , n1492 );
buf ( n6055 , n1860 );
buf ( n6056 , n495 );
buf ( n6057 , n53 );
buf ( n6058 , n262 );
buf ( n6059 , n1718 );
buf ( n6060 , n1109 );
buf ( n6061 , n157 );
buf ( n6062 , n1543 );
buf ( n6063 , n632 );
buf ( n6064 , n1573 );
buf ( n6065 , n188 );
buf ( n6066 , n2004 );
buf ( n6067 , n713 );
buf ( n6068 , n1567 );
buf ( n6069 , n1029 );
buf ( n6070 , n1169 );
buf ( n6071 , n1595 );
buf ( n6072 , n1524 );
buf ( n6073 , n201 );
buf ( n6074 , n2074 );
buf ( n6075 , n866 );
buf ( n6076 , n1102 );
buf ( n6077 , n107 );
buf ( n6078 , n2 );
buf ( n6079 , n931 );
buf ( n6080 , n598 );
buf ( n6081 , n663 );
buf ( n6082 , n2037 );
buf ( n6083 , n179 );
buf ( n6084 , n2160 );
buf ( n6085 , n1775 );
buf ( n6086 , n2180 );
buf ( n6087 , n2052 );
buf ( n6088 , n777 );
buf ( n6089 , n845 );
buf ( n6090 , n1520 );
buf ( n6091 , n2063 );
buf ( n6092 , n1947 );
buf ( n6093 , n1145 );
buf ( n6094 , n1683 );
buf ( n6095 , n1375 );
buf ( n6096 , n1129 );
buf ( n6097 , n209 );
buf ( n6098 , n47 );
buf ( n6099 , n1760 );
buf ( n6100 , n1115 );
buf ( n6101 , n1682 );
buf ( n6102 , n1247 );
buf ( n6103 , n1067 );
buf ( n6104 , n146 );
buf ( n6105 , n1997 );
buf ( n6106 , n973 );
buf ( n6107 , n1830 );
buf ( n6108 , n520 );
buf ( n6109 , n1101 );
buf ( n6110 , n1807 );
buf ( n6111 , n793 );
buf ( n6112 , n662 );
buf ( n6113 , n290 );
buf ( n6114 , n127 );
buf ( n6115 , n1359 );
buf ( n6116 , n1095 );
buf ( n6117 , n776 );
buf ( n6118 , n1161 );
buf ( n6119 , n1689 );
buf ( n6120 , n940 );
buf ( n6121 , n116 );
buf ( n6122 , n2098 );
buf ( n6123 , n1083 );
buf ( n6124 , n109 );
buf ( n6125 , n1854 );
buf ( n6126 , n938 );
buf ( n6127 , n863 );
buf ( n6128 , n1813 );
buf ( n6129 , n38 );
buf ( n6130 , n1962 );
buf ( n6131 , n695 );
buf ( n6132 , n646 );
buf ( n6133 , n1060 );
buf ( n6134 , n1616 );
buf ( n6135 , n1111 );
buf ( n6136 , n634 );
buf ( n6137 , n1894 );
buf ( n6138 , n1899 );
buf ( n6139 , n1233 );
buf ( n6140 , n1097 );
buf ( n6141 , n987 );
buf ( n6142 , n1252 );
buf ( n6143 , n1396 );
buf ( n6144 , n856 );
buf ( n6145 , n2129 );
buf ( n6146 , n220 );
buf ( n6147 , n1921 );
buf ( n6148 , n1069 );
buf ( n6149 , n1042 );
buf ( n6150 , n2035 );
buf ( n6151 , n204 );
buf ( n6152 , n2019 );
buf ( n6153 , n61 );
buf ( n6154 , n1270 );
buf ( n6155 , n2095 );
buf ( n6156 , n775 );
buf ( n6157 , n1449 );
buf ( n6158 , n485 );
buf ( n6159 , n1795 );
buf ( n6160 , n1547 );
buf ( n6161 , n1639 );
buf ( n6162 , n490 );
buf ( n6163 , n2128 );
buf ( n6164 , n2080 );
buf ( n6165 , n1361 );
buf ( n6166 , n1602 );
buf ( n6167 , n689 );
buf ( n6168 , n2059 );
buf ( n6169 , n474 );
buf ( n6170 , n1352 );
buf ( n6171 , n528 );
buf ( n6172 , n1228 );
buf ( n6173 , n1985 );
buf ( n6174 , n1026 );
buf ( n6175 , n2158 );
buf ( n6176 , n1648 );
buf ( n6177 , n1276 );
buf ( n6178 , n128 );
buf ( n6179 , n1617 );
buf ( n6180 , n539 );
buf ( n6181 , n1905 );
buf ( n6182 , n1800 );
buf ( n6183 , n1014 );
buf ( n6184 , n2183 );
buf ( n6185 , n734 );
buf ( n6186 , n1931 );
buf ( n6187 , n1970 );
buf ( n6188 , n1759 );
buf ( n6189 , n1280 );
buf ( n6190 , n759 );
buf ( n6191 , n1941 );
buf ( n6192 , n608 );
buf ( n6193 , n358 );
buf ( n6194 , n497 );
buf ( n6195 , n1339 );
buf ( n6196 , n2068 );
buf ( n6197 , n2057 );
buf ( n6198 , n1842 );
buf ( n6199 , n170 );
buf ( n6200 , n1980 );
buf ( n6201 , n292 );
buf ( n6202 , n185 );
buf ( n6203 , n502 );
buf ( n6204 , n707 );
buf ( n6205 , n126 );
buf ( n6206 , n2131 );
buf ( n6207 , n1920 );
buf ( n6208 , n1593 );
buf ( n6209 , n389 );
buf ( n6210 , n1798 );
buf ( n6211 , n518 );
buf ( n6212 , n508 );
buf ( n6213 , n331 );
buf ( n6214 , n1961 );
buf ( n6215 , n822 );
buf ( n6216 , n611 );
buf ( n6217 , n704 );
buf ( n6218 , n1940 );
buf ( n6219 , n1195 );
buf ( n6220 , n1934 );
buf ( n6221 , n1059 );
buf ( n6222 , n253 );
buf ( n6223 , n1545 );
buf ( n6224 , n2043 );
buf ( n6225 , n1615 );
buf ( n6226 , n1714 );
buf ( n6227 , n1502 );
buf ( n6228 , n1094 );
buf ( n6229 , n234 );
buf ( n6230 , n74 );
buf ( n6231 , n111 );
buf ( n6232 , n1260 );
buf ( n6233 , n183 );
buf ( n6234 , n796 );
buf ( n6235 , n362 );
buf ( n6236 , n784 );
buf ( n6237 , n1131 );
buf ( n6238 , n375 );
buf ( n6239 , n355 );
buf ( n6240 , n828 );
buf ( n6241 , n2081 );
buf ( n6242 , n865 );
buf ( n6243 , n124 );
buf ( n6244 , n670 );
buf ( n6245 , n1445 );
buf ( n6246 , n932 );
buf ( n6247 , n1625 );
buf ( n6248 , n1793 );
buf ( n6249 , n1847 );
buf ( n6250 , n199 );
buf ( n6251 , n364 );
buf ( n6252 , n330 );
buf ( n6253 , n1383 );
buf ( n6254 , n815 );
buf ( n6255 , n509 );
buf ( n6256 , n155 );
buf ( n6257 , n1028 );
buf ( n6258 , n1487 );
buf ( n6259 , n1068 );
buf ( n6260 , n1565 );
buf ( n6261 , n568 );
buf ( n6262 , n468 );
buf ( n6263 , n2072 );
buf ( n6264 , n1531 );
buf ( n6265 , n1254 );
buf ( n6266 , n1387 );
buf ( n6267 , n208 );
buf ( n6268 , n1791 );
buf ( n6269 , n958 );
buf ( n6270 , n990 );
buf ( n6271 , n1845 );
buf ( n6272 , n1653 );
buf ( n6273 , n1517 );
buf ( n6274 , n196 );
buf ( n6275 , n1995 );
buf ( n6276 , n1470 );
buf ( n6277 , n168 );
buf ( n6278 , n105 );
buf ( n6279 , n1381 );
buf ( n6280 , n2123 );
buf ( n6281 , n1799 );
buf ( n6282 , n806 );
buf ( n6283 , n904 );
buf ( n6284 , n119 );
buf ( n6285 , n1875 );
buf ( n6286 , n1297 );
buf ( n6287 , n1663 );
buf ( n6288 , n1469 );
buf ( n6289 , n1624 );
buf ( n6290 , n1015 );
buf ( n6291 , n2125 );
buf ( n6292 , n1211 );
buf ( n6293 , n1027 );
buf ( n6294 , n786 );
buf ( n6295 , n1635 );
buf ( n6296 , n963 );
buf ( n6297 , n1507 );
buf ( n6298 , n52 );
buf ( n6299 , n84 );
buf ( n6300 , n915 );
buf ( n6301 , n1386 );
buf ( n6302 , n1882 );
buf ( n6303 , n164 );
buf ( n6304 , n305 );
buf ( n6305 , n1165 );
buf ( n6306 , n316 );
buf ( n6307 , n1822 );
buf ( n6308 , n998 );
buf ( n6309 , n2064 );
buf ( n6310 , n812 );
buf ( n6311 , n638 );
buf ( n6312 , n1271 );
buf ( n6313 , n1225 );
buf ( n6314 , n807 );
buf ( n6315 , n1415 );
buf ( n6316 , n1406 );
buf ( n6317 , n1020 );
buf ( n6318 , n241 );
buf ( n6319 , n864 );
buf ( n6320 , n683 );
buf ( n6321 , n1411 );
buf ( n6322 , n1440 );
buf ( n6323 , n435 );
buf ( n6324 , n86 );
buf ( n6325 , n1398 );
buf ( n6326 , n403 );
buf ( n6327 , n1600 );
buf ( n6328 , n620 );
buf ( n6329 , n378 );
buf ( n6330 , n1979 );
buf ( n6331 , n1851 );
buf ( n6332 , n1056 );
buf ( n6333 , n2021 );
buf ( n6334 , n1722 );
buf ( n6335 , n2082 );
buf ( n6336 , n967 );
buf ( n6337 , n1971 );
buf ( n6338 , n861 );
buf ( n6339 , n460 );
buf ( n6340 , n70 );
buf ( n6341 , n834 );
buf ( n6342 , n1422 );
buf ( n6343 , n2136 );
buf ( n6344 , n1227 );
buf ( n6345 , n2009 );
buf ( n6346 , n577 );
buf ( n6347 , n2140 );
buf ( n6348 , n1871 );
buf ( n6349 , n1319 );
buf ( n6350 , n537 );
buf ( n6351 , n1641 );
buf ( n6352 , n561 );
buf ( n6353 , n1389 );
buf ( n6354 , n1665 );
buf ( n6355 , n517 );
buf ( n6356 , n1956 );
buf ( n6357 , n1442 );
buf ( n6358 , n1752 );
buf ( n6359 , n1475 );
buf ( n6360 , n391 );
buf ( n6361 , n1032 );
buf ( n6362 , n1532 );
buf ( n6363 , n1538 );
buf ( n6364 , n1677 );
buf ( n6365 , n272 );
buf ( n6366 , n1896 );
buf ( n6367 , n267 );
buf ( n6368 , n404 );
buf ( n6369 , n1368 );
buf ( n6370 , n1933 );
buf ( n6371 , n1785 );
buf ( n6372 , n411 );
buf ( n6373 , n1563 );
buf ( n6374 , n1935 );
buf ( n6375 , n172 );
buf ( n6376 , n1033 );
buf ( n6377 , n1216 );
buf ( n6378 , n1537 );
buf ( n6379 , n1144 );
buf ( n6380 , n522 );
buf ( n6381 , n1840 );
buf ( n6382 , n532 );
buf ( n6383 , n1223 );
buf ( n6384 , n878 );
buf ( n6385 , n724 );
buf ( n6386 , n2114 );
buf ( n6387 , n354 );
buf ( n6388 , n309 );
buf ( n6389 , n100 );
buf ( n6390 , n89 );
buf ( n6391 , n731 );
buf ( n6392 , n467 );
buf ( n6393 , n229 );
buf ( n6394 , n827 );
buf ( n6395 , n913 );
buf ( n6396 , n1717 );
buf ( n6397 , n1402 );
buf ( n6398 , n935 );
buf ( n6399 , n2157 );
buf ( n6400 , n1551 );
buf ( n6401 , n2093 );
buf ( n6402 , n1646 );
buf ( n6403 , n324 );
buf ( n6404 , n2051 );
buf ( n6405 , n1556 );
buf ( n6406 , n381 );
buf ( n6407 , n1957 );
buf ( n6408 , n221 );
buf ( n6409 , n1323 );
buf ( n6410 , n556 );
buf ( n6411 , n419 );
buf ( n6412 , n1105 );
buf ( n6413 , n2056 );
buf ( n6414 , n421 );
buf ( n6415 , n858 );
buf ( n6416 , n73 );
buf ( n6417 , n1660 );
buf ( n6418 , n49 );
buf ( n6419 , n1654 );
buf ( n6420 , n2086 );
buf ( n6421 , n1810 );
buf ( n6422 , n1400 );
buf ( n6423 , n1171 );
buf ( n6424 , n698 );
buf ( n6425 , n1569 );
buf ( n6426 , n1849 );
buf ( n6427 , n312 );
buf ( n6428 , n478 );
buf ( n6429 , n16 );
buf ( n6430 , n284 );
buf ( n6431 , n2090 );
buf ( n6432 , n233 );
buf ( n6433 , n1818 );
buf ( n6434 , n1125 );
buf ( n6435 , n103 );
buf ( n6436 , n951 );
buf ( n6437 , n1640 );
buf ( n6438 , n1732 );
buf ( n6439 , n799 );
buf ( n6440 , n1218 );
buf ( n6441 , n1530 );
buf ( n6442 , n56 );
buf ( n6443 , n590 );
buf ( n6444 , n2017 );
buf ( n6445 , n1269 );
buf ( n6446 , n1454 );
buf ( n6447 , n426 );
buf ( n6448 , n12 );
buf ( n6449 , n1695 );
buf ( n6450 , n546 );
buf ( n6451 , n1009 );
buf ( n6452 , n593 );
buf ( n6453 , n34 );
buf ( n6454 , n564 );
buf ( n6455 , n1139 );
buf ( n6456 , n1497 );
buf ( n6457 , n90 );
buf ( n6458 , n1907 );
buf ( n6459 , n688 );
buf ( n6460 , n377 );
buf ( n6461 , n1608 );
buf ( n6462 , n91 );
buf ( n6463 , n1239 );
buf ( n6464 , n1739 );
buf ( n6465 , n1692 );
buf ( n6466 , n237 );
buf ( n6467 , n1734 );
buf ( n6468 , n1054 );
buf ( n6469 , n325 );
buf ( n6470 , n1919 );
buf ( n6471 , n1924 );
buf ( n6472 , n524 );
buf ( n6473 , n36 );
buf ( n6474 , n2178 );
buf ( n6475 , n1668 );
buf ( n6476 , n2089 );
buf ( n6477 , n881 );
buf ( n6478 , n1834 );
buf ( n6479 , n1604 );
buf ( n6480 , n832 );
buf ( n6481 , n902 );
buf ( n6482 , n1796 );
buf ( n6483 , n2041 );
buf ( n6484 , n487 );
buf ( n6485 , n1501 );
buf ( n6486 , n57 );
buf ( n6487 , n1916 );
buf ( n6488 , n975 );
buf ( n6489 , n2165 );
buf ( n6490 , n97 );
buf ( n6491 , n547 );
buf ( n6492 , n566 );
buf ( n6493 , n543 );
buf ( n6494 , n1788 );
buf ( n6495 , n230 );
buf ( n6496 , n1857 );
buf ( n6497 , n152 );
buf ( n6498 , n252 );
buf ( n6499 , n778 );
buf ( n6500 , n380 );
buf ( n6501 , n770 );
buf ( n6502 , n1690 );
buf ( n6503 , n1913 );
buf ( n6504 , n763 );
buf ( n6505 , n1017 );
buf ( n6506 , n1580 );
buf ( n6507 , n969 );
buf ( n6508 , n1742 );
buf ( n6509 , n336 );
buf ( n6510 , n945 );
buf ( n6511 , n486 );
buf ( n6512 , n571 );
buf ( n6513 , n1064 );
buf ( n6514 , n1679 );
buf ( n6515 , n217 );
buf ( n6516 , n1509 );
buf ( n6517 , n1189 );
buf ( n6518 , n1436 );
buf ( n6519 , n1819 );
buf ( n6520 , n72 );
buf ( n6521 , n231 );
buf ( n6522 , n1733 );
buf ( n6523 , n1809 );
buf ( n6524 , n1209 );
buf ( n6525 , n1427 );
buf ( n6526 , n1780 );
buf ( n6527 , n2173 );
buf ( n6528 , n984 );
buf ( n6529 , n383 );
buf ( n6530 , n661 );
buf ( n6531 , n32 );
buf ( n6532 , n452 );
buf ( n6533 , n24 );
buf ( n6534 , n1883 );
buf ( n6535 , n2060 );
buf ( n6536 , n1443 );
buf ( n6537 , n110 );
buf ( n6538 , n1836 );
buf ( n6539 , n1206 );
buf ( n6540 , n1409 );
buf ( n6541 , n2007 );
buf ( n6542 , n2084 );
buf ( n6543 , n1074 );
buf ( n6544 , n2102 );
buf ( n6545 , n457 );
buf ( n6546 , n410 );
buf ( n6547 , n433 );
buf ( n6548 , n9 );
buf ( n6549 , n261 );
buf ( n6550 , n729 );
buf ( n6551 , n333 );
buf ( n6552 , n804 );
buf ( n6553 , n2126 );
buf ( n6554 , n268 );
buf ( n6555 , n1318 );
buf ( n6556 , n737 );
buf ( n6557 , n909 );
buf ( n6558 , n1761 );
buf ( n6559 , n2027 );
buf ( n6560 , n1783 );
buf ( n6561 , n1210 );
buf ( n6562 , n1273 );
buf ( n6563 , n1281 );
buf ( n6564 , n1955 );
buf ( n6565 , n1178 );
buf ( n6566 , n579 );
buf ( n6567 , n1652 );
buf ( n6568 , n2018 );
buf ( n6569 , n44 );
buf ( n6570 , n1581 );
buf ( n6571 , n2011 );
buf ( n6572 , n1649 );
buf ( n6573 , n993 );
buf ( n6574 , n216 );
buf ( n6575 , n1194 );
buf ( n6576 , n1200 );
buf ( n6577 , n4394 );
buf ( n6578 , n6577 );
not ( n6579 , n6578 );
buf ( n6580 , n4395 );
buf ( n6581 , n4396 );
not ( n6582 , n6580 );
and ( n6583 , n6581 , n6582 );
or ( n6584 , n6580 , n6583 );
not ( n6585 , n6584 );
buf ( n6586 , n4397 );
and ( n6587 , n6585 , n6586 );
not ( n6588 , n6583 );
buf ( n6589 , n4398 );
and ( n6590 , n6588 , n6589 );
buf ( n6591 , n4399 );
xor ( n6592 , n6591 , n6589 );
and ( n6593 , n6592 , n6583 );
or ( n6594 , n6590 , n6593 );
not ( n6595 , n6583 );
buf ( n6596 , n4400 );
and ( n6597 , n6595 , n6596 );
buf ( n6598 , n4401 );
xor ( n6599 , n6598 , n6596 );
and ( n6600 , n6599 , n6583 );
or ( n6601 , n6597 , n6600 );
not ( n6602 , n6583 );
buf ( n6603 , n4402 );
and ( n6604 , n6602 , n6603 );
buf ( n6605 , n4403 );
xor ( n6606 , n6605 , n6603 );
and ( n6607 , n6606 , n6583 );
or ( n6608 , n6604 , n6607 );
xor ( n6609 , n6601 , n6608 );
buf ( n6610 , n4404 );
xor ( n6611 , n6609 , n6610 );
buf ( n6612 , n4405 );
xor ( n6613 , n6611 , n6612 );
buf ( n6614 , n4406 );
xor ( n6615 , n6613 , n6614 );
xor ( n6616 , n6594 , n6615 );
not ( n6617 , n6583 );
buf ( n6618 , n4407 );
and ( n6619 , n6617 , n6618 );
buf ( n6620 , n4408 );
xor ( n6621 , n6620 , n6618 );
and ( n6622 , n6621 , n6583 );
or ( n6623 , n6619 , n6622 );
not ( n6624 , n6583 );
buf ( n6625 , n4409 );
and ( n6626 , n6624 , n6625 );
buf ( n6627 , n4410 );
xor ( n6628 , n6627 , n6625 );
and ( n6629 , n6628 , n6583 );
or ( n6630 , n6626 , n6629 );
xor ( n6631 , n6623 , n6630 );
buf ( n6632 , n4411 );
xor ( n6633 , n6631 , n6632 );
buf ( n6634 , n4412 );
xor ( n6635 , n6633 , n6634 );
not ( n6636 , n6635 );
xor ( n6637 , n6616 , n6636 );
not ( n6638 , n6583 );
buf ( n6639 , n4413 );
and ( n6640 , n6638 , n6639 );
buf ( n6641 , n4414 );
xor ( n6642 , n6641 , n6639 );
and ( n6643 , n6642 , n6583 );
or ( n6644 , n6640 , n6643 );
not ( n6645 , n6583 );
buf ( n6646 , n4415 );
and ( n6647 , n6645 , n6646 );
buf ( n6648 , n4416 );
xor ( n6649 , n6648 , n6646 );
and ( n6650 , n6649 , n6583 );
or ( n6651 , n6647 , n6650 );
buf ( n6652 , n4417 );
xor ( n6653 , n6651 , n6652 );
buf ( n6654 , n4418 );
xor ( n6655 , n6653 , n6654 );
buf ( n6656 , n4419 );
xor ( n6657 , n6655 , n6656 );
buf ( n6658 , n4420 );
xor ( n6659 , n6657 , n6658 );
xor ( n6660 , n6644 , n6659 );
not ( n6661 , n6583 );
buf ( n6662 , n4421 );
and ( n6663 , n6661 , n6662 );
buf ( n6664 , n4422 );
xor ( n6665 , n6664 , n6662 );
and ( n6666 , n6665 , n6583 );
or ( n6667 , n6663 , n6666 );
not ( n6668 , n6583 );
buf ( n6669 , n4423 );
and ( n6670 , n6668 , n6669 );
buf ( n6671 , n4424 );
xor ( n6672 , n6671 , n6669 );
and ( n6673 , n6672 , n6583 );
or ( n6674 , n6670 , n6673 );
xor ( n6675 , n6667 , n6674 );
buf ( n6676 , n4425 );
xor ( n6677 , n6675 , n6676 );
buf ( n6678 , n4426 );
xor ( n6679 , n6677 , n6678 );
buf ( n6680 , n4427 );
xor ( n6681 , n6679 , n6680 );
xor ( n6682 , n6660 , n6681 );
not ( n6683 , n6682 );
buf ( n6684 , n4428 );
not ( n6685 , n6583 );
buf ( n6686 , n4429 );
and ( n6687 , n6685 , n6686 );
buf ( n6688 , n4430 );
xor ( n6689 , n6688 , n6686 );
and ( n6690 , n6689 , n6583 );
or ( n6691 , n6687 , n6690 );
not ( n6692 , n6583 );
buf ( n6693 , n4431 );
and ( n6694 , n6692 , n6693 );
buf ( n6695 , n4432 );
xor ( n6696 , n6695 , n6693 );
and ( n6697 , n6696 , n6583 );
or ( n6698 , n6694 , n6697 );
xor ( n6699 , n6691 , n6698 );
buf ( n6700 , n4433 );
xor ( n6701 , n6699 , n6700 );
buf ( n6702 , n4434 );
xor ( n6703 , n6701 , n6702 );
buf ( n6704 , n4435 );
xor ( n6705 , n6703 , n6704 );
xor ( n6706 , n6684 , n6705 );
not ( n6707 , n6583 );
buf ( n6708 , n4436 );
and ( n6709 , n6707 , n6708 );
buf ( n6710 , n4437 );
xor ( n6711 , n6710 , n6708 );
and ( n6712 , n6711 , n6583 );
or ( n6713 , n6709 , n6712 );
not ( n6714 , n6583 );
buf ( n6715 , n4438 );
and ( n6716 , n6714 , n6715 );
buf ( n6717 , n4439 );
xor ( n6718 , n6717 , n6715 );
and ( n6719 , n6718 , n6583 );
or ( n6720 , n6716 , n6719 );
xor ( n6721 , n6713 , n6720 );
buf ( n6722 , n4440 );
xor ( n6723 , n6721 , n6722 );
buf ( n6724 , n4441 );
xor ( n6725 , n6723 , n6724 );
buf ( n6726 , n4442 );
xor ( n6727 , n6725 , n6726 );
xor ( n6728 , n6706 , n6727 );
and ( n6729 , n6683 , n6728 );
xor ( n6730 , n6637 , n6729 );
buf ( n6731 , n4443 );
not ( n6732 , n6583 );
buf ( n6733 , n4444 );
and ( n6734 , n6732 , n6733 );
buf ( n6735 , n4445 );
xor ( n6736 , n6735 , n6733 );
and ( n6737 , n6736 , n6583 );
or ( n6738 , n6734 , n6737 );
not ( n6739 , n6583 );
buf ( n6740 , n4446 );
and ( n6741 , n6739 , n6740 );
buf ( n6742 , n4447 );
xor ( n6743 , n6742 , n6740 );
and ( n6744 , n6743 , n6583 );
or ( n6745 , n6741 , n6744 );
xor ( n6746 , n6738 , n6745 );
buf ( n6747 , n4448 );
xor ( n6748 , n6746 , n6747 );
buf ( n6749 , n4449 );
xor ( n6750 , n6748 , n6749 );
buf ( n6751 , n4450 );
xor ( n6752 , n6750 , n6751 );
xor ( n6753 , n6731 , n6752 );
not ( n6754 , n6583 );
buf ( n6755 , n4451 );
and ( n6756 , n6754 , n6755 );
buf ( n6757 , n4452 );
xor ( n6758 , n6757 , n6755 );
and ( n6759 , n6758 , n6583 );
or ( n6760 , n6756 , n6759 );
not ( n6761 , n6583 );
buf ( n6762 , n4453 );
and ( n6763 , n6761 , n6762 );
buf ( n6764 , n4454 );
xor ( n6765 , n6764 , n6762 );
and ( n6766 , n6765 , n6583 );
or ( n6767 , n6763 , n6766 );
xor ( n6768 , n6760 , n6767 );
buf ( n6769 , n4455 );
xor ( n6770 , n6768 , n6769 );
buf ( n6771 , n4456 );
xor ( n6772 , n6770 , n6771 );
buf ( n6773 , n4457 );
xor ( n6774 , n6772 , n6773 );
xor ( n6775 , n6753 , n6774 );
not ( n6776 , n6583 );
buf ( n6777 , n4458 );
and ( n6778 , n6776 , n6777 );
buf ( n6779 , n4459 );
xor ( n6780 , n6779 , n6777 );
and ( n6781 , n6780 , n6583 );
or ( n6782 , n6778 , n6781 );
not ( n6783 , n6583 );
buf ( n6784 , n4460 );
and ( n6785 , n6783 , n6784 );
buf ( n6786 , n4461 );
xor ( n6787 , n6786 , n6784 );
and ( n6788 , n6787 , n6583 );
or ( n6789 , n6785 , n6788 );
buf ( n6790 , n4462 );
xor ( n6791 , n6789 , n6790 );
buf ( n6792 , n4463 );
xor ( n6793 , n6791 , n6792 );
buf ( n6794 , n4464 );
xor ( n6795 , n6793 , n6794 );
buf ( n6796 , n4465 );
xor ( n6797 , n6795 , n6796 );
xor ( n6798 , n6782 , n6797 );
not ( n6799 , n6583 );
buf ( n6800 , n4466 );
and ( n6801 , n6799 , n6800 );
buf ( n6802 , n4467 );
xor ( n6803 , n6802 , n6800 );
and ( n6804 , n6803 , n6583 );
or ( n6805 , n6801 , n6804 );
not ( n6806 , n6583 );
buf ( n6807 , n4468 );
and ( n6808 , n6806 , n6807 );
buf ( n6809 , n4469 );
xor ( n6810 , n6809 , n6807 );
and ( n6811 , n6810 , n6583 );
or ( n6812 , n6808 , n6811 );
xor ( n6813 , n6805 , n6812 );
buf ( n6814 , n4470 );
xor ( n6815 , n6813 , n6814 );
buf ( n6816 , n4471 );
xor ( n6817 , n6815 , n6816 );
buf ( n6818 , n4472 );
xor ( n6819 , n6817 , n6818 );
xor ( n6820 , n6798 , n6819 );
not ( n6821 , n6820 );
not ( n6822 , n6583 );
buf ( n6823 , n4473 );
and ( n6824 , n6822 , n6823 );
buf ( n6825 , n4474 );
xor ( n6826 , n6825 , n6823 );
and ( n6827 , n6826 , n6583 );
or ( n6828 , n6824 , n6827 );
not ( n6829 , n6583 );
buf ( n6830 , n4475 );
and ( n6831 , n6829 , n6830 );
buf ( n6832 , n4476 );
xor ( n6833 , n6832 , n6830 );
and ( n6834 , n6833 , n6583 );
or ( n6835 , n6831 , n6834 );
not ( n6836 , n6583 );
buf ( n6837 , n4477 );
and ( n6838 , n6836 , n6837 );
buf ( n6839 , n4478 );
xor ( n6840 , n6839 , n6837 );
and ( n6841 , n6840 , n6583 );
or ( n6842 , n6838 , n6841 );
xor ( n6843 , n6835 , n6842 );
buf ( n6844 , n4479 );
xor ( n6845 , n6843 , n6844 );
buf ( n6846 , n4480 );
xor ( n6847 , n6845 , n6846 );
buf ( n6848 , n4481 );
xor ( n6849 , n6847 , n6848 );
xor ( n6850 , n6828 , n6849 );
not ( n6851 , n6583 );
buf ( n6852 , n4482 );
and ( n6853 , n6851 , n6852 );
buf ( n6854 , n4483 );
xor ( n6855 , n6854 , n6852 );
and ( n6856 , n6855 , n6583 );
or ( n6857 , n6853 , n6856 );
not ( n6858 , n6583 );
buf ( n6859 , n4484 );
and ( n6860 , n6858 , n6859 );
buf ( n6861 , n4485 );
xor ( n6862 , n6861 , n6859 );
and ( n6863 , n6862 , n6583 );
or ( n6864 , n6860 , n6863 );
xor ( n6865 , n6857 , n6864 );
buf ( n6866 , n4486 );
xor ( n6867 , n6865 , n6866 );
buf ( n6868 , n4487 );
xor ( n6869 , n6867 , n6868 );
buf ( n6870 , n4488 );
xor ( n6871 , n6869 , n6870 );
xor ( n6872 , n6850 , n6871 );
and ( n6873 , n6821 , n6872 );
xor ( n6874 , n6775 , n6873 );
buf ( n6875 , n4489 );
not ( n6876 , n6583 );
buf ( n6877 , n4490 );
and ( n6878 , n6876 , n6877 );
buf ( n6879 , n4491 );
xor ( n6880 , n6879 , n6877 );
and ( n6881 , n6880 , n6583 );
or ( n6882 , n6878 , n6881 );
not ( n6883 , n6583 );
buf ( n6884 , n4492 );
and ( n6885 , n6883 , n6884 );
buf ( n6886 , n4493 );
xor ( n6887 , n6886 , n6884 );
and ( n6888 , n6887 , n6583 );
or ( n6889 , n6885 , n6888 );
xor ( n6890 , n6882 , n6889 );
buf ( n6891 , n4494 );
xor ( n6892 , n6890 , n6891 );
buf ( n6893 , n4495 );
xor ( n6894 , n6892 , n6893 );
buf ( n6895 , n4496 );
xor ( n6896 , n6894 , n6895 );
xor ( n6897 , n6875 , n6896 );
not ( n6898 , n6583 );
buf ( n6899 , n4497 );
and ( n6900 , n6898 , n6899 );
buf ( n6901 , n4498 );
xor ( n6902 , n6901 , n6899 );
and ( n6903 , n6902 , n6583 );
or ( n6904 , n6900 , n6903 );
not ( n6905 , n6583 );
buf ( n6906 , n4499 );
and ( n6907 , n6905 , n6906 );
buf ( n6908 , n4500 );
xor ( n6909 , n6908 , n6906 );
and ( n6910 , n6909 , n6583 );
or ( n6911 , n6907 , n6910 );
xor ( n6912 , n6904 , n6911 );
buf ( n6913 , n4501 );
xor ( n6914 , n6912 , n6913 );
buf ( n6915 , n4502 );
xor ( n6916 , n6914 , n6915 );
buf ( n6917 , n4503 );
xor ( n6918 , n6916 , n6917 );
xor ( n6919 , n6897 , n6918 );
not ( n6920 , n6583 );
buf ( n6921 , n4504 );
and ( n6922 , n6920 , n6921 );
buf ( n6923 , n4505 );
xor ( n6924 , n6923 , n6921 );
and ( n6925 , n6924 , n6583 );
or ( n6926 , n6922 , n6925 );
not ( n6927 , n6583 );
buf ( n6928 , n4506 );
and ( n6929 , n6927 , n6928 );
buf ( n6930 , n4507 );
xor ( n6931 , n6930 , n6928 );
and ( n6932 , n6931 , n6583 );
or ( n6933 , n6929 , n6932 );
not ( n6934 , n6583 );
buf ( n6935 , n4508 );
and ( n6936 , n6934 , n6935 );
buf ( n6937 , n4509 );
xor ( n6938 , n6937 , n6935 );
and ( n6939 , n6938 , n6583 );
or ( n6940 , n6936 , n6939 );
xor ( n6941 , n6933 , n6940 );
buf ( n6942 , n4510 );
xor ( n6943 , n6941 , n6942 );
buf ( n6944 , n4511 );
xor ( n6945 , n6943 , n6944 );
buf ( n6946 , n4512 );
xor ( n6947 , n6945 , n6946 );
xor ( n6948 , n6926 , n6947 );
not ( n6949 , n6583 );
buf ( n6950 , n4513 );
and ( n6951 , n6949 , n6950 );
buf ( n6952 , n4514 );
xor ( n6953 , n6952 , n6950 );
and ( n6954 , n6953 , n6583 );
or ( n6955 , n6951 , n6954 );
buf ( n6956 , n4515 );
xor ( n6957 , n6955 , n6956 );
buf ( n6958 , n4516 );
xor ( n6959 , n6957 , n6958 );
buf ( n6960 , n4517 );
xor ( n6961 , n6959 , n6960 );
buf ( n6962 , n4518 );
xor ( n6963 , n6961 , n6962 );
xor ( n6964 , n6948 , n6963 );
not ( n6965 , n6964 );
buf ( n6966 , n4519 );
not ( n6967 , n6583 );
buf ( n6968 , n4520 );
and ( n6969 , n6967 , n6968 );
buf ( n6970 , n4521 );
xor ( n6971 , n6970 , n6968 );
and ( n6972 , n6971 , n6583 );
or ( n6973 , n6969 , n6972 );
not ( n6974 , n6583 );
buf ( n6975 , n4522 );
and ( n6976 , n6974 , n6975 );
buf ( n6977 , n4523 );
xor ( n6978 , n6977 , n6975 );
and ( n6979 , n6978 , n6583 );
or ( n6980 , n6976 , n6979 );
xor ( n6981 , n6973 , n6980 );
buf ( n6982 , n4524 );
xor ( n6983 , n6981 , n6982 );
buf ( n6984 , n4525 );
xor ( n6985 , n6983 , n6984 );
buf ( n6986 , n4526 );
xor ( n6987 , n6985 , n6986 );
xor ( n6988 , n6966 , n6987 );
not ( n6989 , n6583 );
buf ( n6990 , n4527 );
and ( n6991 , n6989 , n6990 );
buf ( n6992 , n4528 );
xor ( n6993 , n6992 , n6990 );
and ( n6994 , n6993 , n6583 );
or ( n6995 , n6991 , n6994 );
not ( n6996 , n6583 );
buf ( n6997 , n4529 );
and ( n6998 , n6996 , n6997 );
buf ( n6999 , n4530 );
xor ( n7000 , n6999 , n6997 );
and ( n7001 , n7000 , n6583 );
or ( n7002 , n6998 , n7001 );
xor ( n7003 , n6995 , n7002 );
buf ( n7004 , n4531 );
xor ( n7005 , n7003 , n7004 );
buf ( n7006 , n4532 );
xor ( n7007 , n7005 , n7006 );
buf ( n7008 , n4533 );
xor ( n7009 , n7007 , n7008 );
xor ( n7010 , n6988 , n7009 );
and ( n7011 , n6965 , n7010 );
xor ( n7012 , n6919 , n7011 );
xor ( n7013 , n6874 , n7012 );
buf ( n7014 , n4534 );
not ( n7015 , n6583 );
buf ( n7016 , n4535 );
and ( n7017 , n7015 , n7016 );
buf ( n7018 , n4536 );
xor ( n7019 , n7018 , n7016 );
and ( n7020 , n7019 , n6583 );
or ( n7021 , n7017 , n7020 );
buf ( n7022 , n4537 );
xor ( n7023 , n7021 , n7022 );
buf ( n7024 , n4538 );
xor ( n7025 , n7023 , n7024 );
buf ( n7026 , n4539 );
xor ( n7027 , n7025 , n7026 );
buf ( n7028 , n4540 );
xor ( n7029 , n7027 , n7028 );
xor ( n7030 , n7014 , n7029 );
not ( n7031 , n6583 );
buf ( n7032 , n4541 );
and ( n7033 , n7031 , n7032 );
buf ( n7034 , n4542 );
xor ( n7035 , n7034 , n7032 );
and ( n7036 , n7035 , n6583 );
or ( n7037 , n7033 , n7036 );
not ( n7038 , n6583 );
buf ( n7039 , n4543 );
and ( n7040 , n7038 , n7039 );
buf ( n7041 , n4544 );
xor ( n7042 , n7041 , n7039 );
and ( n7043 , n7042 , n6583 );
or ( n7044 , n7040 , n7043 );
xor ( n7045 , n7037 , n7044 );
buf ( n7046 , n4545 );
xor ( n7047 , n7045 , n7046 );
buf ( n7048 , n4546 );
xor ( n7049 , n7047 , n7048 );
buf ( n7050 , n4547 );
xor ( n7051 , n7049 , n7050 );
xor ( n7052 , n7030 , n7051 );
not ( n7053 , n6583 );
buf ( n7054 , n4548 );
and ( n7055 , n7053 , n7054 );
buf ( n7056 , n4549 );
xor ( n7057 , n7056 , n7054 );
and ( n7058 , n7057 , n6583 );
or ( n7059 , n7055 , n7058 );
not ( n7060 , n6583 );
buf ( n7061 , n4550 );
and ( n7062 , n7060 , n7061 );
buf ( n7063 , n4551 );
xor ( n7064 , n7063 , n7061 );
and ( n7065 , n7064 , n6583 );
or ( n7066 , n7062 , n7065 );
xor ( n7067 , n7059 , n7066 );
buf ( n7068 , n4552 );
xor ( n7069 , n7067 , n7068 );
buf ( n7070 , n4553 );
xor ( n7071 , n7069 , n7070 );
buf ( n7072 , n4554 );
xor ( n7073 , n7071 , n7072 );
xor ( n7074 , n6805 , n7073 );
not ( n7075 , n6583 );
buf ( n7076 , n4555 );
and ( n7077 , n7075 , n7076 );
buf ( n7078 , n4556 );
xor ( n7079 , n7078 , n7076 );
and ( n7080 , n7079 , n6583 );
or ( n7081 , n7077 , n7080 );
not ( n7082 , n6583 );
buf ( n7083 , n4557 );
and ( n7084 , n7082 , n7083 );
buf ( n7085 , n4558 );
xor ( n7086 , n7085 , n7083 );
and ( n7087 , n7086 , n6583 );
or ( n7088 , n7084 , n7087 );
xor ( n7089 , n7081 , n7088 );
buf ( n7090 , n4559 );
xor ( n7091 , n7089 , n7090 );
buf ( n7092 , n4560 );
xor ( n7093 , n7091 , n7092 );
buf ( n7094 , n4561 );
xor ( n7095 , n7093 , n7094 );
xor ( n7096 , n7074 , n7095 );
not ( n7097 , n7096 );
not ( n7098 , n6583 );
buf ( n7099 , n4562 );
and ( n7100 , n7098 , n7099 );
buf ( n7101 , n4563 );
xor ( n7102 , n7101 , n7099 );
and ( n7103 , n7102 , n6583 );
or ( n7104 , n7100 , n7103 );
not ( n7105 , n6583 );
buf ( n7106 , n4564 );
and ( n7107 , n7105 , n7106 );
buf ( n7108 , n4565 );
xor ( n7109 , n7108 , n7106 );
and ( n7110 , n7109 , n6583 );
or ( n7111 , n7107 , n7110 );
not ( n7112 , n6583 );
buf ( n7113 , n4566 );
and ( n7114 , n7112 , n7113 );
buf ( n7115 , n4567 );
xor ( n7116 , n7115 , n7113 );
and ( n7117 , n7116 , n6583 );
or ( n7118 , n7114 , n7117 );
xor ( n7119 , n7111 , n7118 );
buf ( n7120 , n4568 );
xor ( n7121 , n7119 , n7120 );
buf ( n7122 , n4569 );
xor ( n7123 , n7121 , n7122 );
buf ( n7124 , n4570 );
xor ( n7125 , n7123 , n7124 );
xor ( n7126 , n7104 , n7125 );
not ( n7127 , n6583 );
buf ( n7128 , n4571 );
and ( n7129 , n7127 , n7128 );
buf ( n7130 , n4572 );
xor ( n7131 , n7130 , n7128 );
and ( n7132 , n7131 , n6583 );
or ( n7133 , n7129 , n7132 );
not ( n7134 , n6583 );
buf ( n7135 , n4573 );
and ( n7136 , n7134 , n7135 );
buf ( n7137 , n4574 );
xor ( n7138 , n7137 , n7135 );
and ( n7139 , n7138 , n6583 );
or ( n7140 , n7136 , n7139 );
xor ( n7141 , n7133 , n7140 );
buf ( n7142 , n4575 );
xor ( n7143 , n7141 , n7142 );
buf ( n7144 , n4576 );
xor ( n7145 , n7143 , n7144 );
buf ( n7146 , n4577 );
xor ( n7147 , n7145 , n7146 );
xor ( n7148 , n7126 , n7147 );
and ( n7149 , n7097 , n7148 );
xor ( n7150 , n7052 , n7149 );
xor ( n7151 , n7013 , n7150 );
buf ( n7152 , n4578 );
not ( n7153 , n6583 );
buf ( n7154 , n4579 );
and ( n7155 , n7153 , n7154 );
buf ( n7156 , n4580 );
xor ( n7157 , n7156 , n7154 );
and ( n7158 , n7157 , n6583 );
or ( n7159 , n7155 , n7158 );
not ( n7160 , n6583 );
buf ( n7161 , n4581 );
and ( n7162 , n7160 , n7161 );
buf ( n7163 , n4582 );
xor ( n7164 , n7163 , n7161 );
and ( n7165 , n7164 , n6583 );
or ( n7166 , n7162 , n7165 );
xor ( n7167 , n7159 , n7166 );
buf ( n7168 , n4583 );
xor ( n7169 , n7167 , n7168 );
buf ( n7170 , n4584 );
xor ( n7171 , n7169 , n7170 );
buf ( n7172 , n4585 );
xor ( n7173 , n7171 , n7172 );
xor ( n7174 , n7152 , n7173 );
not ( n7175 , n6583 );
buf ( n7176 , n4586 );
and ( n7177 , n7175 , n7176 );
buf ( n7178 , n4587 );
xor ( n7179 , n7178 , n7176 );
and ( n7180 , n7179 , n6583 );
or ( n7181 , n7177 , n7180 );
buf ( n7182 , n4588 );
xor ( n7183 , n7181 , n7182 );
buf ( n7184 , n4589 );
xor ( n7185 , n7183 , n7184 );
buf ( n7186 , n4590 );
xor ( n7187 , n7185 , n7186 );
buf ( n7188 , n4591 );
xor ( n7189 , n7187 , n7188 );
xor ( n7190 , n7174 , n7189 );
not ( n7191 , n6637 );
and ( n7192 , n7191 , n6682 );
xor ( n7193 , n7190 , n7192 );
xor ( n7194 , n7151 , n7193 );
buf ( n7195 , n4592 );
not ( n7196 , n6583 );
buf ( n7197 , n4593 );
and ( n7198 , n7196 , n7197 );
buf ( n7199 , n4594 );
xor ( n7200 , n7199 , n7197 );
and ( n7201 , n7200 , n6583 );
or ( n7202 , n7198 , n7201 );
not ( n7203 , n6583 );
buf ( n7204 , n4595 );
and ( n7205 , n7203 , n7204 );
buf ( n7206 , n4596 );
xor ( n7207 , n7206 , n7204 );
and ( n7208 , n7207 , n6583 );
or ( n7209 , n7205 , n7208 );
xor ( n7210 , n7202 , n7209 );
buf ( n7211 , n4597 );
xor ( n7212 , n7210 , n7211 );
buf ( n7213 , n4598 );
xor ( n7214 , n7212 , n7213 );
buf ( n7215 , n4599 );
xor ( n7216 , n7214 , n7215 );
xor ( n7217 , n7195 , n7216 );
not ( n7218 , n6583 );
buf ( n7219 , n4600 );
and ( n7220 , n7218 , n7219 );
buf ( n7221 , n4601 );
xor ( n7222 , n7221 , n7219 );
and ( n7223 , n7222 , n6583 );
or ( n7224 , n7220 , n7223 );
not ( n7225 , n6583 );
buf ( n7226 , n4602 );
and ( n7227 , n7225 , n7226 );
buf ( n7228 , n4603 );
xor ( n7229 , n7228 , n7226 );
and ( n7230 , n7229 , n6583 );
or ( n7231 , n7227 , n7230 );
xor ( n7232 , n7224 , n7231 );
buf ( n7233 , n4604 );
xor ( n7234 , n7232 , n7233 );
buf ( n7235 , n4605 );
xor ( n7236 , n7234 , n7235 );
buf ( n7237 , n4606 );
xor ( n7238 , n7236 , n7237 );
xor ( n7239 , n7217 , n7238 );
not ( n7240 , n6583 );
buf ( n7241 , n4607 );
and ( n7242 , n7240 , n7241 );
buf ( n7243 , n4608 );
xor ( n7244 , n7243 , n7241 );
and ( n7245 , n7244 , n6583 );
or ( n7246 , n7242 , n7245 );
not ( n7247 , n6583 );
buf ( n7248 , n4609 );
and ( n7249 , n7247 , n7248 );
buf ( n7250 , n4610 );
xor ( n7251 , n7250 , n7248 );
and ( n7252 , n7251 , n6583 );
or ( n7253 , n7249 , n7252 );
not ( n7254 , n6583 );
buf ( n7255 , n4611 );
and ( n7256 , n7254 , n7255 );
buf ( n7257 , n4612 );
xor ( n7258 , n7257 , n7255 );
and ( n7259 , n7258 , n6583 );
or ( n7260 , n7256 , n7259 );
xor ( n7261 , n7253 , n7260 );
buf ( n7262 , n4613 );
xor ( n7263 , n7261 , n7262 );
buf ( n7264 , n4614 );
xor ( n7265 , n7263 , n7264 );
buf ( n7266 , n4615 );
xor ( n7267 , n7265 , n7266 );
xor ( n7268 , n7246 , n7267 );
not ( n7269 , n6583 );
buf ( n7270 , n4616 );
and ( n7271 , n7269 , n7270 );
buf ( n7272 , n4617 );
xor ( n7273 , n7272 , n7270 );
and ( n7274 , n7273 , n6583 );
or ( n7275 , n7271 , n7274 );
not ( n7276 , n6583 );
buf ( n7277 , n4618 );
and ( n7278 , n7276 , n7277 );
buf ( n7279 , n4619 );
xor ( n7280 , n7279 , n7277 );
and ( n7281 , n7280 , n6583 );
or ( n7282 , n7278 , n7281 );
xor ( n7283 , n7275 , n7282 );
buf ( n7284 , n4620 );
xor ( n7285 , n7283 , n7284 );
buf ( n7286 , n4621 );
xor ( n7287 , n7285 , n7286 );
buf ( n7288 , n4622 );
xor ( n7289 , n7287 , n7288 );
xor ( n7290 , n7268 , n7289 );
not ( n7291 , n7290 );
not ( n7292 , n6583 );
buf ( n7293 , n4623 );
and ( n7294 , n7292 , n7293 );
buf ( n7295 , n4624 );
xor ( n7296 , n7295 , n7293 );
and ( n7297 , n7296 , n6583 );
or ( n7298 , n7294 , n7297 );
not ( n7299 , n6583 );
buf ( n7300 , n4625 );
and ( n7301 , n7299 , n7300 );
buf ( n7302 , n4626 );
xor ( n7303 , n7302 , n7300 );
and ( n7304 , n7303 , n6583 );
or ( n7305 , n7301 , n7304 );
not ( n7306 , n6583 );
buf ( n7307 , n4627 );
and ( n7308 , n7306 , n7307 );
buf ( n7309 , n4628 );
xor ( n7310 , n7309 , n7307 );
and ( n7311 , n7310 , n6583 );
or ( n7312 , n7308 , n7311 );
xor ( n7313 , n7305 , n7312 );
buf ( n7314 , n4629 );
xor ( n7315 , n7313 , n7314 );
buf ( n7316 , n4630 );
xor ( n7317 , n7315 , n7316 );
buf ( n7318 , n4631 );
xor ( n7319 , n7317 , n7318 );
xor ( n7320 , n7298 , n7319 );
not ( n7321 , n6583 );
buf ( n7322 , n4632 );
and ( n7323 , n7321 , n7322 );
buf ( n7324 , n4633 );
xor ( n7325 , n7324 , n7322 );
and ( n7326 , n7325 , n6583 );
or ( n7327 , n7323 , n7326 );
buf ( n7328 , n4634 );
xor ( n7329 , n7327 , n7328 );
buf ( n7330 , n4635 );
xor ( n7331 , n7329 , n7330 );
buf ( n7332 , n4636 );
xor ( n7333 , n7331 , n7332 );
buf ( n7334 , n4637 );
xor ( n7335 , n7333 , n7334 );
xor ( n7336 , n7320 , n7335 );
and ( n7337 , n7291 , n7336 );
xor ( n7338 , n7239 , n7337 );
xor ( n7339 , n7194 , n7338 );
xor ( n7340 , n6730 , n7339 );
not ( n7341 , n6583 );
buf ( n7342 , n4638 );
and ( n7343 , n7341 , n7342 );
buf ( n7344 , n4639 );
xor ( n7345 , n7344 , n7342 );
and ( n7346 , n7345 , n6583 );
or ( n7347 , n7343 , n7346 );
not ( n7348 , n6583 );
buf ( n7349 , n4640 );
and ( n7350 , n7348 , n7349 );
buf ( n7351 , n4641 );
xor ( n7352 , n7351 , n7349 );
and ( n7353 , n7352 , n6583 );
or ( n7354 , n7350 , n7353 );
not ( n7355 , n6583 );
buf ( n7356 , n4642 );
and ( n7357 , n7355 , n7356 );
buf ( n7358 , n4643 );
xor ( n7359 , n7358 , n7356 );
and ( n7360 , n7359 , n6583 );
or ( n7361 , n7357 , n7360 );
xor ( n7362 , n7354 , n7361 );
buf ( n7363 , n4644 );
xor ( n7364 , n7362 , n7363 );
buf ( n7365 , n4645 );
xor ( n7366 , n7364 , n7365 );
buf ( n7367 , n4646 );
xor ( n7368 , n7366 , n7367 );
xor ( n7369 , n7347 , n7368 );
not ( n7370 , n6583 );
buf ( n7371 , n4647 );
and ( n7372 , n7370 , n7371 );
buf ( n7373 , n4648 );
xor ( n7374 , n7373 , n7371 );
and ( n7375 , n7374 , n6583 );
or ( n7376 , n7372 , n7375 );
not ( n7377 , n6583 );
buf ( n7378 , n4649 );
and ( n7379 , n7377 , n7378 );
buf ( n7380 , n4650 );
xor ( n7381 , n7380 , n7378 );
and ( n7382 , n7381 , n6583 );
or ( n7383 , n7379 , n7382 );
xor ( n7384 , n7376 , n7383 );
buf ( n7385 , n4651 );
xor ( n7386 , n7384 , n7385 );
buf ( n7387 , n4652 );
xor ( n7388 , n7386 , n7387 );
buf ( n7389 , n4653 );
xor ( n7390 , n7388 , n7389 );
xor ( n7391 , n7369 , n7390 );
buf ( n7392 , n4654 );
not ( n7393 , n6583 );
buf ( n7394 , n4655 );
and ( n7395 , n7393 , n7394 );
buf ( n7396 , n4656 );
xor ( n7397 , n7396 , n7394 );
and ( n7398 , n7397 , n6583 );
or ( n7399 , n7395 , n7398 );
xor ( n7400 , n7399 , n6828 );
buf ( n7401 , n4657 );
xor ( n7402 , n7400 , n7401 );
buf ( n7403 , n4658 );
xor ( n7404 , n7402 , n7403 );
buf ( n7405 , n4659 );
xor ( n7406 , n7404 , n7405 );
xor ( n7407 , n7392 , n7406 );
not ( n7408 , n6583 );
buf ( n7409 , n4660 );
and ( n7410 , n7408 , n7409 );
buf ( n7411 , n4661 );
xor ( n7412 , n7411 , n7409 );
and ( n7413 , n7412 , n6583 );
or ( n7414 , n7410 , n7413 );
not ( n7415 , n6583 );
buf ( n7416 , n4662 );
and ( n7417 , n7415 , n7416 );
buf ( n7418 , n4663 );
xor ( n7419 , n7418 , n7416 );
and ( n7420 , n7419 , n6583 );
or ( n7421 , n7417 , n7420 );
xor ( n7422 , n7414 , n7421 );
buf ( n7423 , n4664 );
xor ( n7424 , n7422 , n7423 );
buf ( n7425 , n4665 );
xor ( n7426 , n7424 , n7425 );
buf ( n7427 , n4666 );
xor ( n7428 , n7426 , n7427 );
xor ( n7429 , n7407 , n7428 );
not ( n7430 , n7429 );
buf ( n7431 , n4667 );
not ( n7432 , n6583 );
buf ( n7433 , n4668 );
and ( n7434 , n7432 , n7433 );
buf ( n7435 , n4669 );
xor ( n7436 , n7435 , n7433 );
and ( n7437 , n7436 , n6583 );
or ( n7438 , n7434 , n7437 );
not ( n7439 , n6583 );
buf ( n7440 , n4670 );
and ( n7441 , n7439 , n7440 );
buf ( n7442 , n4671 );
xor ( n7443 , n7442 , n7440 );
and ( n7444 , n7443 , n6583 );
or ( n7445 , n7441 , n7444 );
xor ( n7446 , n7438 , n7445 );
buf ( n7447 , n4672 );
xor ( n7448 , n7446 , n7447 );
buf ( n7449 , n4673 );
xor ( n7450 , n7448 , n7449 );
buf ( n7451 , n4674 );
xor ( n7452 , n7450 , n7451 );
xor ( n7453 , n7431 , n7452 );
not ( n7454 , n6583 );
buf ( n7455 , n4675 );
and ( n7456 , n7454 , n7455 );
buf ( n7457 , n4676 );
xor ( n7458 , n7457 , n7455 );
and ( n7459 , n7458 , n6583 );
or ( n7460 , n7456 , n7459 );
buf ( n7461 , n4677 );
xor ( n7462 , n7460 , n7461 );
buf ( n7463 , n4678 );
xor ( n7464 , n7462 , n7463 );
buf ( n7465 , n4679 );
xor ( n7466 , n7464 , n7465 );
buf ( n7467 , n4680 );
buf ( n7468 , n7467 );
xor ( n7469 , n7466 , n7468 );
xor ( n7470 , n7453 , n7469 );
and ( n7471 , n7430 , n7470 );
xor ( n7472 , n7391 , n7471 );
buf ( n7473 , n4681 );
not ( n7474 , n6583 );
buf ( n7475 , n4682 );
and ( n7476 , n7474 , n7475 );
buf ( n7477 , n4683 );
xor ( n7478 , n7477 , n7475 );
and ( n7479 , n7478 , n6583 );
or ( n7480 , n7476 , n7479 );
not ( n7481 , n6583 );
buf ( n7482 , n4684 );
and ( n7483 , n7481 , n7482 );
buf ( n7484 , n4685 );
xor ( n7485 , n7484 , n7482 );
and ( n7486 , n7485 , n6583 );
or ( n7487 , n7483 , n7486 );
xor ( n7488 , n7480 , n7487 );
buf ( n7489 , n4686 );
xor ( n7490 , n7488 , n7489 );
buf ( n7491 , n4687 );
xor ( n7492 , n7490 , n7491 );
buf ( n7493 , n4688 );
xor ( n7494 , n7492 , n7493 );
xor ( n7495 , n7473 , n7494 );
not ( n7496 , n6583 );
buf ( n7497 , n4689 );
and ( n7498 , n7496 , n7497 );
buf ( n7499 , n4690 );
xor ( n7500 , n7499 , n7497 );
and ( n7501 , n7500 , n6583 );
or ( n7502 , n7498 , n7501 );
not ( n7503 , n6583 );
buf ( n7504 , n4691 );
and ( n7505 , n7503 , n7504 );
buf ( n7506 , n4692 );
xor ( n7507 , n7506 , n7504 );
and ( n7508 , n7507 , n6583 );
or ( n7509 , n7505 , n7508 );
xor ( n7510 , n7502 , n7509 );
buf ( n7511 , n4693 );
xor ( n7512 , n7510 , n7511 );
buf ( n7513 , n4694 );
xor ( n7514 , n7512 , n7513 );
buf ( n7515 , n4695 );
xor ( n7516 , n7514 , n7515 );
xor ( n7517 , n7495 , n7516 );
buf ( n7518 , n4696 );
not ( n7519 , n6583 );
buf ( n7520 , n4697 );
and ( n7521 , n7519 , n7520 );
buf ( n7522 , n4698 );
xor ( n7523 , n7522 , n7520 );
and ( n7524 , n7523 , n6583 );
or ( n7525 , n7521 , n7524 );
buf ( n7526 , n4699 );
xor ( n7527 , n7525 , n7526 );
buf ( n7528 , n4700 );
xor ( n7529 , n7527 , n7528 );
buf ( n7530 , n4701 );
xor ( n7531 , n7529 , n7530 );
buf ( n7532 , n4702 );
xor ( n7533 , n7531 , n7532 );
xor ( n7534 , n7518 , n7533 );
not ( n7535 , n6583 );
buf ( n7536 , n4703 );
and ( n7537 , n7535 , n7536 );
buf ( n7538 , n4704 );
xor ( n7539 , n7538 , n7536 );
and ( n7540 , n7539 , n6583 );
or ( n7541 , n7537 , n7540 );
not ( n7542 , n6583 );
buf ( n7543 , n4705 );
and ( n7544 , n7542 , n7543 );
buf ( n7545 , n4706 );
xor ( n7546 , n7545 , n7543 );
and ( n7547 , n7546 , n6583 );
or ( n7548 , n7544 , n7547 );
xor ( n7549 , n7541 , n7548 );
buf ( n7550 , n4707 );
xor ( n7551 , n7549 , n7550 );
buf ( n7552 , n4708 );
xor ( n7553 , n7551 , n7552 );
buf ( n7554 , n4709 );
xor ( n7555 , n7553 , n7554 );
xor ( n7556 , n7534 , n7555 );
not ( n7557 , n7556 );
buf ( n7558 , n4710 );
not ( n7559 , n6583 );
buf ( n7560 , n4711 );
and ( n7561 , n7559 , n7560 );
buf ( n7562 , n4712 );
xor ( n7563 , n7562 , n7560 );
and ( n7564 , n7563 , n6583 );
or ( n7565 , n7561 , n7564 );
not ( n7566 , n6583 );
buf ( n7567 , n4713 );
and ( n7568 , n7566 , n7567 );
buf ( n7569 , n4714 );
xor ( n7570 , n7569 , n7567 );
and ( n7571 , n7570 , n6583 );
or ( n7572 , n7568 , n7571 );
xor ( n7573 , n7565 , n7572 );
buf ( n7574 , n4715 );
xor ( n7575 , n7573 , n7574 );
buf ( n7576 , n4716 );
xor ( n7577 , n7575 , n7576 );
buf ( n7578 , n4717 );
xor ( n7579 , n7577 , n7578 );
xor ( n7580 , n7558 , n7579 );
not ( n7581 , n6583 );
buf ( n7582 , n4718 );
and ( n7583 , n7581 , n7582 );
buf ( n7584 , n4719 );
xor ( n7585 , n7584 , n7582 );
and ( n7586 , n7585 , n6583 );
or ( n7587 , n7583 , n7586 );
not ( n7588 , n6583 );
buf ( n7589 , n4720 );
and ( n7590 , n7588 , n7589 );
buf ( n7591 , n4721 );
xor ( n7592 , n7591 , n7589 );
and ( n7593 , n7592 , n6583 );
or ( n7594 , n7590 , n7593 );
xor ( n7595 , n7587 , n7594 );
buf ( n7596 , n7595 );
buf ( n7597 , n4722 );
xor ( n7598 , n7596 , n7597 );
buf ( n7599 , n4723 );
xor ( n7600 , n7598 , n7599 );
xor ( n7601 , n7580 , n7600 );
and ( n7602 , n7557 , n7601 );
xor ( n7603 , n7517 , n7602 );
xor ( n7604 , n7472 , n7603 );
not ( n7605 , n6583 );
buf ( n7606 , n4724 );
and ( n7607 , n7605 , n7606 );
buf ( n7608 , n4725 );
xor ( n7609 , n7608 , n7606 );
and ( n7610 , n7609 , n6583 );
or ( n7611 , n7607 , n7610 );
not ( n7612 , n6583 );
buf ( n7613 , n4726 );
and ( n7614 , n7612 , n7613 );
buf ( n7615 , n4727 );
xor ( n7616 , n7615 , n7613 );
and ( n7617 , n7616 , n6583 );
or ( n7618 , n7614 , n7617 );
not ( n7619 , n6583 );
buf ( n7620 , n4728 );
and ( n7621 , n7619 , n7620 );
buf ( n7622 , n4729 );
xor ( n7623 , n7622 , n7620 );
and ( n7624 , n7623 , n6583 );
or ( n7625 , n7621 , n7624 );
xor ( n7626 , n7618 , n7625 );
buf ( n7627 , n4730 );
xor ( n7628 , n7626 , n7627 );
buf ( n7629 , n4731 );
xor ( n7630 , n7628 , n7629 );
buf ( n7631 , n4732 );
xor ( n7632 , n7630 , n7631 );
xor ( n7633 , n7611 , n7632 );
not ( n7634 , n6583 );
buf ( n7635 , n4733 );
and ( n7636 , n7634 , n7635 );
buf ( n7637 , n4734 );
xor ( n7638 , n7637 , n7635 );
and ( n7639 , n7638 , n6583 );
or ( n7640 , n7636 , n7639 );
not ( n7641 , n6583 );
buf ( n7642 , n4735 );
and ( n7643 , n7641 , n7642 );
buf ( n7644 , n4736 );
xor ( n7645 , n7644 , n7642 );
and ( n7646 , n7645 , n6583 );
or ( n7647 , n7643 , n7646 );
xor ( n7648 , n7640 , n7647 );
buf ( n7649 , n4737 );
xor ( n7650 , n7648 , n7649 );
buf ( n7651 , n4738 );
xor ( n7652 , n7650 , n7651 );
buf ( n7653 , n4739 );
xor ( n7654 , n7652 , n7653 );
xor ( n7655 , n7633 , n7654 );
buf ( n7656 , n4740 );
not ( n7657 , n6583 );
buf ( n7658 , n4741 );
and ( n7659 , n7657 , n7658 );
buf ( n7660 , n4742 );
xor ( n7661 , n7660 , n7658 );
and ( n7662 , n7661 , n6583 );
or ( n7663 , n7659 , n7662 );
not ( n7664 , n6583 );
buf ( n7665 , n4743 );
and ( n7666 , n7664 , n7665 );
buf ( n7667 , n4744 );
xor ( n7668 , n7667 , n7665 );
and ( n7669 , n7668 , n6583 );
or ( n7670 , n7666 , n7669 );
xor ( n7671 , n7663 , n7670 );
buf ( n7672 , n4745 );
xor ( n7673 , n7671 , n7672 );
buf ( n7674 , n4746 );
xor ( n7675 , n7673 , n7674 );
buf ( n7676 , n4747 );
xor ( n7677 , n7675 , n7676 );
xor ( n7678 , n7656 , n7677 );
buf ( n7679 , n4748 );
xor ( n7680 , n6594 , n7679 );
buf ( n7681 , n4749 );
xor ( n7682 , n7680 , n7681 );
buf ( n7683 , n4750 );
xor ( n7684 , n7682 , n7683 );
buf ( n7685 , n4751 );
xor ( n7686 , n7684 , n7685 );
xor ( n7687 , n7678 , n7686 );
not ( n7688 , n7687 );
buf ( n7689 , n4752 );
not ( n7690 , n6583 );
buf ( n7691 , n4753 );
and ( n7692 , n7690 , n7691 );
buf ( n7693 , n4754 );
xor ( n7694 , n7693 , n7691 );
and ( n7695 , n7694 , n6583 );
or ( n7696 , n7692 , n7695 );
not ( n7697 , n6583 );
buf ( n7698 , n4755 );
and ( n7699 , n7697 , n7698 );
buf ( n7700 , n4756 );
xor ( n7701 , n7700 , n7698 );
and ( n7702 , n7701 , n6583 );
or ( n7703 , n7699 , n7702 );
xor ( n7704 , n7696 , n7703 );
buf ( n7705 , n4757 );
xor ( n7706 , n7704 , n7705 );
buf ( n7707 , n4758 );
xor ( n7708 , n7706 , n7707 );
buf ( n7709 , n4759 );
xor ( n7710 , n7708 , n7709 );
xor ( n7711 , n7689 , n7710 );
xor ( n7712 , n7711 , n6705 );
and ( n7713 , n7688 , n7712 );
xor ( n7714 , n7655 , n7713 );
xor ( n7715 , n7604 , n7714 );
not ( n7716 , n6583 );
buf ( n7717 , n4760 );
and ( n7718 , n7716 , n7717 );
buf ( n7719 , n4761 );
xor ( n7720 , n7719 , n7717 );
and ( n7721 , n7720 , n6583 );
or ( n7722 , n7718 , n7721 );
not ( n7723 , n6583 );
buf ( n7724 , n4762 );
and ( n7725 , n7723 , n7724 );
buf ( n7726 , n4763 );
xor ( n7727 , n7726 , n7724 );
and ( n7728 , n7727 , n6583 );
or ( n7729 , n7725 , n7728 );
buf ( n7730 , n4764 );
xor ( n7731 , n7729 , n7730 );
buf ( n7732 , n4765 );
xor ( n7733 , n7731 , n7732 );
buf ( n7734 , n4766 );
xor ( n7735 , n7733 , n7734 );
buf ( n7736 , n4767 );
xor ( n7737 , n7735 , n7736 );
xor ( n7738 , n7722 , n7737 );
not ( n7739 , n6583 );
buf ( n7740 , n4768 );
and ( n7741 , n7739 , n7740 );
buf ( n7742 , n4769 );
xor ( n7743 , n7742 , n7740 );
and ( n7744 , n7743 , n6583 );
or ( n7745 , n7741 , n7744 );
not ( n7746 , n6583 );
buf ( n7747 , n4770 );
and ( n7748 , n7746 , n7747 );
buf ( n7749 , n4771 );
xor ( n7750 , n7749 , n7747 );
and ( n7751 , n7750 , n6583 );
or ( n7752 , n7748 , n7751 );
xor ( n7753 , n7745 , n7752 );
buf ( n7754 , n4772 );
xor ( n7755 , n7753 , n7754 );
buf ( n7756 , n4773 );
xor ( n7757 , n7755 , n7756 );
buf ( n7758 , n4774 );
xor ( n7759 , n7757 , n7758 );
xor ( n7760 , n7738 , n7759 );
buf ( n7761 , n4775 );
not ( n7762 , n6583 );
buf ( n7763 , n4776 );
and ( n7764 , n7762 , n7763 );
buf ( n7765 , n4777 );
xor ( n7766 , n7765 , n7763 );
and ( n7767 , n7766 , n6583 );
or ( n7768 , n7764 , n7767 );
not ( n7769 , n6583 );
buf ( n7770 , n4778 );
and ( n7771 , n7769 , n7770 );
buf ( n7772 , n4779 );
xor ( n7773 , n7772 , n7770 );
and ( n7774 , n7773 , n6583 );
or ( n7775 , n7771 , n7774 );
xor ( n7776 , n7768 , n7775 );
buf ( n7777 , n4780 );
xor ( n7778 , n7776 , n7777 );
buf ( n7779 , n4781 );
xor ( n7780 , n7778 , n7779 );
buf ( n7781 , n4782 );
xor ( n7782 , n7780 , n7781 );
xor ( n7783 , n7761 , n7782 );
not ( n7784 , n6583 );
buf ( n7785 , n4783 );
and ( n7786 , n7784 , n7785 );
buf ( n7787 , n4784 );
xor ( n7788 , n7787 , n7785 );
and ( n7789 , n7788 , n6583 );
or ( n7790 , n7786 , n7789 );
not ( n7791 , n6583 );
buf ( n7792 , n4785 );
and ( n7793 , n7791 , n7792 );
buf ( n7794 , n4786 );
xor ( n7795 , n7794 , n7792 );
and ( n7796 , n7795 , n6583 );
or ( n7797 , n7793 , n7796 );
xor ( n7798 , n7790 , n7797 );
buf ( n7799 , n4787 );
xor ( n7800 , n7798 , n7799 );
buf ( n7801 , n4788 );
xor ( n7802 , n7800 , n7801 );
buf ( n7803 , n4789 );
xor ( n7804 , n7802 , n7803 );
xor ( n7805 , n7783 , n7804 );
not ( n7806 , n7805 );
buf ( n7807 , n4790 );
not ( n7808 , n6583 );
buf ( n7809 , n4791 );
and ( n7810 , n7808 , n7809 );
buf ( n7811 , n4792 );
xor ( n7812 , n7811 , n7809 );
and ( n7813 , n7812 , n6583 );
or ( n7814 , n7810 , n7813 );
not ( n7815 , n6583 );
buf ( n7816 , n4793 );
and ( n7817 , n7815 , n7816 );
buf ( n7818 , n4794 );
xor ( n7819 , n7818 , n7816 );
and ( n7820 , n7819 , n6583 );
or ( n7821 , n7817 , n7820 );
xor ( n7822 , n7814 , n7821 );
buf ( n7823 , n4795 );
xor ( n7824 , n7822 , n7823 );
buf ( n7825 , n4796 );
xor ( n7826 , n7824 , n7825 );
buf ( n7827 , n4797 );
xor ( n7828 , n7826 , n7827 );
xor ( n7829 , n7807 , n7828 );
not ( n7830 , n6583 );
buf ( n7831 , n4798 );
and ( n7832 , n7830 , n7831 );
buf ( n7833 , n4799 );
xor ( n7834 , n7833 , n7831 );
and ( n7835 , n7834 , n6583 );
or ( n7836 , n7832 , n7835 );
not ( n7837 , n6583 );
buf ( n7838 , n4800 );
and ( n7839 , n7837 , n7838 );
buf ( n7840 , n4801 );
xor ( n7841 , n7840 , n7838 );
and ( n7842 , n7841 , n6583 );
or ( n7843 , n7839 , n7842 );
xor ( n7844 , n7836 , n7843 );
buf ( n7845 , n4802 );
buf ( n7846 , n7845 );
xor ( n7847 , n7844 , n7846 );
buf ( n7848 , n4803 );
xor ( n7849 , n7847 , n7848 );
buf ( n7850 , n4804 );
xor ( n7851 , n7849 , n7850 );
xor ( n7852 , n7829 , n7851 );
and ( n7853 , n7806 , n7852 );
xor ( n7854 , n7760 , n7853 );
xor ( n7855 , n7715 , n7854 );
not ( n7856 , n6583 );
buf ( n7857 , n4805 );
and ( n7858 , n7856 , n7857 );
buf ( n7859 , n4806 );
xor ( n7860 , n7859 , n7857 );
and ( n7861 , n7860 , n6583 );
or ( n7862 , n7858 , n7861 );
xor ( n7863 , n7862 , n7173 );
xor ( n7864 , n7863 , n7189 );
buf ( n7865 , n4807 );
not ( n7866 , n6583 );
buf ( n7867 , n4808 );
and ( n7868 , n7866 , n7867 );
buf ( n7869 , n4809 );
xor ( n7870 , n7869 , n7867 );
and ( n7871 , n7870 , n6583 );
or ( n7872 , n7868 , n7871 );
not ( n7873 , n6583 );
buf ( n7874 , n4810 );
and ( n7875 , n7873 , n7874 );
buf ( n7876 , n4811 );
xor ( n7877 , n7876 , n7874 );
and ( n7878 , n7877 , n6583 );
or ( n7879 , n7875 , n7878 );
xor ( n7880 , n7872 , n7879 );
buf ( n7881 , n4812 );
xor ( n7882 , n7880 , n7881 );
buf ( n7883 , n4813 );
xor ( n7884 , n7882 , n7883 );
buf ( n7885 , n4814 );
xor ( n7886 , n7884 , n7885 );
xor ( n7887 , n7865 , n7886 );
not ( n7888 , n6583 );
buf ( n7889 , n4815 );
and ( n7890 , n7888 , n7889 );
buf ( n7891 , n4816 );
xor ( n7892 , n7891 , n7889 );
and ( n7893 , n7892 , n6583 );
or ( n7894 , n7890 , n7893 );
not ( n7895 , n6583 );
buf ( n7896 , n4817 );
and ( n7897 , n7895 , n7896 );
buf ( n7898 , n4818 );
xor ( n7899 , n7898 , n7896 );
and ( n7900 , n7899 , n6583 );
or ( n7901 , n7897 , n7900 );
xor ( n7902 , n7894 , n7901 );
buf ( n7903 , n4819 );
xor ( n7904 , n7902 , n7903 );
buf ( n7905 , n4820 );
xor ( n7906 , n7904 , n7905 );
buf ( n7907 , n4821 );
xor ( n7908 , n7906 , n7907 );
xor ( n7909 , n7887 , n7908 );
not ( n7910 , n7909 );
buf ( n7911 , n4822 );
not ( n7912 , n6583 );
buf ( n7913 , n4823 );
and ( n7914 , n7912 , n7913 );
buf ( n7915 , n4824 );
xor ( n7916 , n7915 , n7913 );
and ( n7917 , n7916 , n6583 );
or ( n7918 , n7914 , n7917 );
buf ( n7919 , n4825 );
xor ( n7920 , n7918 , n7919 );
buf ( n7921 , n4826 );
xor ( n7922 , n7920 , n7921 );
buf ( n7923 , n4827 );
xor ( n7924 , n7922 , n7923 );
buf ( n7925 , n4828 );
xor ( n7926 , n7924 , n7925 );
xor ( n7927 , n7911 , n7926 );
not ( n7928 , n6583 );
buf ( n7929 , n4829 );
and ( n7930 , n7928 , n7929 );
buf ( n7931 , n4830 );
xor ( n7932 , n7931 , n7929 );
and ( n7933 , n7932 , n6583 );
or ( n7934 , n7930 , n7933 );
not ( n7935 , n6583 );
buf ( n7936 , n4831 );
and ( n7937 , n7935 , n7936 );
buf ( n7938 , n4832 );
xor ( n7939 , n7938 , n7936 );
and ( n7940 , n7939 , n6583 );
or ( n7941 , n7937 , n7940 );
xor ( n7942 , n7934 , n7941 );
buf ( n7943 , n4833 );
xor ( n7944 , n7942 , n7943 );
buf ( n7945 , n4834 );
xor ( n7946 , n7944 , n7945 );
buf ( n7947 , n4835 );
xor ( n7948 , n7946 , n7947 );
xor ( n7949 , n7927 , n7948 );
and ( n7950 , n7910 , n7949 );
xor ( n7951 , n7864 , n7950 );
xor ( n7952 , n7855 , n7951 );
xor ( n7953 , n7340 , n7952 );
not ( n7954 , n6583 );
buf ( n7955 , n4836 );
and ( n7956 , n7954 , n7955 );
buf ( n7957 , n4837 );
xor ( n7958 , n7957 , n7955 );
and ( n7959 , n7958 , n6583 );
or ( n7960 , n7956 , n7959 );
not ( n7961 , n6583 );
buf ( n7962 , n4838 );
and ( n7963 , n7961 , n7962 );
buf ( n7964 , n4839 );
xor ( n7965 , n7964 , n7962 );
and ( n7966 , n7965 , n6583 );
or ( n7967 , n7963 , n7966 );
not ( n7968 , n6583 );
buf ( n7969 , n4840 );
and ( n7970 , n7968 , n7969 );
buf ( n7971 , n4841 );
xor ( n7972 , n7971 , n7969 );
and ( n7973 , n7972 , n6583 );
or ( n7974 , n7970 , n7973 );
xor ( n7975 , n7967 , n7974 );
buf ( n7976 , n4842 );
xor ( n7977 , n7975 , n7976 );
xor ( n7978 , n7977 , n7807 );
buf ( n7979 , n4843 );
xor ( n7980 , n7978 , n7979 );
xor ( n7981 , n7960 , n7980 );
not ( n7982 , n6583 );
buf ( n7983 , n4844 );
and ( n7984 , n7982 , n7983 );
buf ( n7985 , n4845 );
xor ( n7986 , n7985 , n7983 );
and ( n7987 , n7986 , n6583 );
or ( n7988 , n7984 , n7987 );
buf ( n7989 , n4846 );
xor ( n7990 , n7988 , n7989 );
buf ( n7991 , n4847 );
xor ( n7992 , n7990 , n7991 );
buf ( n7993 , n4848 );
xor ( n7994 , n7992 , n7993 );
buf ( n7995 , n4849 );
xor ( n7996 , n7994 , n7995 );
xor ( n7997 , n7981 , n7996 );
not ( n7998 , n6583 );
buf ( n7999 , n4850 );
and ( n8000 , n7998 , n7999 );
buf ( n8001 , n4851 );
xor ( n8002 , n8001 , n7999 );
and ( n8003 , n8002 , n6583 );
or ( n8004 , n8000 , n8003 );
not ( n8005 , n6583 );
buf ( n8006 , n4852 );
and ( n8007 , n8005 , n8006 );
buf ( n8008 , n4853 );
xor ( n8009 , n8008 , n8006 );
and ( n8010 , n8009 , n6583 );
or ( n8011 , n8007 , n8010 );
xor ( n8012 , n8004 , n8011 );
buf ( n8013 , n4854 );
xor ( n8014 , n8012 , n8013 );
buf ( n8015 , n4855 );
xor ( n8016 , n8014 , n8015 );
buf ( n8017 , n4856 );
xor ( n8018 , n8016 , n8017 );
xor ( n8019 , n6792 , n8018 );
xor ( n8020 , n8019 , n7073 );
not ( n8021 , n8020 );
not ( n8022 , n6583 );
buf ( n8023 , n4857 );
and ( n8024 , n8022 , n8023 );
buf ( n8025 , n4858 );
xor ( n8026 , n8025 , n8023 );
and ( n8027 , n8026 , n6583 );
or ( n8028 , n8024 , n8027 );
buf ( n8029 , n4859 );
xor ( n8030 , n8028 , n8029 );
buf ( n8031 , n4860 );
xor ( n8032 , n8030 , n8031 );
buf ( n8033 , n4861 );
xor ( n8034 , n8032 , n8033 );
buf ( n8035 , n4862 );
xor ( n8036 , n8034 , n8035 );
xor ( n8037 , n7213 , n8036 );
not ( n8038 , n6583 );
buf ( n8039 , n4863 );
and ( n8040 , n8038 , n8039 );
buf ( n8041 , n4864 );
xor ( n8042 , n8041 , n8039 );
and ( n8043 , n8042 , n6583 );
or ( n8044 , n8040 , n8043 );
not ( n8045 , n6583 );
buf ( n8046 , n4865 );
and ( n8047 , n8045 , n8046 );
buf ( n8048 , n4866 );
xor ( n8049 , n8048 , n8046 );
and ( n8050 , n8049 , n6583 );
or ( n8051 , n8047 , n8050 );
xor ( n8052 , n8044 , n8051 );
buf ( n8053 , n4867 );
xor ( n8054 , n8052 , n8053 );
buf ( n8055 , n4868 );
xor ( n8056 , n8054 , n8055 );
buf ( n8057 , n4869 );
xor ( n8058 , n8056 , n8057 );
xor ( n8059 , n8037 , n8058 );
and ( n8060 , n8021 , n8059 );
xor ( n8061 , n7997 , n8060 );
not ( n8062 , n6583 );
buf ( n8063 , n4870 );
and ( n8064 , n8062 , n8063 );
buf ( n8065 , n4871 );
xor ( n8066 , n8065 , n8063 );
and ( n8067 , n8066 , n6583 );
or ( n8068 , n8064 , n8067 );
not ( n8069 , n6583 );
buf ( n8070 , n4872 );
and ( n8071 , n8069 , n8070 );
buf ( n8072 , n4873 );
xor ( n8073 , n8072 , n8070 );
and ( n8074 , n8073 , n6583 );
or ( n8075 , n8071 , n8074 );
buf ( n8076 , n4874 );
xor ( n8077 , n8075 , n8076 );
buf ( n8078 , n4875 );
xor ( n8079 , n8077 , n8078 );
buf ( n8080 , n4876 );
xor ( n8081 , n8079 , n8080 );
buf ( n8082 , n4877 );
xor ( n8083 , n8081 , n8082 );
xor ( n8084 , n8068 , n8083 );
not ( n8085 , n6583 );
buf ( n8086 , n4878 );
and ( n8087 , n8085 , n8086 );
buf ( n8088 , n4879 );
xor ( n8089 , n8088 , n8086 );
and ( n8090 , n8089 , n6583 );
or ( n8091 , n8087 , n8090 );
not ( n8092 , n6583 );
buf ( n8093 , n4880 );
and ( n8094 , n8092 , n8093 );
buf ( n8095 , n4881 );
xor ( n8096 , n8095 , n8093 );
and ( n8097 , n8096 , n6583 );
or ( n8098 , n8094 , n8097 );
xor ( n8099 , n8091 , n8098 );
buf ( n8100 , n4882 );
xor ( n8101 , n8099 , n8100 );
buf ( n8102 , n4883 );
xor ( n8103 , n8101 , n8102 );
buf ( n8104 , n4884 );
xor ( n8105 , n8103 , n8104 );
xor ( n8106 , n8084 , n8105 );
not ( n8107 , n6583 );
buf ( n8108 , n4885 );
and ( n8109 , n8107 , n8108 );
buf ( n8110 , n4886 );
xor ( n8111 , n8110 , n8108 );
and ( n8112 , n8111 , n6583 );
or ( n8113 , n8109 , n8112 );
not ( n8114 , n6583 );
buf ( n8115 , n4887 );
and ( n8116 , n8114 , n8115 );
buf ( n8117 , n4888 );
xor ( n8118 , n8117 , n8115 );
and ( n8119 , n8118 , n6583 );
or ( n8120 , n8116 , n8119 );
xor ( n8121 , n8113 , n8120 );
buf ( n8122 , n4889 );
xor ( n8123 , n8121 , n8122 );
buf ( n8124 , n4890 );
xor ( n8125 , n8123 , n8124 );
buf ( n8126 , n4891 );
xor ( n8127 , n8125 , n8126 );
xor ( n8128 , n7548 , n8127 );
not ( n8129 , n6583 );
buf ( n8130 , n4892 );
and ( n8131 , n8129 , n8130 );
buf ( n8132 , n4893 );
xor ( n8133 , n8132 , n8130 );
and ( n8134 , n8133 , n6583 );
or ( n8135 , n8131 , n8134 );
xor ( n8136 , n8135 , n7104 );
buf ( n8137 , n4894 );
xor ( n8138 , n8136 , n8137 );
buf ( n8139 , n4895 );
xor ( n8140 , n8138 , n8139 );
buf ( n8141 , n4896 );
xor ( n8142 , n8140 , n8141 );
xor ( n8143 , n8128 , n8142 );
not ( n8144 , n8143 );
buf ( n8145 , n4897 );
not ( n8146 , n6583 );
buf ( n8147 , n4898 );
and ( n8148 , n8146 , n8147 );
buf ( n8149 , n4899 );
xor ( n8150 , n8149 , n8147 );
and ( n8151 , n8150 , n6583 );
or ( n8152 , n8148 , n8151 );
not ( n8153 , n6583 );
buf ( n8154 , n4900 );
and ( n8155 , n8153 , n8154 );
buf ( n8156 , n4901 );
xor ( n8157 , n8156 , n8154 );
and ( n8158 , n8157 , n6583 );
or ( n8159 , n8155 , n8158 );
xor ( n8160 , n8152 , n8159 );
buf ( n8161 , n4902 );
xor ( n8162 , n8160 , n8161 );
buf ( n8163 , n4903 );
xor ( n8164 , n8162 , n8163 );
buf ( n8165 , n4904 );
buf ( n8166 , n8165 );
xor ( n8167 , n8164 , n8166 );
xor ( n8168 , n8145 , n8167 );
not ( n8169 , n6583 );
buf ( n8170 , n4905 );
and ( n8171 , n8169 , n8170 );
buf ( n8172 , n4906 );
xor ( n8173 , n8172 , n8170 );
and ( n8174 , n8173 , n6583 );
or ( n8175 , n8171 , n8174 );
not ( n8176 , n6583 );
buf ( n8177 , n4907 );
and ( n8178 , n8176 , n8177 );
buf ( n8179 , n4908 );
xor ( n8180 , n8179 , n8177 );
and ( n8181 , n8180 , n6583 );
or ( n8182 , n8178 , n8181 );
xor ( n8183 , n8175 , n8182 );
buf ( n8184 , n4909 );
xor ( n8185 , n8183 , n8184 );
buf ( n8186 , n4910 );
xor ( n8187 , n8185 , n8186 );
buf ( n8188 , n4911 );
xor ( n8189 , n8187 , n8188 );
xor ( n8190 , n8168 , n8189 );
and ( n8191 , n8144 , n8190 );
xor ( n8192 , n8106 , n8191 );
buf ( n8193 , n4912 );
buf ( n8194 , n4913 );
or ( n8195 , n8193 , n8194 );
buf ( n8196 , n4914 );
or ( n8197 , n8195 , n8196 );
buf ( n8198 , n4915 );
or ( n8199 , n8197 , n8198 );
buf ( n8200 , n4916 );
or ( n8201 , n8199 , n8200 );
buf ( n8202 , n4917 );
or ( n8203 , n8201 , n8202 );
buf ( n8204 , n4918 );
or ( n8205 , n8203 , n8204 );
xor ( n8206 , n8192 , n8205 );
not ( n8207 , n6583 );
buf ( n8208 , n4919 );
and ( n8209 , n8207 , n8208 );
buf ( n8210 , n4920 );
xor ( n8211 , n8210 , n8208 );
and ( n8212 , n8211 , n6583 );
or ( n8213 , n8209 , n8212 );
not ( n8214 , n6583 );
buf ( n8215 , n4921 );
and ( n8216 , n8214 , n8215 );
buf ( n8217 , n4922 );
xor ( n8218 , n8217 , n8215 );
and ( n8219 , n8218 , n6583 );
or ( n8220 , n8216 , n8219 );
not ( n8221 , n6583 );
buf ( n8222 , n4923 );
and ( n8223 , n8221 , n8222 );
buf ( n8224 , n4924 );
xor ( n8225 , n8224 , n8222 );
and ( n8226 , n8225 , n6583 );
or ( n8227 , n8223 , n8226 );
xor ( n8228 , n8220 , n8227 );
buf ( n8229 , n4925 );
xor ( n8230 , n8228 , n8229 );
buf ( n8231 , n4926 );
xor ( n8232 , n8230 , n8231 );
buf ( n8233 , n4927 );
xor ( n8234 , n8232 , n8233 );
xor ( n8235 , n8213 , n8234 );
not ( n8236 , n6583 );
buf ( n8237 , n4928 );
and ( n8238 , n8236 , n8237 );
buf ( n8239 , n4929 );
xor ( n8240 , n8239 , n8237 );
and ( n8241 , n8240 , n6583 );
or ( n8242 , n8238 , n8241 );
buf ( n8243 , n4930 );
xor ( n8244 , n8242 , n8243 );
buf ( n8245 , n4931 );
xor ( n8246 , n8244 , n8245 );
buf ( n8247 , n4932 );
xor ( n8248 , n8246 , n8247 );
buf ( n8249 , n4933 );
xor ( n8250 , n8248 , n8249 );
xor ( n8251 , n8235 , n8250 );
buf ( n8252 , n4934 );
xor ( n8253 , n8252 , n7428 );
xor ( n8254 , n8253 , n7579 );
not ( n8255 , n8254 );
not ( n8256 , n6583 );
buf ( n8257 , n4935 );
and ( n8258 , n8256 , n8257 );
buf ( n8259 , n4936 );
xor ( n8260 , n8259 , n8257 );
and ( n8261 , n8260 , n6583 );
or ( n8262 , n8258 , n8261 );
buf ( n8263 , n4937 );
xor ( n8264 , n8262 , n8263 );
buf ( n8265 , n4938 );
xor ( n8266 , n8264 , n8265 );
buf ( n8267 , n4939 );
xor ( n8268 , n8266 , n8267 );
buf ( n8269 , n4940 );
xor ( n8270 , n8268 , n8269 );
xor ( n8271 , n6632 , n8270 );
not ( n8272 , n6583 );
buf ( n8273 , n4941 );
and ( n8274 , n8272 , n8273 );
buf ( n8275 , n4942 );
xor ( n8276 , n8275 , n8273 );
and ( n8277 , n8276 , n6583 );
or ( n8278 , n8274 , n8277 );
not ( n8279 , n6583 );
buf ( n8280 , n4943 );
and ( n8281 , n8279 , n8280 );
buf ( n8282 , n4944 );
xor ( n8283 , n8282 , n8280 );
and ( n8284 , n8283 , n6583 );
or ( n8285 , n8281 , n8284 );
xor ( n8286 , n8278 , n8285 );
buf ( n8287 , n4945 );
xor ( n8288 , n8286 , n8287 );
buf ( n8289 , n4946 );
xor ( n8290 , n8288 , n8289 );
buf ( n8291 , n4947 );
xor ( n8292 , n8290 , n8291 );
xor ( n8293 , n8271 , n8292 );
and ( n8294 , n8255 , n8293 );
xor ( n8295 , n8251 , n8294 );
xor ( n8296 , n8206 , n8295 );
not ( n8297 , n6583 );
buf ( n8298 , n4948 );
and ( n8299 , n8297 , n8298 );
buf ( n8300 , n4949 );
xor ( n8301 , n8300 , n8298 );
and ( n8302 , n8301 , n6583 );
or ( n8303 , n8299 , n8302 );
not ( n8304 , n6583 );
buf ( n8305 , n4950 );
and ( n8306 , n8304 , n8305 );
buf ( n8307 , n4951 );
xor ( n8308 , n8307 , n8305 );
and ( n8309 , n8308 , n6583 );
or ( n8310 , n8306 , n8309 );
xor ( n8311 , n8303 , n8310 );
buf ( n8312 , n4952 );
xor ( n8313 , n8311 , n8312 );
buf ( n8314 , n4953 );
xor ( n8315 , n8313 , n8314 );
buf ( n8316 , n4954 );
buf ( n8317 , n8316 );
xor ( n8318 , n8315 , n8317 );
xor ( n8319 , n8091 , n8318 );
not ( n8320 , n6583 );
buf ( n8321 , n4955 );
and ( n8322 , n8320 , n8321 );
buf ( n8323 , n4956 );
xor ( n8324 , n8323 , n8321 );
and ( n8325 , n8324 , n6583 );
or ( n8326 , n8322 , n8325 );
not ( n8327 , n6583 );
buf ( n8328 , n4957 );
and ( n8329 , n8327 , n8328 );
buf ( n8330 , n4958 );
xor ( n8331 , n8330 , n8328 );
and ( n8332 , n8331 , n6583 );
or ( n8333 , n8329 , n8332 );
xor ( n8334 , n8326 , n8333 );
buf ( n8335 , n4959 );
xor ( n8336 , n8334 , n8335 );
buf ( n8337 , n4960 );
xor ( n8338 , n8336 , n8337 );
buf ( n8339 , n4961 );
xor ( n8340 , n8338 , n8339 );
xor ( n8341 , n8319 , n8340 );
not ( n8342 , n6583 );
buf ( n8343 , n4962 );
and ( n8344 , n8342 , n8343 );
buf ( n8345 , n4963 );
xor ( n8346 , n8345 , n8343 );
and ( n8347 , n8346 , n6583 );
or ( n8348 , n8344 , n8347 );
not ( n8349 , n6583 );
buf ( n8350 , n4964 );
and ( n8351 , n8349 , n8350 );
buf ( n8352 , n4965 );
xor ( n8353 , n8352 , n8350 );
and ( n8354 , n8353 , n6583 );
or ( n8355 , n8351 , n8354 );
not ( n8356 , n6583 );
buf ( n8357 , n4966 );
and ( n8358 , n8356 , n8357 );
buf ( n8359 , n4967 );
xor ( n8360 , n8359 , n8357 );
and ( n8361 , n8360 , n6583 );
or ( n8362 , n8358 , n8361 );
xor ( n8363 , n8355 , n8362 );
buf ( n8364 , n4968 );
xor ( n8365 , n8363 , n8364 );
buf ( n8366 , n4969 );
xor ( n8367 , n8365 , n8366 );
buf ( n8368 , n4970 );
xor ( n8369 , n8367 , n8368 );
xor ( n8370 , n8348 , n8369 );
not ( n8371 , n6583 );
buf ( n8372 , n4971 );
and ( n8373 , n8371 , n8372 );
buf ( n8374 , n8373 );
not ( n8375 , n6583 );
buf ( n8376 , n4972 );
and ( n8377 , n8375 , n8376 );
buf ( n8378 , n4973 );
xor ( n8379 , n8378 , n8376 );
and ( n8380 , n8379 , n6583 );
or ( n8381 , n8377 , n8380 );
xor ( n8382 , n8374 , n8381 );
buf ( n8383 , n4974 );
xor ( n8384 , n8382 , n8383 );
buf ( n8385 , n4975 );
xor ( n8386 , n8384 , n8385 );
buf ( n8387 , n4976 );
xor ( n8388 , n8386 , n8387 );
xor ( n8389 , n8370 , n8388 );
not ( n8390 , n8389 );
buf ( n8391 , n4977 );
not ( n8392 , n6583 );
buf ( n8393 , n4978 );
and ( n8394 , n8392 , n8393 );
buf ( n8395 , n4979 );
xor ( n8396 , n8395 , n8393 );
and ( n8397 , n8396 , n6583 );
or ( n8398 , n8394 , n8397 );
not ( n8399 , n6583 );
buf ( n8400 , n4980 );
and ( n8401 , n8399 , n8400 );
buf ( n8402 , n4981 );
xor ( n8403 , n8402 , n8400 );
and ( n8404 , n8403 , n6583 );
or ( n8405 , n8401 , n8404 );
xor ( n8406 , n8398 , n8405 );
buf ( n8407 , n4982 );
xor ( n8408 , n8406 , n8407 );
buf ( n8409 , n4983 );
xor ( n8410 , n8408 , n8409 );
buf ( n8411 , n4984 );
xor ( n8412 , n8410 , n8411 );
xor ( n8413 , n8391 , n8412 );
not ( n8414 , n6583 );
buf ( n8415 , n4985 );
and ( n8416 , n8414 , n8415 );
buf ( n8417 , n4986 );
xor ( n8418 , n8417 , n8415 );
and ( n8419 , n8418 , n6583 );
or ( n8420 , n8416 , n8419 );
buf ( n8421 , n4987 );
xor ( n8422 , n8420 , n8421 );
buf ( n8423 , n4988 );
xor ( n8424 , n8422 , n8423 );
buf ( n8425 , n4989 );
xor ( n8426 , n8424 , n8425 );
buf ( n8427 , n4990 );
xor ( n8428 , n8426 , n8427 );
xor ( n8429 , n8413 , n8428 );
and ( n8430 , n8390 , n8429 );
xor ( n8431 , n8341 , n8430 );
xor ( n8432 , n8296 , n8431 );
not ( n8433 , n6583 );
buf ( n8434 , n4991 );
and ( n8435 , n8433 , n8434 );
buf ( n8436 , n4992 );
xor ( n8437 , n8436 , n8434 );
and ( n8438 , n8437 , n6583 );
or ( n8439 , n8435 , n8438 );
not ( n8440 , n6583 );
buf ( n8441 , n4993 );
and ( n8442 , n8440 , n8441 );
buf ( n8443 , n4994 );
xor ( n8444 , n8443 , n8441 );
and ( n8445 , n8444 , n6583 );
or ( n8446 , n8442 , n8445 );
not ( n8447 , n6583 );
buf ( n8448 , n4995 );
and ( n8449 , n8447 , n8448 );
buf ( n8450 , n4996 );
xor ( n8451 , n8450 , n8448 );
and ( n8452 , n8451 , n6583 );
or ( n8453 , n8449 , n8452 );
xor ( n8454 , n8446 , n8453 );
buf ( n8455 , n4997 );
xor ( n8456 , n8454 , n8455 );
buf ( n8457 , n4998 );
xor ( n8458 , n8456 , n8457 );
buf ( n8459 , n4999 );
xor ( n8460 , n8458 , n8459 );
xor ( n8461 , n8439 , n8460 );
not ( n8462 , n6583 );
buf ( n8463 , n5000 );
and ( n8464 , n8462 , n8463 );
buf ( n8465 , n5001 );
xor ( n8466 , n8465 , n8463 );
and ( n8467 , n8466 , n6583 );
or ( n8468 , n8464 , n8467 );
not ( n8469 , n6583 );
buf ( n8470 , n5002 );
and ( n8471 , n8469 , n8470 );
buf ( n8472 , n5003 );
xor ( n8473 , n8472 , n8470 );
and ( n8474 , n8473 , n6583 );
or ( n8475 , n8471 , n8474 );
xor ( n8476 , n8468 , n8475 );
buf ( n8477 , n5004 );
xor ( n8478 , n8476 , n8477 );
buf ( n8479 , n5005 );
xor ( n8480 , n8478 , n8479 );
buf ( n8481 , n5006 );
xor ( n8482 , n8480 , n8481 );
xor ( n8483 , n8461 , n8482 );
not ( n8484 , n6583 );
buf ( n8485 , n5007 );
and ( n8486 , n8484 , n8485 );
buf ( n8487 , n5008 );
xor ( n8488 , n8487 , n8485 );
and ( n8489 , n8488 , n6583 );
or ( n8490 , n8486 , n8489 );
not ( n8491 , n6583 );
buf ( n8492 , n5009 );
and ( n8493 , n8491 , n8492 );
buf ( n8494 , n5010 );
xor ( n8495 , n8494 , n8492 );
and ( n8496 , n8495 , n6583 );
or ( n8497 , n8493 , n8496 );
buf ( n8498 , n5011 );
xor ( n8499 , n8497 , n8498 );
buf ( n8500 , n5012 );
xor ( n8501 , n8499 , n8500 );
buf ( n8502 , n5013 );
xor ( n8503 , n8501 , n8502 );
buf ( n8504 , n5014 );
xor ( n8505 , n8503 , n8504 );
xor ( n8506 , n8490 , n8505 );
xor ( n8507 , n8506 , n7267 );
not ( n8508 , n8507 );
buf ( n8509 , n5015 );
not ( n8510 , n6583 );
buf ( n8511 , n5016 );
and ( n8512 , n8510 , n8511 );
buf ( n8513 , n5017 );
xor ( n8514 , n8513 , n8511 );
and ( n8515 , n8514 , n6583 );
or ( n8516 , n8512 , n8515 );
not ( n8517 , n6583 );
buf ( n8518 , n5018 );
and ( n8519 , n8517 , n8518 );
buf ( n8520 , n5019 );
xor ( n8521 , n8520 , n8518 );
and ( n8522 , n8521 , n6583 );
or ( n8523 , n8519 , n8522 );
xor ( n8524 , n8516 , n8523 );
buf ( n8525 , n5020 );
xor ( n8526 , n8524 , n8525 );
buf ( n8527 , n5021 );
xor ( n8528 , n8526 , n8527 );
buf ( n8529 , n5022 );
xor ( n8530 , n8528 , n8529 );
xor ( n8531 , n8509 , n8530 );
not ( n8532 , n6583 );
buf ( n8533 , n5023 );
and ( n8534 , n8532 , n8533 );
buf ( n8535 , n5024 );
xor ( n8536 , n8535 , n8533 );
and ( n8537 , n8536 , n6583 );
or ( n8538 , n8534 , n8537 );
not ( n8539 , n6583 );
buf ( n8540 , n5025 );
and ( n8541 , n8539 , n8540 );
buf ( n8542 , n5026 );
xor ( n8543 , n8542 , n8540 );
and ( n8544 , n8543 , n6583 );
or ( n8545 , n8541 , n8544 );
xor ( n8546 , n8538 , n8545 );
buf ( n8547 , n5027 );
xor ( n8548 , n8546 , n8547 );
buf ( n8549 , n5028 );
xor ( n8550 , n8548 , n8549 );
buf ( n8551 , n5029 );
xor ( n8552 , n8550 , n8551 );
xor ( n8553 , n8531 , n8552 );
and ( n8554 , n8508 , n8553 );
xor ( n8555 , n8483 , n8554 );
xor ( n8556 , n8432 , n8555 );
not ( n8557 , n6583 );
buf ( n8558 , n5030 );
and ( n8559 , n8557 , n8558 );
buf ( n8560 , n5031 );
xor ( n8561 , n8560 , n8558 );
and ( n8562 , n8561 , n6583 );
or ( n8563 , n8559 , n8562 );
not ( n8564 , n6583 );
buf ( n8565 , n5032 );
and ( n8566 , n8564 , n8565 );
buf ( n8567 , n5033 );
xor ( n8568 , n8567 , n8565 );
and ( n8569 , n8568 , n6583 );
or ( n8570 , n8566 , n8569 );
not ( n8571 , n6583 );
buf ( n8572 , n5034 );
and ( n8573 , n8571 , n8572 );
buf ( n8574 , n5035 );
xor ( n8575 , n8574 , n8572 );
and ( n8576 , n8575 , n6583 );
or ( n8577 , n8573 , n8576 );
xor ( n8578 , n8570 , n8577 );
buf ( n8579 , n5036 );
xor ( n8580 , n8578 , n8579 );
buf ( n8581 , n5037 );
xor ( n8582 , n8580 , n8581 );
buf ( n8583 , n5038 );
xor ( n8584 , n8582 , n8583 );
xor ( n8585 , n8563 , n8584 );
not ( n8586 , n6583 );
buf ( n8587 , n5039 );
and ( n8588 , n8586 , n8587 );
buf ( n8589 , n5040 );
xor ( n8590 , n8589 , n8587 );
and ( n8591 , n8590 , n6583 );
or ( n8592 , n8588 , n8591 );
not ( n8593 , n6583 );
buf ( n8594 , n5041 );
and ( n8595 , n8593 , n8594 );
buf ( n8596 , n5042 );
xor ( n8597 , n8596 , n8594 );
and ( n8598 , n8597 , n6583 );
or ( n8599 , n8595 , n8598 );
xor ( n8600 , n8592 , n8599 );
buf ( n8601 , n5043 );
xor ( n8602 , n8600 , n8601 );
buf ( n8603 , n5044 );
xor ( n8604 , n8602 , n8603 );
buf ( n8605 , n5045 );
xor ( n8606 , n8604 , n8605 );
xor ( n8607 , n8585 , n8606 );
not ( n8608 , n7997 );
and ( n8609 , n8608 , n8020 );
xor ( n8610 , n8607 , n8609 );
xor ( n8611 , n8556 , n8610 );
xor ( n8612 , n8061 , n8611 );
buf ( n8613 , n5046 );
xor ( n8614 , n8613 , n7555 );
not ( n8615 , n6583 );
buf ( n8616 , n5047 );
and ( n8617 , n8615 , n8616 );
buf ( n8618 , n5048 );
xor ( n8619 , n8618 , n8616 );
and ( n8620 , n8619 , n6583 );
or ( n8621 , n8617 , n8620 );
not ( n8622 , n6583 );
buf ( n8623 , n5049 );
and ( n8624 , n8622 , n8623 );
buf ( n8625 , n5050 );
xor ( n8626 , n8625 , n8623 );
and ( n8627 , n8626 , n6583 );
or ( n8628 , n8624 , n8627 );
xor ( n8629 , n8621 , n8628 );
buf ( n8630 , n5051 );
xor ( n8631 , n8629 , n8630 );
buf ( n8632 , n5052 );
xor ( n8633 , n8631 , n8632 );
buf ( n8634 , n5053 );
xor ( n8635 , n8633 , n8634 );
xor ( n8636 , n8614 , n8635 );
buf ( n8637 , n5054 );
xor ( n8638 , n8637 , n7600 );
not ( n8639 , n6583 );
buf ( n8640 , n5055 );
and ( n8641 , n8639 , n8640 );
buf ( n8642 , n5056 );
xor ( n8643 , n8642 , n8640 );
and ( n8644 , n8643 , n6583 );
or ( n8645 , n8641 , n8644 );
buf ( n8646 , n5057 );
xor ( n8647 , n8645 , n8646 );
buf ( n8648 , n5058 );
xor ( n8649 , n8647 , n8648 );
buf ( n8650 , n5059 );
xor ( n8651 , n8649 , n8650 );
buf ( n8652 , n5060 );
xor ( n8653 , n8651 , n8652 );
xor ( n8654 , n8638 , n8653 );
not ( n8655 , n8654 );
buf ( n8656 , n5061 );
xor ( n8657 , n8656 , n7886 );
xor ( n8658 , n8657 , n7908 );
and ( n8659 , n8655 , n8658 );
xor ( n8660 , n8636 , n8659 );
buf ( n8661 , n5062 );
xor ( n8662 , n8661 , n6963 );
not ( n8663 , n6583 );
buf ( n8664 , n5063 );
and ( n8665 , n8663 , n8664 );
buf ( n8666 , n5064 );
xor ( n8667 , n8666 , n8664 );
and ( n8668 , n8667 , n6583 );
or ( n8669 , n8665 , n8668 );
not ( n8670 , n6583 );
buf ( n8671 , n5065 );
and ( n8672 , n8670 , n8671 );
buf ( n8673 , n5066 );
xor ( n8674 , n8673 , n8671 );
and ( n8675 , n8674 , n6583 );
or ( n8676 , n8672 , n8675 );
xor ( n8677 , n8669 , n8676 );
buf ( n8678 , n5067 );
xor ( n8679 , n8677 , n8678 );
buf ( n8680 , n5068 );
xor ( n8681 , n8679 , n8680 );
buf ( n8682 , n5069 );
xor ( n8683 , n8681 , n8682 );
xor ( n8684 , n8662 , n8683 );
not ( n8685 , n6583 );
buf ( n8686 , n5070 );
and ( n8687 , n8685 , n8686 );
buf ( n8688 , n5071 );
xor ( n8689 , n8688 , n8686 );
and ( n8690 , n8689 , n6583 );
or ( n8691 , n8687 , n8690 );
not ( n8692 , n6583 );
buf ( n8693 , n5072 );
and ( n8694 , n8692 , n8693 );
buf ( n8695 , n5073 );
xor ( n8696 , n8695 , n8693 );
and ( n8697 , n8696 , n6583 );
or ( n8698 , n8694 , n8697 );
xor ( n8699 , n8691 , n8698 );
buf ( n8700 , n5074 );
xor ( n8701 , n8699 , n8700 );
buf ( n8702 , n5075 );
xor ( n8703 , n8701 , n8702 );
buf ( n8704 , n5076 );
xor ( n8705 , n8703 , n8704 );
xor ( n8706 , n7629 , n8705 );
not ( n8707 , n6583 );
buf ( n8708 , n5077 );
and ( n8709 , n8707 , n8708 );
buf ( n8710 , n5078 );
xor ( n8711 , n8710 , n8708 );
and ( n8712 , n8711 , n6583 );
or ( n8713 , n8709 , n8712 );
not ( n8714 , n6583 );
buf ( n8715 , n5079 );
and ( n8716 , n8714 , n8715 );
buf ( n8717 , n5080 );
xor ( n8718 , n8717 , n8715 );
and ( n8719 , n8718 , n6583 );
or ( n8720 , n8716 , n8719 );
xor ( n8721 , n8713 , n8720 );
buf ( n8722 , n5081 );
xor ( n8723 , n8721 , n8722 );
buf ( n8724 , n5082 );
xor ( n8725 , n8723 , n8724 );
buf ( n8726 , n5083 );
xor ( n8727 , n8725 , n8726 );
xor ( n8728 , n8706 , n8727 );
not ( n8729 , n8728 );
buf ( n8730 , n5084 );
xor ( n8731 , n8730 , n8584 );
xor ( n8732 , n8731 , n8606 );
and ( n8733 , n8729 , n8732 );
xor ( n8734 , n8684 , n8733 );
xor ( n8735 , n8660 , n8734 );
buf ( n8736 , n5085 );
not ( n8737 , n6583 );
buf ( n8738 , n5086 );
and ( n8739 , n8737 , n8738 );
buf ( n8740 , n5087 );
xor ( n8741 , n8740 , n8738 );
and ( n8742 , n8741 , n6583 );
or ( n8743 , n8739 , n8742 );
not ( n8744 , n6583 );
buf ( n8745 , n5088 );
and ( n8746 , n8744 , n8745 );
buf ( n8747 , n5089 );
xor ( n8748 , n8747 , n8745 );
and ( n8749 , n8748 , n6583 );
or ( n8750 , n8746 , n8749 );
xor ( n8751 , n8743 , n8750 );
buf ( n8752 , n5090 );
xor ( n8753 , n8751 , n8752 );
buf ( n8754 , n5091 );
xor ( n8755 , n8753 , n8754 );
buf ( n8756 , n5092 );
xor ( n8757 , n8755 , n8756 );
xor ( n8758 , n8736 , n8757 );
buf ( n8759 , n5093 );
xor ( n8760 , n8439 , n8759 );
buf ( n8761 , n5094 );
xor ( n8762 , n8760 , n8761 );
buf ( n8763 , n5095 );
xor ( n8764 , n8762 , n8763 );
buf ( n8765 , n5096 );
xor ( n8766 , n8764 , n8765 );
xor ( n8767 , n8758 , n8766 );
buf ( n8768 , n5097 );
not ( n8769 , n6583 );
buf ( n8770 , n5098 );
and ( n8771 , n8769 , n8770 );
buf ( n8772 , n5099 );
xor ( n8773 , n8772 , n8770 );
and ( n8774 , n8773 , n6583 );
or ( n8775 , n8771 , n8774 );
not ( n8776 , n6583 );
buf ( n8777 , n5100 );
and ( n8778 , n8776 , n8777 );
buf ( n8779 , n5101 );
xor ( n8780 , n8779 , n8777 );
and ( n8781 , n8780 , n6583 );
or ( n8782 , n8778 , n8781 );
xor ( n8783 , n8775 , n8782 );
buf ( n8784 , n5102 );
xor ( n8785 , n8783 , n8784 );
buf ( n8786 , n5103 );
xor ( n8787 , n8785 , n8786 );
buf ( n8788 , n5104 );
xor ( n8789 , n8787 , n8788 );
xor ( n8790 , n8768 , n8789 );
xor ( n8791 , n8790 , n8530 );
not ( n8792 , n8791 );
not ( n8793 , n6583 );
buf ( n8794 , n5105 );
and ( n8795 , n8793 , n8794 );
buf ( n8796 , n5106 );
xor ( n8797 , n8796 , n8794 );
and ( n8798 , n8797 , n6583 );
or ( n8799 , n8795 , n8798 );
buf ( n8800 , n5107 );
xor ( n8801 , n8799 , n8800 );
buf ( n8802 , n5108 );
xor ( n8803 , n8801 , n8802 );
buf ( n8804 , n5109 );
xor ( n8805 , n8803 , n8804 );
buf ( n8806 , n5110 );
xor ( n8807 , n8805 , n8806 );
xor ( n8808 , n6848 , n8807 );
not ( n8809 , n6583 );
buf ( n8810 , n5111 );
and ( n8811 , n8809 , n8810 );
buf ( n8812 , n5112 );
xor ( n8813 , n8812 , n8810 );
and ( n8814 , n8813 , n6583 );
or ( n8815 , n8811 , n8814 );
xor ( n8816 , n8815 , n7347 );
buf ( n8817 , n5113 );
xor ( n8818 , n8816 , n8817 );
buf ( n8819 , n5114 );
xor ( n8820 , n8818 , n8819 );
buf ( n8821 , n5115 );
xor ( n8822 , n8820 , n8821 );
xor ( n8823 , n8808 , n8822 );
and ( n8824 , n8792 , n8823 );
xor ( n8825 , n8767 , n8824 );
xor ( n8826 , n8735 , n8825 );
buf ( n8827 , n5116 );
not ( n8828 , n6583 );
buf ( n8829 , n5117 );
and ( n8830 , n8828 , n8829 );
buf ( n8831 , n5118 );
xor ( n8832 , n8831 , n8829 );
and ( n8833 , n8832 , n6583 );
or ( n8834 , n8830 , n8833 );
xor ( n8835 , n8834 , n6644 );
buf ( n8836 , n5119 );
xor ( n8837 , n8835 , n8836 );
buf ( n8838 , n5120 );
xor ( n8839 , n8837 , n8838 );
buf ( n8840 , n5121 );
xor ( n8841 , n8839 , n8840 );
xor ( n8842 , n8827 , n8841 );
not ( n8843 , n6583 );
buf ( n8844 , n5122 );
and ( n8845 , n8843 , n8844 );
buf ( n8846 , n5123 );
xor ( n8847 , n8846 , n8844 );
and ( n8848 , n8847 , n6583 );
or ( n8849 , n8845 , n8848 );
not ( n8850 , n6583 );
buf ( n8851 , n5124 );
and ( n8852 , n8850 , n8851 );
buf ( n8853 , n5125 );
xor ( n8854 , n8853 , n8851 );
and ( n8855 , n8854 , n6583 );
or ( n8856 , n8852 , n8855 );
xor ( n8857 , n8849 , n8856 );
buf ( n8858 , n5126 );
xor ( n8859 , n8857 , n8858 );
buf ( n8860 , n5127 );
xor ( n8861 , n8859 , n8860 );
buf ( n8862 , n5128 );
xor ( n8863 , n8861 , n8862 );
xor ( n8864 , n8842 , n8863 );
buf ( n8865 , n5129 );
not ( n8866 , n6583 );
buf ( n8867 , n5130 );
and ( n8868 , n8866 , n8867 );
buf ( n8869 , n5131 );
xor ( n8870 , n8869 , n8867 );
and ( n8871 , n8870 , n6583 );
or ( n8872 , n8868 , n8871 );
not ( n8873 , n6583 );
buf ( n8874 , n5132 );
and ( n8875 , n8873 , n8874 );
buf ( n8876 , n5133 );
xor ( n8877 , n8876 , n8874 );
and ( n8878 , n8877 , n6583 );
or ( n8879 , n8875 , n8878 );
xor ( n8880 , n8872 , n8879 );
buf ( n8881 , n5134 );
xor ( n8882 , n8880 , n8881 );
buf ( n8883 , n5135 );
xor ( n8884 , n8882 , n8883 );
buf ( n8885 , n5136 );
xor ( n8886 , n8884 , n8885 );
xor ( n8887 , n8865 , n8886 );
not ( n8888 , n6583 );
buf ( n8889 , n5137 );
and ( n8890 , n8888 , n8889 );
buf ( n8891 , n5138 );
xor ( n8892 , n8891 , n8889 );
and ( n8893 , n8892 , n6583 );
or ( n8894 , n8890 , n8893 );
not ( n8895 , n6583 );
buf ( n8896 , n5139 );
and ( n8897 , n8895 , n8896 );
buf ( n8898 , n5140 );
xor ( n8899 , n8898 , n8896 );
and ( n8900 , n8899 , n6583 );
or ( n8901 , n8897 , n8900 );
xor ( n8902 , n8894 , n8901 );
buf ( n8903 , n5141 );
xor ( n8904 , n8902 , n8903 );
buf ( n8905 , n5142 );
xor ( n8906 , n8904 , n8905 );
buf ( n8907 , n5143 );
xor ( n8908 , n8906 , n8907 );
xor ( n8909 , n8887 , n8908 );
not ( n8910 , n8909 );
buf ( n8911 , n5144 );
not ( n8912 , n6583 );
buf ( n8913 , n5145 );
and ( n8914 , n8912 , n8913 );
buf ( n8915 , n5146 );
xor ( n8916 , n8915 , n8913 );
and ( n8917 , n8916 , n6583 );
or ( n8918 , n8914 , n8917 );
not ( n8919 , n6583 );
buf ( n8920 , n5147 );
and ( n8921 , n8919 , n8920 );
buf ( n8922 , n5148 );
xor ( n8923 , n8922 , n8920 );
and ( n8924 , n8923 , n6583 );
or ( n8925 , n8921 , n8924 );
xor ( n8926 , n8918 , n8925 );
buf ( n8927 , n5149 );
xor ( n8928 , n8926 , n8927 );
buf ( n8929 , n5150 );
xor ( n8930 , n8928 , n8929 );
buf ( n8931 , n5151 );
xor ( n8932 , n8930 , n8931 );
xor ( n8933 , n8911 , n8932 );
not ( n8934 , n6583 );
buf ( n8935 , n5152 );
and ( n8936 , n8934 , n8935 );
buf ( n8937 , n5153 );
xor ( n8938 , n8937 , n8935 );
and ( n8939 , n8938 , n6583 );
or ( n8940 , n8936 , n8939 );
buf ( n8941 , n5154 );
xor ( n8942 , n8940 , n8941 );
buf ( n8943 , n5155 );
xor ( n8944 , n8942 , n8943 );
buf ( n8945 , n5156 );
xor ( n8946 , n8944 , n8945 );
buf ( n8947 , n5157 );
xor ( n8948 , n8946 , n8947 );
xor ( n8949 , n8933 , n8948 );
and ( n8950 , n8910 , n8949 );
xor ( n8951 , n8864 , n8950 );
xor ( n8952 , n8826 , n8951 );
buf ( n8953 , n5158 );
not ( n8954 , n6583 );
buf ( n8955 , n5159 );
and ( n8956 , n8954 , n8955 );
buf ( n8957 , n5160 );
xor ( n8958 , n8957 , n8955 );
and ( n8959 , n8958 , n6583 );
or ( n8960 , n8956 , n8959 );
not ( n8961 , n6583 );
buf ( n8962 , n5161 );
and ( n8963 , n8961 , n8962 );
buf ( n8964 , n5162 );
xor ( n8965 , n8964 , n8962 );
and ( n8966 , n8965 , n6583 );
or ( n8967 , n8963 , n8966 );
xor ( n8968 , n8960 , n8967 );
buf ( n8969 , n5163 );
xor ( n8970 , n8968 , n8969 );
buf ( n8971 , n5164 );
xor ( n8972 , n8970 , n8971 );
buf ( n8973 , n5165 );
xor ( n8974 , n8972 , n8973 );
xor ( n8975 , n8953 , n8974 );
xor ( n8976 , n8975 , n7216 );
buf ( n8977 , n5166 );
not ( n8978 , n6583 );
buf ( n8979 , n5167 );
and ( n8980 , n8978 , n8979 );
buf ( n8981 , n5168 );
xor ( n8982 , n8981 , n8979 );
and ( n8983 , n8982 , n6583 );
or ( n8984 , n8980 , n8983 );
buf ( n8985 , n5169 );
xor ( n8986 , n8984 , n8985 );
buf ( n8987 , n5170 );
xor ( n8988 , n8986 , n8987 );
buf ( n8989 , n5171 );
xor ( n8990 , n8988 , n8989 );
buf ( n8991 , n5172 );
xor ( n8992 , n8990 , n8991 );
xor ( n8993 , n8977 , n8992 );
xor ( n8994 , n8993 , n8167 );
not ( n8995 , n8994 );
buf ( n8996 , n5173 );
xor ( n8997 , n8996 , n6636 );
not ( n8998 , n6583 );
buf ( n8999 , n5174 );
and ( n9000 , n8998 , n8999 );
buf ( n9001 , n5175 );
xor ( n9002 , n9001 , n8999 );
and ( n9003 , n9002 , n6583 );
or ( n9004 , n9000 , n9003 );
not ( n9005 , n6583 );
buf ( n9006 , n5176 );
and ( n9007 , n9005 , n9006 );
buf ( n9008 , n5177 );
xor ( n9009 , n9008 , n9006 );
and ( n9010 , n9009 , n6583 );
or ( n9011 , n9007 , n9010 );
xor ( n9012 , n9004 , n9011 );
buf ( n9013 , n5178 );
xor ( n9014 , n9012 , n9013 );
buf ( n9015 , n5179 );
xor ( n9016 , n9014 , n9015 );
buf ( n9017 , n5180 );
xor ( n9018 , n9016 , n9017 );
xor ( n9019 , n8997 , n9018 );
and ( n9020 , n8995 , n9019 );
xor ( n9021 , n8976 , n9020 );
xor ( n9022 , n8952 , n9021 );
xor ( n9023 , n8612 , n9022 );
not ( n9024 , n9023 );
buf ( n9025 , n5181 );
not ( n9026 , n6583 );
buf ( n9027 , n5182 );
and ( n9028 , n9026 , n9027 );
buf ( n9029 , n5183 );
xor ( n9030 , n9029 , n9027 );
and ( n9031 , n9030 , n6583 );
or ( n9032 , n9028 , n9031 );
not ( n9033 , n6583 );
buf ( n9034 , n5184 );
and ( n9035 , n9033 , n9034 );
buf ( n9036 , n5185 );
xor ( n9037 , n9036 , n9034 );
and ( n9038 , n9037 , n6583 );
or ( n9039 , n9035 , n9038 );
xor ( n9040 , n9032 , n9039 );
buf ( n9041 , n5186 );
xor ( n9042 , n9040 , n9041 );
buf ( n9043 , n5187 );
xor ( n9044 , n9042 , n9043 );
buf ( n9045 , n5188 );
xor ( n9046 , n9044 , n9045 );
xor ( n9047 , n9025 , n9046 );
xor ( n9048 , n9047 , n8974 );
not ( n9049 , n6583 );
buf ( n9050 , n5189 );
and ( n9051 , n9049 , n9050 );
buf ( n9052 , n5190 );
xor ( n9053 , n9052 , n9050 );
and ( n9054 , n9053 , n6583 );
or ( n9055 , n9051 , n9054 );
not ( n9056 , n6583 );
buf ( n9057 , n5191 );
and ( n9058 , n9056 , n9057 );
buf ( n9059 , n5192 );
xor ( n9060 , n9059 , n9057 );
and ( n9061 , n9060 , n6583 );
or ( n9062 , n9058 , n9061 );
xor ( n9063 , n9055 , n9062 );
buf ( n9064 , n5193 );
xor ( n9065 , n9063 , n9064 );
buf ( n9066 , n5194 );
xor ( n9067 , n9065 , n9066 );
buf ( n9068 , n5195 );
xor ( n9069 , n9067 , n9068 );
xor ( n9070 , n8905 , n9069 );
not ( n9071 , n6583 );
buf ( n9072 , n5196 );
and ( n9073 , n9071 , n9072 );
buf ( n9074 , n5197 );
xor ( n9075 , n9074 , n9072 );
and ( n9076 , n9075 , n6583 );
or ( n9077 , n9073 , n9076 );
buf ( n9078 , n5198 );
xor ( n9079 , n9077 , n9078 );
buf ( n9080 , n5199 );
xor ( n9081 , n9079 , n9080 );
buf ( n9082 , n5200 );
xor ( n9083 , n9081 , n9082 );
buf ( n9084 , n5201 );
xor ( n9085 , n9083 , n9084 );
xor ( n9086 , n9070 , n9085 );
not ( n9087 , n9086 );
buf ( n9088 , n5202 );
not ( n9089 , n6583 );
buf ( n9090 , n5203 );
and ( n9091 , n9089 , n9090 );
buf ( n9092 , n5204 );
xor ( n9093 , n9092 , n9090 );
and ( n9094 , n9093 , n6583 );
or ( n9095 , n9091 , n9094 );
not ( n9096 , n6583 );
buf ( n9097 , n5205 );
and ( n9098 , n9096 , n9097 );
buf ( n9099 , n5206 );
xor ( n9100 , n9099 , n9097 );
and ( n9101 , n9100 , n6583 );
or ( n9102 , n9098 , n9101 );
xor ( n9103 , n9095 , n9102 );
buf ( n9104 , n5207 );
xor ( n9105 , n9103 , n9104 );
buf ( n9106 , n5208 );
xor ( n9107 , n9105 , n9106 );
buf ( n9108 , n5209 );
xor ( n9109 , n9107 , n9108 );
xor ( n9110 , n9088 , n9109 );
xor ( n9111 , n9110 , n8841 );
and ( n9112 , n9087 , n9111 );
xor ( n9113 , n9048 , n9112 );
xor ( n9114 , n6812 , n7073 );
xor ( n9115 , n9114 , n7095 );
not ( n9116 , n9048 );
and ( n9117 , n9116 , n9086 );
xor ( n9118 , n9115 , n9117 );
buf ( n9119 , n5210 );
not ( n9120 , n6583 );
buf ( n9121 , n5211 );
and ( n9122 , n9120 , n9121 );
buf ( n9123 , n5212 );
xor ( n9124 , n9123 , n9121 );
and ( n9125 , n9124 , n6583 );
or ( n9126 , n9122 , n9125 );
not ( n9127 , n6583 );
buf ( n9128 , n5213 );
and ( n9129 , n9127 , n9128 );
buf ( n9130 , n5214 );
xor ( n9131 , n9130 , n9128 );
and ( n9132 , n9131 , n6583 );
or ( n9133 , n9129 , n9132 );
xor ( n9134 , n9126 , n9133 );
buf ( n9135 , n5215 );
xor ( n9136 , n9134 , n9135 );
buf ( n9137 , n5216 );
xor ( n9138 , n9136 , n9137 );
buf ( n9139 , n5217 );
xor ( n9140 , n9138 , n9139 );
xor ( n9141 , n9119 , n9140 );
not ( n9142 , n6583 );
buf ( n9143 , n5218 );
and ( n9144 , n9142 , n9143 );
buf ( n9145 , n5219 );
xor ( n9146 , n9145 , n9143 );
and ( n9147 , n9146 , n6583 );
or ( n9148 , n9144 , n9147 );
not ( n9149 , n6583 );
buf ( n9150 , n5220 );
and ( n9151 , n9149 , n9150 );
buf ( n9152 , n5221 );
xor ( n9153 , n9152 , n9150 );
and ( n9154 , n9153 , n6583 );
or ( n9155 , n9151 , n9154 );
xor ( n9156 , n9148 , n9155 );
buf ( n9157 , n5222 );
xor ( n9158 , n9156 , n9157 );
xor ( n9159 , n9158 , n7911 );
buf ( n9160 , n5223 );
xor ( n9161 , n9159 , n9160 );
xor ( n9162 , n9141 , n9161 );
buf ( n9163 , n5224 );
not ( n9164 , n6583 );
buf ( n9165 , n5225 );
and ( n9166 , n9164 , n9165 );
buf ( n9167 , n5226 );
xor ( n9168 , n9167 , n9165 );
and ( n9169 , n9168 , n6583 );
or ( n9170 , n9166 , n9169 );
buf ( n9171 , n5227 );
xor ( n9172 , n9170 , n9171 );
buf ( n9173 , n5228 );
xor ( n9174 , n9172 , n9173 );
buf ( n9175 , n5229 );
xor ( n9176 , n9174 , n9175 );
buf ( n9177 , n5230 );
xor ( n9178 , n9176 , n9177 );
xor ( n9179 , n9163 , n9178 );
not ( n9180 , n6583 );
buf ( n9181 , n5231 );
and ( n9182 , n9180 , n9181 );
buf ( n9183 , n5232 );
xor ( n9184 , n9183 , n9181 );
and ( n9185 , n9184 , n6583 );
or ( n9186 , n9182 , n9185 );
not ( n9187 , n6583 );
buf ( n9188 , n5233 );
and ( n9189 , n9187 , n9188 );
buf ( n9190 , n5234 );
xor ( n9191 , n9190 , n9188 );
and ( n9192 , n9191 , n6583 );
or ( n9193 , n9189 , n9192 );
xor ( n9194 , n9186 , n9193 );
buf ( n9195 , n5235 );
xor ( n9196 , n9194 , n9195 );
buf ( n9197 , n5236 );
xor ( n9198 , n9196 , n9197 );
buf ( n9199 , n5237 );
xor ( n9200 , n9198 , n9199 );
xor ( n9201 , n9179 , n9200 );
not ( n9202 , n9201 );
buf ( n9203 , n5238 );
xor ( n9204 , n9203 , n7216 );
xor ( n9205 , n9204 , n7238 );
and ( n9206 , n9202 , n9205 );
xor ( n9207 , n9162 , n9206 );
xor ( n9208 , n9118 , n9207 );
not ( n9209 , n6583 );
buf ( n9210 , n5239 );
and ( n9211 , n9209 , n9210 );
buf ( n9212 , n5240 );
xor ( n9213 , n9212 , n9210 );
and ( n9214 , n9213 , n6583 );
or ( n9215 , n9211 , n9214 );
not ( n9216 , n6583 );
buf ( n9217 , n5241 );
and ( n9218 , n9216 , n9217 );
buf ( n9219 , n5242 );
xor ( n9220 , n9219 , n9217 );
and ( n9221 , n9220 , n6583 );
or ( n9222 , n9218 , n9221 );
xor ( n9223 , n9215 , n9222 );
buf ( n9224 , n5243 );
xor ( n9225 , n9223 , n9224 );
buf ( n9226 , n5244 );
xor ( n9227 , n9225 , n9226 );
buf ( n9228 , n5245 );
xor ( n9229 , n9227 , n9228 );
xor ( n9230 , n8333 , n9229 );
not ( n9231 , n6583 );
buf ( n9232 , n5246 );
and ( n9233 , n9231 , n9232 );
buf ( n9234 , n5247 );
xor ( n9235 , n9234 , n9232 );
and ( n9236 , n9235 , n6583 );
or ( n9237 , n9233 , n9236 );
xor ( n9238 , n6926 , n9237 );
buf ( n9239 , n5248 );
xor ( n9240 , n9238 , n9239 );
buf ( n9241 , n5249 );
xor ( n9242 , n9240 , n9241 );
buf ( n9243 , n5250 );
xor ( n9244 , n9242 , n9243 );
xor ( n9245 , n9230 , n9244 );
buf ( n9246 , n5251 );
xor ( n9247 , n9246 , n7390 );
not ( n9248 , n6583 );
buf ( n9249 , n5252 );
and ( n9250 , n9248 , n9249 );
buf ( n9251 , n5253 );
xor ( n9252 , n9251 , n9249 );
and ( n9253 , n9252 , n6583 );
or ( n9254 , n9250 , n9253 );
buf ( n9255 , n5254 );
xor ( n9256 , n9254 , n9255 );
buf ( n9257 , n5255 );
xor ( n9258 , n9256 , n9257 );
buf ( n9259 , n5256 );
xor ( n9260 , n9258 , n9259 );
buf ( n9261 , n5257 );
xor ( n9262 , n9260 , n9261 );
xor ( n9263 , n9247 , n9262 );
not ( n9264 , n9263 );
not ( n9265 , n6583 );
buf ( n9266 , n5258 );
and ( n9267 , n9265 , n9266 );
buf ( n9268 , n5259 );
xor ( n9269 , n9268 , n9266 );
and ( n9270 , n9269 , n6583 );
or ( n9271 , n9267 , n9270 );
not ( n9272 , n6583 );
buf ( n9273 , n5260 );
and ( n9274 , n9272 , n9273 );
buf ( n9275 , n5261 );
xor ( n9276 , n9275 , n9273 );
and ( n9277 , n9276 , n6583 );
or ( n9278 , n9274 , n9277 );
xor ( n9279 , n9271 , n9278 );
buf ( n9280 , n5262 );
xor ( n9281 , n9279 , n9280 );
buf ( n9282 , n5263 );
xor ( n9283 , n9281 , n9282 );
buf ( n9284 , n5264 );
xor ( n9285 , n9283 , n9284 );
xor ( n9286 , n6960 , n9285 );
not ( n9287 , n6583 );
buf ( n9288 , n5265 );
and ( n9289 , n9287 , n9288 );
buf ( n9290 , n5266 );
xor ( n9291 , n9290 , n9288 );
and ( n9292 , n9291 , n6583 );
or ( n9293 , n9289 , n9292 );
not ( n9294 , n6583 );
buf ( n9295 , n5267 );
and ( n9296 , n9294 , n9295 );
buf ( n9297 , n5268 );
xor ( n9298 , n9297 , n9295 );
and ( n9299 , n9298 , n6583 );
or ( n9300 , n9296 , n9299 );
xor ( n9301 , n9293 , n9300 );
buf ( n9302 , n5269 );
xor ( n9303 , n9301 , n9302 );
buf ( n9304 , n5270 );
xor ( n9305 , n9303 , n9304 );
buf ( n9306 , n5271 );
xor ( n9307 , n9305 , n9306 );
xor ( n9308 , n9286 , n9307 );
and ( n9309 , n9264 , n9308 );
xor ( n9310 , n9245 , n9309 );
xor ( n9311 , n9208 , n9310 );
not ( n9312 , n6583 );
buf ( n9313 , n5272 );
and ( n9314 , n9312 , n9313 );
buf ( n9315 , n5273 );
xor ( n9316 , n9315 , n9313 );
and ( n9317 , n9316 , n6583 );
or ( n9318 , n9314 , n9317 );
xor ( n9319 , n9318 , n7189 );
not ( n9320 , n6583 );
buf ( n9321 , n5274 );
and ( n9322 , n9320 , n9321 );
buf ( n9323 , n5275 );
xor ( n9324 , n9323 , n9321 );
and ( n9325 , n9324 , n6583 );
or ( n9326 , n9322 , n9325 );
not ( n9327 , n6583 );
buf ( n9328 , n5276 );
and ( n9329 , n9327 , n9328 );
buf ( n9330 , n5277 );
xor ( n9331 , n9330 , n9328 );
and ( n9332 , n9331 , n6583 );
or ( n9333 , n9329 , n9332 );
xor ( n9334 , n9326 , n9333 );
buf ( n9335 , n5278 );
xor ( n9336 , n9334 , n9335 );
buf ( n9337 , n5279 );
xor ( n9338 , n9336 , n9337 );
buf ( n9339 , n5280 );
xor ( n9340 , n9338 , n9339 );
xor ( n9341 , n9319 , n9340 );
not ( n9342 , n6583 );
buf ( n9343 , n5281 );
and ( n9344 , n9342 , n9343 );
buf ( n9345 , n5282 );
xor ( n9346 , n9345 , n9343 );
and ( n9347 , n9346 , n6583 );
or ( n9348 , n9344 , n9347 );
not ( n9349 , n6583 );
buf ( n9350 , n5283 );
and ( n9351 , n9349 , n9350 );
buf ( n9352 , n5284 );
xor ( n9353 , n9352 , n9350 );
and ( n9354 , n9353 , n6583 );
or ( n9355 , n9351 , n9354 );
xor ( n9356 , n9348 , n9355 );
buf ( n9357 , n5285 );
xor ( n9358 , n9356 , n9357 );
buf ( n9359 , n5286 );
xor ( n9360 , n9358 , n9359 );
buf ( n9361 , n5287 );
xor ( n9362 , n9360 , n9361 );
xor ( n9363 , n8364 , n9362 );
not ( n9364 , n6583 );
buf ( n9365 , n5288 );
and ( n9366 , n9364 , n9365 );
buf ( n9367 , n5289 );
xor ( n9368 , n9367 , n9365 );
and ( n9369 , n9368 , n6583 );
or ( n9370 , n9366 , n9369 );
not ( n9371 , n6583 );
buf ( n9372 , n5290 );
and ( n9373 , n9371 , n9372 );
buf ( n9374 , n5291 );
xor ( n9375 , n9374 , n9372 );
and ( n9376 , n9375 , n6583 );
or ( n9377 , n9373 , n9376 );
xor ( n9378 , n9370 , n9377 );
buf ( n9379 , n5292 );
xor ( n9380 , n9378 , n9379 );
buf ( n9381 , n5293 );
xor ( n9382 , n9380 , n9381 );
buf ( n9383 , n5294 );
xor ( n9384 , n9382 , n9383 );
xor ( n9385 , n9363 , n9384 );
not ( n9386 , n9385 );
not ( n9387 , n6583 );
buf ( n9388 , n5295 );
and ( n9389 , n9387 , n9388 );
buf ( n9390 , n5296 );
xor ( n9391 , n9390 , n9388 );
and ( n9392 , n9391 , n6583 );
or ( n9393 , n9389 , n9392 );
not ( n9394 , n6583 );
buf ( n9395 , n5297 );
and ( n9396 , n9394 , n9395 );
buf ( n9397 , n5298 );
xor ( n9398 , n9397 , n9395 );
and ( n9399 , n9398 , n6583 );
or ( n9400 , n9396 , n9399 );
xor ( n9401 , n9393 , n9400 );
xor ( n9402 , n9401 , n8827 );
buf ( n9403 , n5299 );
xor ( n9404 , n9402 , n9403 );
buf ( n9405 , n5300 );
xor ( n9406 , n9404 , n9405 );
xor ( n9407 , n8549 , n9406 );
not ( n9408 , n6583 );
buf ( n9409 , n5301 );
and ( n9410 , n9408 , n9409 );
buf ( n9411 , n5302 );
xor ( n9412 , n9411 , n9409 );
and ( n9413 , n9412 , n6583 );
or ( n9414 , n9410 , n9413 );
not ( n9415 , n6583 );
buf ( n9416 , n5303 );
and ( n9417 , n9415 , n9416 );
buf ( n9418 , n5304 );
xor ( n9419 , n9418 , n9416 );
and ( n9420 , n9419 , n6583 );
or ( n9421 , n9417 , n9420 );
xor ( n9422 , n9414 , n9421 );
buf ( n9423 , n5305 );
xor ( n9424 , n9422 , n9423 );
buf ( n9425 , n5306 );
xor ( n9426 , n9424 , n9425 );
buf ( n9427 , n5307 );
xor ( n9428 , n9426 , n9427 );
xor ( n9429 , n9407 , n9428 );
and ( n9430 , n9386 , n9429 );
xor ( n9431 , n9341 , n9430 );
xor ( n9432 , n9311 , n9431 );
not ( n9433 , n6583 );
buf ( n9434 , n5308 );
and ( n9435 , n9433 , n9434 );
buf ( n9436 , n5309 );
xor ( n9437 , n9436 , n9434 );
and ( n9438 , n9437 , n6583 );
or ( n9439 , n9435 , n9438 );
xor ( n9440 , n9439 , n7804 );
not ( n9441 , n6583 );
buf ( n9442 , n5310 );
and ( n9443 , n9441 , n9442 );
buf ( n9444 , n5311 );
xor ( n9445 , n9444 , n9442 );
and ( n9446 , n9445 , n6583 );
or ( n9447 , n9443 , n9446 );
buf ( n9448 , n5312 );
xor ( n9449 , n9447 , n9448 );
buf ( n9450 , n5313 );
xor ( n9451 , n9449 , n9450 );
buf ( n9452 , n5314 );
xor ( n9453 , n9451 , n9452 );
buf ( n9454 , n5315 );
xor ( n9455 , n9453 , n9454 );
xor ( n9456 , n9440 , n9455 );
buf ( n9457 , n5316 );
not ( n9458 , n6583 );
buf ( n9459 , n5317 );
and ( n9460 , n9458 , n9459 );
buf ( n9461 , n5318 );
xor ( n9462 , n9461 , n9459 );
and ( n9463 , n9462 , n6583 );
or ( n9464 , n9460 , n9463 );
not ( n9465 , n6583 );
buf ( n9466 , n5319 );
and ( n9467 , n9465 , n9466 );
buf ( n9468 , n5320 );
xor ( n9469 , n9468 , n9466 );
and ( n9470 , n9469 , n6583 );
or ( n9471 , n9467 , n9470 );
xor ( n9472 , n9464 , n9471 );
buf ( n9473 , n5321 );
xor ( n9474 , n9472 , n9473 );
buf ( n9475 , n5322 );
xor ( n9476 , n9474 , n9475 );
buf ( n9477 , n5323 );
xor ( n9478 , n9476 , n9477 );
xor ( n9479 , n9457 , n9478 );
not ( n9480 , n6583 );
buf ( n9481 , n5324 );
and ( n9482 , n9480 , n9481 );
buf ( n9483 , n5325 );
xor ( n9484 , n9483 , n9481 );
and ( n9485 , n9484 , n6583 );
or ( n9486 , n9482 , n9485 );
xor ( n9487 , n9486 , n8490 );
buf ( n9488 , n5326 );
xor ( n9489 , n9487 , n9488 );
buf ( n9490 , n5327 );
xor ( n9491 , n9489 , n9490 );
buf ( n9492 , n5328 );
xor ( n9493 , n9491 , n9492 );
xor ( n9494 , n9479 , n9493 );
not ( n9495 , n9494 );
buf ( n9496 , n5329 );
not ( n9497 , n6583 );
buf ( n9498 , n5330 );
and ( n9499 , n9497 , n9498 );
buf ( n9500 , n5331 );
xor ( n9501 , n9500 , n9498 );
and ( n9502 , n9501 , n6583 );
or ( n9503 , n9499 , n9502 );
buf ( n9504 , n5332 );
xor ( n9505 , n9503 , n9504 );
buf ( n9506 , n5333 );
xor ( n9507 , n9505 , n9506 );
buf ( n9508 , n5334 );
xor ( n9509 , n9507 , n9508 );
buf ( n9510 , n5335 );
xor ( n9511 , n9509 , n9510 );
xor ( n9512 , n9496 , n9511 );
not ( n9513 , n6583 );
buf ( n9514 , n5336 );
and ( n9515 , n9513 , n9514 );
buf ( n9516 , n5337 );
xor ( n9517 , n9516 , n9514 );
and ( n9518 , n9517 , n6583 );
or ( n9519 , n9515 , n9518 );
not ( n9520 , n6583 );
buf ( n9521 , n5338 );
and ( n9522 , n9520 , n9521 );
buf ( n9523 , n5339 );
xor ( n9524 , n9523 , n9521 );
and ( n9525 , n9524 , n6583 );
or ( n9526 , n9522 , n9525 );
xor ( n9527 , n9519 , n9526 );
buf ( n9528 , n5340 );
xor ( n9529 , n9527 , n9528 );
buf ( n9530 , n5341 );
xor ( n9531 , n9529 , n9530 );
buf ( n9532 , n5342 );
xor ( n9533 , n9531 , n9532 );
xor ( n9534 , n9512 , n9533 );
and ( n9535 , n9495 , n9534 );
xor ( n9536 , n9456 , n9535 );
xor ( n9537 , n9432 , n9536 );
xor ( n9538 , n9113 , n9537 );
buf ( n9539 , n5343 );
not ( n9540 , n6583 );
buf ( n9541 , n5344 );
and ( n9542 , n9540 , n9541 );
buf ( n9543 , n5345 );
xor ( n9544 , n9543 , n9541 );
and ( n9545 , n9544 , n6583 );
or ( n9546 , n9542 , n9545 );
not ( n9547 , n6583 );
buf ( n9548 , n5346 );
and ( n9549 , n9547 , n9548 );
buf ( n9550 , n5347 );
xor ( n9551 , n9550 , n9548 );
and ( n9552 , n9551 , n6583 );
or ( n9553 , n9549 , n9552 );
xor ( n9554 , n9546 , n9553 );
buf ( n9555 , n5348 );
xor ( n9556 , n9554 , n9555 );
buf ( n9557 , n5349 );
xor ( n9558 , n9556 , n9557 );
buf ( n9559 , n5350 );
xor ( n9560 , n9558 , n9559 );
xor ( n9561 , n9539 , n9560 );
xor ( n9562 , n9561 , n8807 );
not ( n9563 , n6583 );
buf ( n9564 , n5351 );
and ( n9565 , n9563 , n9564 );
buf ( n9566 , n5352 );
xor ( n9567 , n9566 , n9564 );
and ( n9568 , n9567 , n6583 );
or ( n9569 , n9565 , n9568 );
not ( n9570 , n6583 );
buf ( n9571 , n5353 );
and ( n9572 , n9570 , n9571 );
buf ( n9573 , n5354 );
xor ( n9574 , n9573 , n9571 );
and ( n9575 , n9574 , n6583 );
or ( n9576 , n9572 , n9575 );
xor ( n9577 , n9569 , n9576 );
buf ( n9578 , n5355 );
xor ( n9579 , n9577 , n9578 );
buf ( n9580 , n5356 );
xor ( n9581 , n9579 , n9580 );
buf ( n9582 , n5357 );
xor ( n9583 , n9581 , n9582 );
xor ( n9584 , n6658 , n9583 );
not ( n9585 , n6583 );
buf ( n9586 , n5358 );
and ( n9587 , n9585 , n9586 );
buf ( n9588 , n5359 );
xor ( n9589 , n9588 , n9586 );
and ( n9590 , n9589 , n6583 );
or ( n9591 , n9587 , n9590 );
xor ( n9592 , n9591 , n7722 );
buf ( n9593 , n5360 );
xor ( n9594 , n9592 , n9593 );
buf ( n9595 , n5361 );
xor ( n9596 , n9594 , n9595 );
buf ( n9597 , n5362 );
xor ( n9598 , n9596 , n9597 );
xor ( n9599 , n9584 , n9598 );
not ( n9600 , n9599 );
not ( n9601 , n6583 );
buf ( n9602 , n5363 );
and ( n9603 , n9601 , n9602 );
buf ( n9604 , n5364 );
xor ( n9605 , n9604 , n9602 );
and ( n9606 , n9605 , n6583 );
or ( n9607 , n9603 , n9606 );
buf ( n9608 , n5365 );
xor ( n9609 , n9607 , n9608 );
buf ( n9610 , n5366 );
xor ( n9611 , n9609 , n9610 );
buf ( n9612 , n5367 );
xor ( n9613 , n9611 , n9612 );
buf ( n9614 , n5368 );
xor ( n9615 , n9613 , n9614 );
xor ( n9616 , n7502 , n9615 );
xor ( n9617 , n9616 , n8584 );
and ( n9618 , n9600 , n9617 );
xor ( n9619 , n9562 , n9618 );
not ( n9620 , n6583 );
buf ( n9621 , n5369 );
and ( n9622 , n9620 , n9621 );
buf ( n9623 , n5370 );
xor ( n9624 , n9623 , n9621 );
and ( n9625 , n9624 , n6583 );
or ( n9626 , n9622 , n9625 );
not ( n9627 , n6583 );
buf ( n9628 , n5371 );
and ( n9629 , n9627 , n9628 );
buf ( n9630 , n5372 );
xor ( n9631 , n9630 , n9628 );
and ( n9632 , n9631 , n6583 );
or ( n9633 , n9629 , n9632 );
xor ( n9634 , n9626 , n9633 );
buf ( n9635 , n5373 );
xor ( n9636 , n9634 , n9635 );
xor ( n9637 , n9636 , n8977 );
buf ( n9638 , n5374 );
xor ( n9639 , n9637 , n9638 );
xor ( n9640 , n8055 , n9639 );
not ( n9641 , n6583 );
buf ( n9642 , n5375 );
and ( n9643 , n9641 , n9642 );
buf ( n9644 , n5376 );
xor ( n9645 , n9644 , n9642 );
and ( n9646 , n9645 , n6583 );
or ( n9647 , n9643 , n9646 );
not ( n9648 , n6583 );
buf ( n9649 , n5377 );
and ( n9650 , n9648 , n9649 );
buf ( n9651 , n5378 );
xor ( n9652 , n9651 , n9649 );
and ( n9653 , n9652 , n6583 );
or ( n9654 , n9650 , n9653 );
xor ( n9655 , n9647 , n9654 );
xor ( n9656 , n9655 , n8145 );
buf ( n9657 , n5379 );
xor ( n9658 , n9656 , n9657 );
buf ( n9659 , n5380 );
xor ( n9660 , n9658 , n9659 );
xor ( n9661 , n9640 , n9660 );
buf ( n9662 , n5381 );
xor ( n9663 , n9662 , n7051 );
xor ( n9664 , n9663 , n6987 );
not ( n9665 , n9664 );
not ( n9666 , n6583 );
buf ( n9667 , n5382 );
and ( n9668 , n9666 , n9667 );
buf ( n9669 , n5383 );
xor ( n9670 , n9669 , n9667 );
and ( n9671 , n9670 , n6583 );
or ( n9672 , n9668 , n9671 );
xor ( n9673 , n9672 , n8412 );
xor ( n9674 , n9673 , n8428 );
and ( n9675 , n9665 , n9674 );
xor ( n9676 , n9661 , n9675 );
xor ( n9677 , n9619 , n9676 );
buf ( n9678 , n5384 );
not ( n9679 , n6583 );
buf ( n9680 , n5385 );
and ( n9681 , n9679 , n9680 );
buf ( n9682 , n5386 );
xor ( n9683 , n9682 , n9680 );
and ( n9684 , n9683 , n6583 );
or ( n9685 , n9681 , n9684 );
not ( n9686 , n6583 );
buf ( n9687 , n5387 );
and ( n9688 , n9686 , n9687 );
buf ( n9689 , n5388 );
xor ( n9690 , n9689 , n9687 );
and ( n9691 , n9690 , n6583 );
or ( n9692 , n9688 , n9691 );
xor ( n9693 , n9685 , n9692 );
buf ( n9694 , n5389 );
xor ( n9695 , n9693 , n9694 );
buf ( n9696 , n5390 );
xor ( n9697 , n9695 , n9696 );
buf ( n9698 , n5391 );
xor ( n9699 , n9697 , n9698 );
xor ( n9700 , n9678 , n9699 );
xor ( n9701 , n9700 , n9362 );
buf ( n9702 , n5392 );
not ( n9703 , n6583 );
buf ( n9704 , n5393 );
and ( n9705 , n9703 , n9704 );
buf ( n9706 , n5394 );
xor ( n9707 , n9706 , n9704 );
and ( n9708 , n9707 , n6583 );
or ( n9709 , n9705 , n9708 );
buf ( n9710 , n5395 );
xor ( n9711 , n9709 , n9710 );
xor ( n9712 , n9711 , n7865 );
buf ( n9713 , n5396 );
xor ( n9714 , n9712 , n9713 );
xor ( n9715 , n9714 , n8656 );
xor ( n9716 , n9702 , n9715 );
xor ( n9717 , n9716 , n8886 );
not ( n9718 , n9717 );
not ( n9719 , n6583 );
buf ( n9720 , n5397 );
and ( n9721 , n9719 , n9720 );
buf ( n9722 , n5398 );
xor ( n9723 , n9722 , n9720 );
and ( n9724 , n9723 , n6583 );
or ( n9725 , n9721 , n9724 );
not ( n9726 , n6583 );
buf ( n9727 , n5399 );
and ( n9728 , n9726 , n9727 );
buf ( n9729 , n5400 );
xor ( n9730 , n9729 , n9727 );
and ( n9731 , n9730 , n6583 );
or ( n9732 , n9728 , n9731 );
xor ( n9733 , n9725 , n9732 );
buf ( n9734 , n5401 );
xor ( n9735 , n9733 , n9734 );
buf ( n9736 , n5402 );
xor ( n9737 , n9735 , n9736 );
buf ( n9738 , n5403 );
xor ( n9739 , n9737 , n9738 );
xor ( n9740 , n8570 , n9739 );
not ( n9741 , n6583 );
buf ( n9742 , n5404 );
and ( n9743 , n9741 , n9742 );
buf ( n9744 , n5405 );
xor ( n9745 , n9744 , n9742 );
and ( n9746 , n9745 , n6583 );
or ( n9747 , n9743 , n9746 );
not ( n9748 , n6583 );
buf ( n9749 , n5406 );
and ( n9750 , n9748 , n9749 );
buf ( n9751 , n5407 );
xor ( n9752 , n9751 , n9749 );
and ( n9753 , n9752 , n6583 );
or ( n9754 , n9750 , n9753 );
xor ( n9755 , n9747 , n9754 );
buf ( n9756 , n5408 );
xor ( n9757 , n9755 , n9756 );
buf ( n9758 , n5409 );
xor ( n9759 , n9757 , n9758 );
buf ( n9760 , n5410 );
xor ( n9761 , n9759 , n9760 );
xor ( n9762 , n9740 , n9761 );
and ( n9763 , n9718 , n9762 );
xor ( n9764 , n9701 , n9763 );
xor ( n9765 , n9677 , n9764 );
xor ( n9766 , n8860 , n6681 );
not ( n9767 , n6583 );
buf ( n9768 , n5411 );
and ( n9769 , n9767 , n9768 );
buf ( n9770 , n5412 );
xor ( n9771 , n9770 , n9768 );
and ( n9772 , n9771 , n6583 );
or ( n9773 , n9769 , n9772 );
not ( n9774 , n6583 );
buf ( n9775 , n5413 );
and ( n9776 , n9774 , n9775 );
buf ( n9777 , n5414 );
xor ( n9778 , n9777 , n9775 );
and ( n9779 , n9778 , n6583 );
or ( n9780 , n9776 , n9779 );
xor ( n9781 , n9773 , n9780 );
buf ( n9782 , n5415 );
xor ( n9783 , n9781 , n9782 );
buf ( n9784 , n5416 );
xor ( n9785 , n9783 , n9784 );
buf ( n9786 , n5417 );
xor ( n9787 , n9785 , n9786 );
xor ( n9788 , n9766 , n9787 );
not ( n9789 , n6583 );
buf ( n9790 , n5418 );
and ( n9791 , n9789 , n9790 );
buf ( n9792 , n5419 );
xor ( n9793 , n9792 , n9790 );
and ( n9794 , n9793 , n6583 );
or ( n9795 , n9791 , n9794 );
not ( n9796 , n6583 );
buf ( n9797 , n5420 );
and ( n9798 , n9796 , n9797 );
buf ( n9799 , n5421 );
xor ( n9800 , n9799 , n9797 );
and ( n9801 , n9800 , n6583 );
or ( n9802 , n9798 , n9801 );
xor ( n9803 , n9795 , n9802 );
buf ( n9804 , n5422 );
xor ( n9805 , n9803 , n9804 );
buf ( n9806 , n5423 );
xor ( n9807 , n9805 , n9806 );
buf ( n9808 , n5424 );
xor ( n9809 , n9807 , n9808 );
xor ( n9810 , n6751 , n9809 );
not ( n9811 , n6583 );
buf ( n9812 , n5425 );
and ( n9813 , n9811 , n9812 );
buf ( n9814 , n5426 );
xor ( n9815 , n9814 , n9812 );
and ( n9816 , n9815 , n6583 );
or ( n9817 , n9813 , n9816 );
buf ( n9818 , n5427 );
xor ( n9819 , n9817 , n9818 );
buf ( n9820 , n5428 );
xor ( n9821 , n9819 , n9820 );
buf ( n9822 , n5429 );
xor ( n9823 , n9821 , n9822 );
buf ( n9824 , n5430 );
xor ( n9825 , n9823 , n9824 );
xor ( n9826 , n9810 , n9825 );
not ( n9827 , n9826 );
not ( n9828 , n6583 );
buf ( n9829 , n5431 );
and ( n9830 , n9828 , n9829 );
buf ( n9831 , n5432 );
xor ( n9832 , n9831 , n9829 );
and ( n9833 , n9832 , n6583 );
or ( n9834 , n9830 , n9833 );
not ( n9835 , n6583 );
buf ( n9836 , n5433 );
and ( n9837 , n9835 , n9836 );
buf ( n9838 , n5434 );
xor ( n9839 , n9838 , n9836 );
and ( n9840 , n9839 , n6583 );
or ( n9841 , n9837 , n9840 );
not ( n9842 , n6583 );
buf ( n9843 , n5435 );
and ( n9844 , n9842 , n9843 );
buf ( n9845 , n5436 );
xor ( n9846 , n9845 , n9843 );
and ( n9847 , n9846 , n6583 );
or ( n9848 , n9844 , n9847 );
xor ( n9849 , n9841 , n9848 );
buf ( n9850 , n5437 );
xor ( n9851 , n9849 , n9850 );
buf ( n9852 , n5438 );
xor ( n9853 , n9851 , n9852 );
buf ( n9854 , n5439 );
xor ( n9855 , n9853 , n9854 );
xor ( n9856 , n9834 , n9855 );
not ( n9857 , n6583 );
buf ( n9858 , n5440 );
and ( n9859 , n9857 , n9858 );
buf ( n9860 , n5441 );
xor ( n9861 , n9860 , n9858 );
and ( n9862 , n9861 , n6583 );
or ( n9863 , n9859 , n9862 );
not ( n9864 , n6583 );
buf ( n9865 , n5442 );
and ( n9866 , n9864 , n9865 );
buf ( n9867 , n5443 );
xor ( n9868 , n9867 , n9865 );
and ( n9869 , n9868 , n6583 );
or ( n9870 , n9866 , n9869 );
xor ( n9871 , n9863 , n9870 );
buf ( n9872 , n5444 );
xor ( n9873 , n9871 , n9872 );
buf ( n9874 , n5445 );
xor ( n9875 , n9873 , n9874 );
buf ( n9876 , n5446 );
xor ( n9877 , n9875 , n9876 );
xor ( n9878 , n9856 , n9877 );
and ( n9879 , n9827 , n9878 );
xor ( n9880 , n9788 , n9879 );
xor ( n9881 , n9765 , n9880 );
buf ( n9882 , n5447 );
not ( n9883 , n6583 );
buf ( n9884 , n5448 );
and ( n9885 , n9883 , n9884 );
buf ( n9886 , n5449 );
xor ( n9887 , n9886 , n9884 );
and ( n9888 , n9887 , n6583 );
or ( n9889 , n9885 , n9888 );
buf ( n9890 , n5450 );
xor ( n9891 , n9889 , n9890 );
buf ( n9892 , n5451 );
xor ( n9893 , n9891 , n9892 );
buf ( n9894 , n5452 );
xor ( n9895 , n9893 , n9894 );
buf ( n9896 , n5453 );
xor ( n9897 , n9895 , n9896 );
xor ( n9898 , n9882 , n9897 );
xor ( n9899 , n9898 , n9046 );
buf ( n9900 , n5454 );
not ( n9901 , n6583 );
buf ( n9902 , n5455 );
and ( n9903 , n9901 , n9902 );
buf ( n9904 , n5456 );
xor ( n9905 , n9904 , n9902 );
and ( n9906 , n9905 , n6583 );
or ( n9907 , n9903 , n9906 );
not ( n9908 , n6583 );
buf ( n9909 , n5457 );
and ( n9910 , n9908 , n9909 );
buf ( n9911 , n5458 );
xor ( n9912 , n9911 , n9909 );
and ( n9913 , n9912 , n6583 );
or ( n9914 , n9910 , n9913 );
xor ( n9915 , n9907 , n9914 );
xor ( n9916 , n9915 , n9163 );
buf ( n9917 , n5459 );
xor ( n9918 , n9916 , n9917 );
buf ( n9919 , n5460 );
xor ( n9920 , n9918 , n9919 );
xor ( n9921 , n9900 , n9920 );
not ( n9922 , n6583 );
buf ( n9923 , n5461 );
and ( n9924 , n9922 , n9923 );
buf ( n9925 , n5462 );
xor ( n9926 , n9925 , n9923 );
and ( n9927 , n9926 , n6583 );
or ( n9928 , n9924 , n9927 );
not ( n9929 , n6583 );
buf ( n9930 , n5463 );
and ( n9931 , n9929 , n9930 );
buf ( n9932 , n5464 );
xor ( n9933 , n9932 , n9930 );
and ( n9934 , n9933 , n6583 );
or ( n9935 , n9931 , n9934 );
xor ( n9936 , n9928 , n9935 );
buf ( n9937 , n5465 );
xor ( n9938 , n9936 , n9937 );
buf ( n9939 , n5466 );
xor ( n9940 , n9938 , n9939 );
buf ( n9941 , n5467 );
xor ( n9942 , n9940 , n9941 );
xor ( n9943 , n9921 , n9942 );
not ( n9944 , n9943 );
not ( n9945 , n6583 );
buf ( n9946 , n5468 );
and ( n9947 , n9945 , n9946 );
buf ( n9948 , n5469 );
xor ( n9949 , n9948 , n9946 );
and ( n9950 , n9949 , n6583 );
or ( n9951 , n9947 , n9950 );
not ( n9952 , n6583 );
buf ( n9953 , n5470 );
and ( n9954 , n9952 , n9953 );
buf ( n9955 , n5471 );
xor ( n9956 , n9955 , n9953 );
and ( n9957 , n9956 , n6583 );
or ( n9958 , n9954 , n9957 );
not ( n9959 , n6583 );
buf ( n9960 , n5472 );
and ( n9961 , n9959 , n9960 );
buf ( n9962 , n5473 );
xor ( n9963 , n9962 , n9960 );
and ( n9964 , n9963 , n6583 );
or ( n9965 , n9961 , n9964 );
xor ( n9966 , n9958 , n9965 );
buf ( n9967 , n5474 );
xor ( n9968 , n9966 , n9967 );
buf ( n9969 , n5475 );
xor ( n9970 , n9968 , n9969 );
buf ( n9971 , n5476 );
xor ( n9972 , n9970 , n9971 );
xor ( n9973 , n9951 , n9972 );
xor ( n9974 , n9973 , n7494 );
and ( n9975 , n9944 , n9974 );
xor ( n9976 , n9899 , n9975 );
xor ( n9977 , n9881 , n9976 );
xor ( n9978 , n9538 , n9977 );
and ( n9979 , n9024 , n9978 );
xor ( n9980 , n7953 , n9979 );
and ( n9981 , n9980 , n6584 );
or ( n9982 , n6587 , n9981 );
and ( n9983 , n6579 , n9982 );
buf ( n9984 , n9983 );
buf ( n9985 , n9984 );
buf ( n9986 , n6577 );
not ( n9987 , n9986 );
not ( n9988 , n6584 );
and ( n9989 , n9988 , n7467 );
not ( n9990 , n9978 );
buf ( n9991 , n5477 );
not ( n9992 , n6583 );
buf ( n9993 , n5478 );
and ( n9994 , n9992 , n9993 );
buf ( n9995 , n5479 );
xor ( n9996 , n9995 , n9993 );
and ( n9997 , n9996 , n6583 );
or ( n9998 , n9994 , n9997 );
not ( n9999 , n6583 );
buf ( n10000 , n5480 );
and ( n10001 , n9999 , n10000 );
buf ( n10002 , n5481 );
xor ( n10003 , n10002 , n10000 );
and ( n10004 , n10003 , n6583 );
or ( n10005 , n10001 , n10004 );
xor ( n10006 , n9998 , n10005 );
buf ( n10007 , n5482 );
xor ( n10008 , n10006 , n10007 );
buf ( n10009 , n5483 );
xor ( n10010 , n10008 , n10009 );
buf ( n10011 , n5484 );
xor ( n10012 , n10010 , n10011 );
xor ( n10013 , n9991 , n10012 );
not ( n10014 , n6583 );
buf ( n10015 , n5485 );
and ( n10016 , n10014 , n10015 );
buf ( n10017 , n5486 );
xor ( n10018 , n10017 , n10015 );
and ( n10019 , n10018 , n6583 );
or ( n10020 , n10016 , n10019 );
not ( n10021 , n6583 );
buf ( n10022 , n5487 );
and ( n10023 , n10021 , n10022 );
buf ( n10024 , n5488 );
xor ( n10025 , n10024 , n10022 );
and ( n10026 , n10025 , n6583 );
or ( n10027 , n10023 , n10026 );
xor ( n10028 , n10020 , n10027 );
buf ( n10029 , n5489 );
xor ( n10030 , n10028 , n10029 );
buf ( n10031 , n5490 );
xor ( n10032 , n10030 , n10031 );
buf ( n10033 , n5491 );
xor ( n10034 , n10032 , n10033 );
xor ( n10035 , n10013 , n10034 );
not ( n10036 , n6583 );
buf ( n10037 , n5492 );
and ( n10038 , n10036 , n10037 );
buf ( n10039 , n5493 );
xor ( n10040 , n10039 , n10037 );
and ( n10041 , n10040 , n6583 );
or ( n10042 , n10038 , n10041 );
not ( n10043 , n6583 );
buf ( n10044 , n5494 );
and ( n10045 , n10043 , n10044 );
buf ( n10046 , n5495 );
xor ( n10047 , n10046 , n10044 );
and ( n10048 , n10047 , n6583 );
or ( n10049 , n10045 , n10048 );
xor ( n10050 , n10042 , n10049 );
xor ( n10051 , n10050 , n7761 );
buf ( n10052 , n5496 );
xor ( n10053 , n10051 , n10052 );
buf ( n10054 , n5497 );
xor ( n10055 , n10053 , n10054 );
xor ( n10056 , n6726 , n10055 );
not ( n10057 , n6583 );
buf ( n10058 , n5498 );
and ( n10059 , n10057 , n10058 );
buf ( n10060 , n5499 );
xor ( n10061 , n10060 , n10058 );
and ( n10062 , n10061 , n6583 );
or ( n10063 , n10059 , n10062 );
xor ( n10064 , n10063 , n9439 );
buf ( n10065 , n5500 );
xor ( n10066 , n10064 , n10065 );
buf ( n10067 , n5501 );
xor ( n10068 , n10066 , n10067 );
buf ( n10069 , n5502 );
xor ( n10070 , n10068 , n10069 );
xor ( n10071 , n10056 , n10070 );
not ( n10072 , n10071 );
xor ( n10073 , n8894 , n9069 );
xor ( n10074 , n10073 , n9085 );
and ( n10075 , n10072 , n10074 );
xor ( n10076 , n10035 , n10075 );
buf ( n10077 , n5503 );
not ( n10078 , n6583 );
buf ( n10079 , n5504 );
and ( n10080 , n10078 , n10079 );
buf ( n10081 , n5505 );
xor ( n10082 , n10081 , n10079 );
and ( n10083 , n10082 , n6583 );
or ( n10084 , n10080 , n10083 );
not ( n10085 , n6583 );
buf ( n10086 , n5506 );
and ( n10087 , n10085 , n10086 );
buf ( n10088 , n5507 );
xor ( n10089 , n10088 , n10086 );
and ( n10090 , n10089 , n6583 );
or ( n10091 , n10087 , n10090 );
xor ( n10092 , n10084 , n10091 );
buf ( n10093 , n5508 );
xor ( n10094 , n10092 , n10093 );
buf ( n10095 , n5509 );
xor ( n10096 , n10094 , n10095 );
buf ( n10097 , n5510 );
xor ( n10098 , n10096 , n10097 );
xor ( n10099 , n10077 , n10098 );
not ( n10100 , n6583 );
buf ( n10101 , n5511 );
and ( n10102 , n10100 , n10101 );
buf ( n10103 , n5512 );
xor ( n10104 , n10103 , n10101 );
and ( n10105 , n10104 , n6583 );
or ( n10106 , n10102 , n10105 );
not ( n10107 , n6583 );
buf ( n10108 , n5513 );
and ( n10109 , n10107 , n10108 );
buf ( n10110 , n5514 );
xor ( n10111 , n10110 , n10108 );
and ( n10112 , n10111 , n6583 );
or ( n10113 , n10109 , n10112 );
xor ( n10114 , n10106 , n10113 );
buf ( n10115 , n5515 );
xor ( n10116 , n10114 , n10115 );
buf ( n10117 , n5516 );
xor ( n10118 , n10116 , n10117 );
buf ( n10119 , n5517 );
xor ( n10120 , n10118 , n10119 );
xor ( n10121 , n10099 , n10120 );
not ( n10122 , n6583 );
buf ( n10123 , n5518 );
and ( n10124 , n10122 , n10123 );
buf ( n10125 , n5519 );
xor ( n10126 , n10125 , n10123 );
and ( n10127 , n10126 , n6583 );
or ( n10128 , n10124 , n10127 );
not ( n10129 , n6583 );
buf ( n10130 , n5520 );
and ( n10131 , n10129 , n10130 );
buf ( n10132 , n5521 );
xor ( n10133 , n10132 , n10130 );
and ( n10134 , n10133 , n6583 );
or ( n10135 , n10131 , n10134 );
xor ( n10136 , n10128 , n10135 );
buf ( n10137 , n5522 );
xor ( n10138 , n10136 , n10137 );
buf ( n10139 , n5523 );
xor ( n10140 , n10138 , n10139 );
buf ( n10141 , n5524 );
xor ( n10142 , n10140 , n10141 );
xor ( n10143 , n9106 , n10142 );
xor ( n10144 , n10143 , n6659 );
not ( n10145 , n10144 );
xor ( n10146 , n8269 , n9244 );
not ( n10147 , n6583 );
buf ( n10148 , n5525 );
and ( n10149 , n10147 , n10148 );
buf ( n10150 , n5526 );
xor ( n10151 , n10150 , n10148 );
and ( n10152 , n10151 , n6583 );
or ( n10153 , n10149 , n10152 );
not ( n10154 , n6583 );
buf ( n10155 , n5527 );
and ( n10156 , n10154 , n10155 );
buf ( n10157 , n5528 );
xor ( n10158 , n10157 , n10155 );
and ( n10159 , n10158 , n6583 );
or ( n10160 , n10156 , n10159 );
xor ( n10161 , n10153 , n10160 );
xor ( n10162 , n10161 , n8661 );
buf ( n10163 , n5529 );
xor ( n10164 , n10162 , n10163 );
buf ( n10165 , n5530 );
xor ( n10166 , n10164 , n10165 );
xor ( n10167 , n10146 , n10166 );
and ( n10168 , n10145 , n10167 );
xor ( n10169 , n10121 , n10168 );
buf ( n10170 , n5531 );
xor ( n10171 , n10170 , n7996 );
not ( n10172 , n6583 );
buf ( n10173 , n5532 );
and ( n10174 , n10172 , n10173 );
buf ( n10175 , n5533 );
xor ( n10176 , n10175 , n10173 );
and ( n10177 , n10176 , n6583 );
or ( n10178 , n10174 , n10177 );
not ( n10179 , n6583 );
buf ( n10180 , n5534 );
and ( n10181 , n10179 , n10180 );
buf ( n10182 , n5535 );
xor ( n10183 , n10182 , n10180 );
and ( n10184 , n10183 , n6583 );
or ( n10185 , n10181 , n10184 );
xor ( n10186 , n10178 , n10185 );
buf ( n10187 , n5536 );
xor ( n10188 , n10186 , n10187 );
buf ( n10189 , n5537 );
xor ( n10190 , n10188 , n10189 );
buf ( n10191 , n5538 );
xor ( n10192 , n10190 , n10191 );
xor ( n10193 , n10171 , n10192 );
not ( n10194 , n10035 );
and ( n10195 , n10194 , n10071 );
xor ( n10196 , n10193 , n10195 );
xor ( n10197 , n10169 , n10196 );
buf ( n10198 , n5539 );
not ( n10199 , n6583 );
buf ( n10200 , n5540 );
and ( n10201 , n10199 , n10200 );
buf ( n10202 , n5541 );
xor ( n10203 , n10202 , n10200 );
and ( n10204 , n10203 , n6583 );
or ( n10205 , n10201 , n10204 );
not ( n10206 , n6583 );
buf ( n10207 , n5542 );
and ( n10208 , n10206 , n10207 );
buf ( n10209 , n5543 );
xor ( n10210 , n10209 , n10207 );
and ( n10211 , n10210 , n6583 );
or ( n10212 , n10208 , n10211 );
xor ( n10213 , n10205 , n10212 );
buf ( n10214 , n5544 );
xor ( n10215 , n10213 , n10214 );
buf ( n10216 , n5545 );
xor ( n10217 , n10215 , n10216 );
buf ( n10218 , n5546 );
xor ( n10219 , n10217 , n10218 );
xor ( n10220 , n10198 , n10219 );
xor ( n10221 , n10220 , n9715 );
not ( n10222 , n6583 );
buf ( n10223 , n5547 );
and ( n10224 , n10222 , n10223 );
buf ( n10225 , n5548 );
xor ( n10226 , n10225 , n10223 );
and ( n10227 , n10226 , n6583 );
or ( n10228 , n10224 , n10227 );
not ( n10229 , n6583 );
buf ( n10230 , n5549 );
and ( n10231 , n10229 , n10230 );
buf ( n10232 , n5550 );
xor ( n10233 , n10232 , n10230 );
and ( n10234 , n10233 , n6583 );
or ( n10235 , n10231 , n10234 );
xor ( n10236 , n10228 , n10235 );
buf ( n10237 , n5551 );
xor ( n10238 , n10236 , n10237 );
xor ( n10239 , n10238 , n7431 );
buf ( n10240 , n5552 );
xor ( n10241 , n10239 , n10240 );
xor ( n10242 , n9612 , n10241 );
xor ( n10243 , n10242 , n9739 );
not ( n10244 , n10243 );
buf ( n10245 , n5553 );
not ( n10246 , n6583 );
buf ( n10247 , n5554 );
and ( n10248 , n10246 , n10247 );
buf ( n10249 , n5555 );
xor ( n10250 , n10249 , n10247 );
and ( n10251 , n10250 , n6583 );
or ( n10252 , n10248 , n10251 );
buf ( n10253 , n5556 );
xor ( n10254 , n10252 , n10253 );
buf ( n10255 , n5557 );
xor ( n10256 , n10254 , n10255 );
buf ( n10257 , n5558 );
xor ( n10258 , n10256 , n10257 );
buf ( n10259 , n5559 );
xor ( n10260 , n10258 , n10259 );
xor ( n10261 , n10245 , n10260 );
not ( n10262 , n6583 );
buf ( n10263 , n5560 );
and ( n10264 , n10262 , n10263 );
buf ( n10265 , n5561 );
xor ( n10266 , n10265 , n10263 );
and ( n10267 , n10266 , n6583 );
or ( n10268 , n10264 , n10267 );
not ( n10269 , n6583 );
buf ( n10270 , n5562 );
and ( n10271 , n10269 , n10270 );
buf ( n10272 , n5563 );
xor ( n10273 , n10272 , n10270 );
and ( n10274 , n10273 , n6583 );
or ( n10275 , n10271 , n10274 );
xor ( n10276 , n10268 , n10275 );
buf ( n10277 , n5564 );
xor ( n10278 , n10276 , n10277 );
buf ( n10279 , n5565 );
xor ( n10280 , n10278 , n10279 );
buf ( n10281 , n5566 );
xor ( n10282 , n10280 , n10281 );
xor ( n10283 , n10261 , n10282 );
and ( n10284 , n10244 , n10283 );
xor ( n10285 , n10221 , n10284 );
xor ( n10286 , n10197 , n10285 );
buf ( n10287 , n5567 );
xor ( n10288 , n10287 , n9920 );
xor ( n10289 , n10288 , n9942 );
xor ( n10290 , n9015 , n8292 );
xor ( n10291 , n10290 , n9699 );
not ( n10292 , n10291 );
xor ( n10293 , n8634 , n8142 );
not ( n10294 , n6583 );
buf ( n10295 , n5568 );
and ( n10296 , n10294 , n10295 );
buf ( n10297 , n5569 );
xor ( n10298 , n10297 , n10295 );
and ( n10299 , n10298 , n6583 );
or ( n10300 , n10296 , n10299 );
buf ( n10301 , n5570 );
xor ( n10302 , n10300 , n10301 );
buf ( n10303 , n5571 );
xor ( n10304 , n10302 , n10303 );
buf ( n10305 , n5572 );
xor ( n10306 , n10304 , n10305 );
buf ( n10307 , n5573 );
xor ( n10308 , n10306 , n10307 );
xor ( n10309 , n10293 , n10308 );
and ( n10310 , n10292 , n10309 );
xor ( n10311 , n10289 , n10310 );
xor ( n10312 , n10286 , n10311 );
buf ( n10313 , n5574 );
not ( n10314 , n6583 );
buf ( n10315 , n5575 );
and ( n10316 , n10314 , n10315 );
buf ( n10317 , n5576 );
xor ( n10318 , n10317 , n10315 );
and ( n10319 , n10318 , n6583 );
or ( n10320 , n10316 , n10319 );
xor ( n10321 , n8213 , n10320 );
buf ( n10322 , n5577 );
xor ( n10323 , n10321 , n10322 );
buf ( n10324 , n5578 );
xor ( n10325 , n10323 , n10324 );
buf ( n10326 , n5579 );
xor ( n10327 , n10325 , n10326 );
xor ( n10328 , n10313 , n10327 );
not ( n10329 , n6583 );
buf ( n10330 , n5580 );
and ( n10331 , n10329 , n10330 );
buf ( n10332 , n5581 );
xor ( n10333 , n10332 , n10330 );
and ( n10334 , n10333 , n6583 );
or ( n10335 , n10331 , n10334 );
not ( n10336 , n6583 );
buf ( n10337 , n5582 );
and ( n10338 , n10336 , n10337 );
buf ( n10339 , n5583 );
xor ( n10340 , n10339 , n10337 );
and ( n10341 , n10340 , n6583 );
or ( n10342 , n10338 , n10341 );
xor ( n10343 , n10335 , n10342 );
buf ( n10344 , n5584 );
xor ( n10345 , n10343 , n10344 );
buf ( n10346 , n5585 );
xor ( n10347 , n10345 , n10346 );
buf ( n10348 , n5586 );
xor ( n10349 , n10347 , n10348 );
xor ( n10350 , n10328 , n10349 );
buf ( n10351 , n5587 );
not ( n10352 , n6583 );
buf ( n10353 , n5588 );
and ( n10354 , n10352 , n10353 );
buf ( n10355 , n5589 );
xor ( n10356 , n10355 , n10353 );
and ( n10357 , n10356 , n6583 );
or ( n10358 , n10354 , n10357 );
buf ( n10359 , n5590 );
xor ( n10360 , n10358 , n10359 );
buf ( n10361 , n5591 );
xor ( n10362 , n10360 , n10361 );
buf ( n10363 , n5592 );
xor ( n10364 , n10362 , n10363 );
buf ( n10365 , n5593 );
xor ( n10366 , n10364 , n10365 );
xor ( n10367 , n10351 , n10366 );
not ( n10368 , n6583 );
buf ( n10369 , n5594 );
and ( n10370 , n10368 , n10369 );
buf ( n10371 , n5595 );
xor ( n10372 , n10371 , n10369 );
and ( n10373 , n10372 , n6583 );
or ( n10374 , n10370 , n10373 );
not ( n10375 , n6583 );
buf ( n10376 , n5596 );
and ( n10377 , n10375 , n10376 );
buf ( n10378 , n5597 );
xor ( n10379 , n10378 , n10376 );
and ( n10380 , n10379 , n6583 );
or ( n10381 , n10377 , n10380 );
xor ( n10382 , n10374 , n10381 );
buf ( n10383 , n5598 );
xor ( n10384 , n10382 , n10383 );
buf ( n10385 , n5599 );
xor ( n10386 , n10384 , n10385 );
buf ( n10387 , n5600 );
xor ( n10388 , n10386 , n10387 );
xor ( n10389 , n10367 , n10388 );
not ( n10390 , n10389 );
not ( n10391 , n6583 );
buf ( n10392 , n5601 );
and ( n10393 , n10391 , n10392 );
buf ( n10394 , n5602 );
xor ( n10395 , n10394 , n10392 );
and ( n10396 , n10395 , n6583 );
or ( n10397 , n10393 , n10396 );
not ( n10398 , n6583 );
buf ( n10399 , n5603 );
and ( n10400 , n10398 , n10399 );
buf ( n10401 , n5604 );
xor ( n10402 , n10401 , n10399 );
and ( n10403 , n10402 , n6583 );
or ( n10404 , n10400 , n10403 );
xor ( n10405 , n10397 , n10404 );
buf ( n10406 , n5605 );
xor ( n10407 , n10405 , n10406 );
buf ( n10408 , n5606 );
xor ( n10409 , n10407 , n10408 );
buf ( n10410 , n5607 );
xor ( n10411 , n10409 , n10410 );
xor ( n10412 , n7827 , n10411 );
not ( n10413 , n6583 );
buf ( n10414 , n5608 );
and ( n10415 , n10413 , n10414 );
buf ( n10416 , n5609 );
xor ( n10417 , n10416 , n10414 );
and ( n10418 , n10417 , n6583 );
or ( n10419 , n10415 , n10418 );
not ( n10420 , n6583 );
buf ( n10421 , n5610 );
and ( n10422 , n10420 , n10421 );
buf ( n10423 , n5611 );
xor ( n10424 , n10423 , n10421 );
and ( n10425 , n10424 , n6583 );
or ( n10426 , n10422 , n10425 );
xor ( n10427 , n10419 , n10426 );
buf ( n10428 , n5612 );
xor ( n10429 , n10427 , n10428 );
buf ( n10430 , n5613 );
xor ( n10431 , n10429 , n10430 );
buf ( n10432 , n5614 );
xor ( n10433 , n10431 , n10432 );
xor ( n10434 , n10412 , n10433 );
and ( n10435 , n10390 , n10434 );
xor ( n10436 , n10350 , n10435 );
xor ( n10437 , n10312 , n10436 );
xor ( n10438 , n10076 , n10437 );
xor ( n10439 , n6962 , n9285 );
xor ( n10440 , n10439 , n9307 );
xor ( n10441 , n6760 , n9825 );
xor ( n10442 , n10441 , n7828 );
not ( n10443 , n10442 );
not ( n10444 , n6583 );
buf ( n10445 , n5615 );
and ( n10446 , n10444 , n10445 );
buf ( n10447 , n5616 );
xor ( n10448 , n10447 , n10445 );
and ( n10449 , n10448 , n6583 );
or ( n10450 , n10446 , n10449 );
xor ( n10451 , n10450 , n10012 );
xor ( n10452 , n10451 , n10034 );
and ( n10453 , n10443 , n10452 );
xor ( n10454 , n10440 , n10453 );
not ( n10455 , n6583 );
buf ( n10456 , n5617 );
and ( n10457 , n10455 , n10456 );
buf ( n10458 , n5618 );
xor ( n10459 , n10458 , n10456 );
and ( n10460 , n10459 , n6583 );
or ( n10461 , n10457 , n10460 );
not ( n10462 , n6583 );
buf ( n10463 , n5619 );
and ( n10464 , n10462 , n10463 );
buf ( n10465 , n5620 );
xor ( n10466 , n10465 , n10463 );
and ( n10467 , n10466 , n6583 );
or ( n10468 , n10464 , n10467 );
xor ( n10469 , n10461 , n10468 );
buf ( n10470 , n5621 );
xor ( n10471 , n10469 , n10470 );
buf ( n10472 , n5622 );
xor ( n10473 , n10471 , n10472 );
buf ( n10474 , n5623 );
xor ( n10475 , n10473 , n10474 );
xor ( n10476 , n7803 , n10475 );
not ( n10477 , n6583 );
buf ( n10478 , n5624 );
and ( n10479 , n10477 , n10478 );
buf ( n10480 , n5625 );
xor ( n10481 , n10480 , n10478 );
and ( n10482 , n10481 , n6583 );
or ( n10483 , n10479 , n10482 );
not ( n10484 , n6583 );
buf ( n10485 , n5626 );
and ( n10486 , n10484 , n10485 );
buf ( n10487 , n5627 );
xor ( n10488 , n10487 , n10485 );
and ( n10489 , n10488 , n6583 );
or ( n10490 , n10486 , n10489 );
xor ( n10491 , n10483 , n10490 );
buf ( n10492 , n5628 );
xor ( n10493 , n10491 , n10492 );
buf ( n10494 , n5629 );
xor ( n10495 , n10493 , n10494 );
buf ( n10496 , n5630 );
xor ( n10497 , n10495 , n10496 );
xor ( n10498 , n10476 , n10497 );
not ( n10499 , n6583 );
buf ( n10500 , n5631 );
and ( n10501 , n10499 , n10500 );
buf ( n10502 , n5632 );
xor ( n10503 , n10502 , n10500 );
and ( n10504 , n10503 , n6583 );
or ( n10505 , n10501 , n10504 );
xor ( n10506 , n10505 , n9560 );
xor ( n10507 , n10506 , n8807 );
not ( n10508 , n10507 );
buf ( n10509 , n5633 );
xor ( n10510 , n10509 , n9109 );
xor ( n10511 , n10510 , n8841 );
and ( n10512 , n10508 , n10511 );
xor ( n10513 , n10498 , n10512 );
xor ( n10514 , n10454 , n10513 );
buf ( n10515 , n5634 );
not ( n10516 , n6583 );
buf ( n10517 , n5635 );
and ( n10518 , n10516 , n10517 );
buf ( n10519 , n5636 );
xor ( n10520 , n10519 , n10517 );
and ( n10521 , n10520 , n6583 );
or ( n10522 , n10518 , n10521 );
buf ( n10523 , n5637 );
xor ( n10524 , n10522 , n10523 );
buf ( n10525 , n5638 );
xor ( n10526 , n10524 , n10525 );
buf ( n10527 , n5639 );
xor ( n10528 , n10526 , n10527 );
buf ( n10529 , n5640 );
xor ( n10530 , n10528 , n10529 );
xor ( n10531 , n10515 , n10530 );
not ( n10532 , n6583 );
buf ( n10533 , n5641 );
and ( n10534 , n10532 , n10533 );
buf ( n10535 , n5642 );
xor ( n10536 , n10535 , n10533 );
and ( n10537 , n10536 , n6583 );
or ( n10538 , n10534 , n10537 );
not ( n10539 , n6583 );
buf ( n10540 , n5643 );
and ( n10541 , n10539 , n10540 );
buf ( n10542 , n5644 );
xor ( n10543 , n10542 , n10540 );
and ( n10544 , n10543 , n6583 );
or ( n10545 , n10541 , n10544 );
xor ( n10546 , n10538 , n10545 );
buf ( n10547 , n5645 );
xor ( n10548 , n10546 , n10547 );
buf ( n10549 , n5646 );
xor ( n10550 , n10548 , n10549 );
buf ( n10551 , n5647 );
xor ( n10552 , n10550 , n10551 );
xor ( n10553 , n10531 , n10552 );
xor ( n10554 , n7814 , n10411 );
xor ( n10555 , n10554 , n10433 );
not ( n10556 , n10555 );
not ( n10557 , n6583 );
buf ( n10558 , n5648 );
and ( n10559 , n10557 , n10558 );
buf ( n10560 , n5649 );
xor ( n10561 , n10560 , n10558 );
and ( n10562 , n10561 , n6583 );
or ( n10563 , n10559 , n10562 );
not ( n10564 , n6583 );
buf ( n10565 , n5650 );
and ( n10566 , n10564 , n10565 );
buf ( n10567 , n5651 );
xor ( n10568 , n10567 , n10565 );
and ( n10569 , n10568 , n6583 );
or ( n10570 , n10566 , n10569 );
not ( n10571 , n6583 );
buf ( n10572 , n5652 );
and ( n10573 , n10571 , n10572 );
buf ( n10574 , n5653 );
xor ( n10575 , n10574 , n10572 );
and ( n10576 , n10575 , n6583 );
or ( n10577 , n10573 , n10576 );
xor ( n10578 , n10570 , n10577 );
buf ( n10579 , n5654 );
xor ( n10580 , n10578 , n10579 );
buf ( n10581 , n5655 );
xor ( n10582 , n10580 , n10581 );
buf ( n10583 , n5656 );
xor ( n10584 , n10582 , n10583 );
xor ( n10585 , n10563 , n10584 );
xor ( n10586 , n10585 , n10241 );
and ( n10587 , n10556 , n10586 );
xor ( n10588 , n10553 , n10587 );
xor ( n10589 , n10514 , n10588 );
not ( n10590 , n6583 );
buf ( n10591 , n5657 );
and ( n10592 , n10590 , n10591 );
buf ( n10593 , n5658 );
xor ( n10594 , n10593 , n10591 );
and ( n10595 , n10594 , n6583 );
or ( n10596 , n10592 , n10595 );
xor ( n10597 , n10596 , n7611 );
buf ( n10598 , n5659 );
xor ( n10599 , n10597 , n10598 );
buf ( n10600 , n5660 );
xor ( n10601 , n10599 , n10600 );
buf ( n10602 , n5661 );
xor ( n10603 , n10601 , n10602 );
xor ( n10604 , n7146 , n10603 );
not ( n10605 , n6583 );
buf ( n10606 , n5662 );
and ( n10607 , n10605 , n10606 );
buf ( n10608 , n5663 );
xor ( n10609 , n10608 , n10606 );
and ( n10610 , n10609 , n6583 );
or ( n10611 , n10607 , n10610 );
buf ( n10612 , n5664 );
xor ( n10613 , n10611 , n10612 );
buf ( n10614 , n5665 );
xor ( n10615 , n10613 , n10614 );
buf ( n10616 , n5666 );
xor ( n10617 , n10615 , n10616 );
buf ( n10618 , n5667 );
xor ( n10619 , n10617 , n10618 );
xor ( n10620 , n10604 , n10619 );
xor ( n10621 , n7918 , n8908 );
not ( n10622 , n6583 );
buf ( n10623 , n5668 );
and ( n10624 , n10622 , n10623 );
buf ( n10625 , n5669 );
xor ( n10626 , n10625 , n10623 );
and ( n10627 , n10626 , n6583 );
or ( n10628 , n10624 , n10627 );
not ( n10629 , n6583 );
buf ( n10630 , n5670 );
and ( n10631 , n10629 , n10630 );
buf ( n10632 , n5671 );
xor ( n10633 , n10632 , n10630 );
and ( n10634 , n10633 , n6583 );
or ( n10635 , n10631 , n10634 );
xor ( n10636 , n10628 , n10635 );
buf ( n10637 , n5672 );
xor ( n10638 , n10636 , n10637 );
buf ( n10639 , n5673 );
xor ( n10640 , n10638 , n10639 );
buf ( n10641 , n5674 );
xor ( n10642 , n10640 , n10641 );
xor ( n10643 , n10621 , n10642 );
not ( n10644 , n10643 );
not ( n10645 , n6583 );
buf ( n10646 , n5675 );
and ( n10647 , n10645 , n10646 );
buf ( n10648 , n5676 );
xor ( n10649 , n10648 , n10646 );
and ( n10650 , n10649 , n6583 );
or ( n10651 , n10647 , n10650 );
xor ( n10652 , n10651 , n8428 );
not ( n10653 , n6583 );
buf ( n10654 , n5677 );
and ( n10655 , n10653 , n10654 );
buf ( n10656 , n5678 );
xor ( n10657 , n10656 , n10654 );
and ( n10658 , n10657 , n6583 );
or ( n10659 , n10655 , n10658 );
not ( n10660 , n6583 );
buf ( n10661 , n5679 );
and ( n10662 , n10660 , n10661 );
buf ( n10663 , n5680 );
xor ( n10664 , n10663 , n10661 );
and ( n10665 , n10664 , n6583 );
or ( n10666 , n10662 , n10665 );
xor ( n10667 , n10659 , n10666 );
buf ( n10668 , n5681 );
xor ( n10669 , n10667 , n10668 );
buf ( n10670 , n5682 );
xor ( n10671 , n10669 , n10670 );
buf ( n10672 , n5683 );
xor ( n10673 , n10671 , n10672 );
xor ( n10674 , n10652 , n10673 );
and ( n10675 , n10644 , n10674 );
xor ( n10676 , n10620 , n10675 );
xor ( n10677 , n10589 , n10676 );
buf ( n10678 , n5684 );
not ( n10679 , n6583 );
buf ( n10680 , n5685 );
and ( n10681 , n10679 , n10680 );
buf ( n10682 , n5686 );
xor ( n10683 , n10682 , n10680 );
and ( n10684 , n10683 , n6583 );
or ( n10685 , n10681 , n10684 );
not ( n10686 , n6583 );
buf ( n10687 , n5687 );
and ( n10688 , n10686 , n10687 );
buf ( n10689 , n5688 );
xor ( n10690 , n10689 , n10687 );
and ( n10691 , n10690 , n6583 );
or ( n10692 , n10688 , n10691 );
xor ( n10693 , n10685 , n10692 );
xor ( n10694 , n10693 , n10170 );
buf ( n10695 , n5689 );
xor ( n10696 , n10694 , n10695 );
buf ( n10697 , n5690 );
xor ( n10698 , n10696 , n10697 );
xor ( n10699 , n10678 , n10698 );
xor ( n10700 , n10699 , n8932 );
not ( n10701 , n6583 );
buf ( n10702 , n5691 );
and ( n10703 , n10701 , n10702 );
buf ( n10704 , n5692 );
xor ( n10705 , n10704 , n10702 );
and ( n10706 , n10705 , n6583 );
or ( n10707 , n10703 , n10706 );
not ( n10708 , n6583 );
buf ( n10709 , n5693 );
and ( n10710 , n10708 , n10709 );
buf ( n10711 , n5694 );
xor ( n10712 , n10711 , n10709 );
and ( n10713 , n10712 , n6583 );
or ( n10714 , n10710 , n10713 );
not ( n10715 , n6583 );
buf ( n10716 , n5695 );
and ( n10717 , n10715 , n10716 );
buf ( n10718 , n5696 );
xor ( n10719 , n10718 , n10716 );
and ( n10720 , n10719 , n6583 );
or ( n10721 , n10717 , n10720 );
xor ( n10722 , n10714 , n10721 );
buf ( n10723 , n5697 );
xor ( n10724 , n10722 , n10723 );
buf ( n10725 , n5698 );
xor ( n10726 , n10724 , n10725 );
buf ( n10727 , n5699 );
xor ( n10728 , n10726 , n10727 );
xor ( n10729 , n10707 , n10728 );
xor ( n10730 , n10729 , n6752 );
not ( n10731 , n10730 );
xor ( n10732 , n8628 , n8142 );
xor ( n10733 , n10732 , n10308 );
and ( n10734 , n10731 , n10733 );
xor ( n10735 , n10700 , n10734 );
xor ( n10736 , n10677 , n10735 );
xor ( n10737 , n10438 , n10736 );
and ( n10738 , n9990 , n10737 );
xor ( n10739 , n9023 , n10738 );
and ( n10740 , n10739 , n6584 );
or ( n10741 , n9989 , n10740 );
and ( n10742 , n9987 , n10741 );
buf ( n10743 , n10742 );
buf ( n10744 , n10743 );
not ( n10745 , n6578 );
not ( n10746 , n6584 );
and ( n10747 , n10746 , n7845 );
xor ( n10748 , n7850 , n10433 );
xor ( n10749 , n10748 , n7029 );
not ( n10750 , n8483 );
and ( n10751 , n10750 , n8507 );
xor ( n10752 , n10749 , n10751 );
buf ( n10753 , n5700 );
xor ( n10754 , n10753 , n7390 );
xor ( n10755 , n10754 , n9262 );
buf ( n10756 , n5701 );
not ( n10757 , n6583 );
buf ( n10758 , n5702 );
and ( n10759 , n10757 , n10758 );
buf ( n10760 , n5703 );
xor ( n10761 , n10760 , n10758 );
and ( n10762 , n10761 , n6583 );
or ( n10763 , n10759 , n10762 );
not ( n10764 , n6583 );
buf ( n10765 , n5704 );
and ( n10766 , n10764 , n10765 );
buf ( n10767 , n5705 );
xor ( n10768 , n10767 , n10765 );
and ( n10769 , n10768 , n6583 );
or ( n10770 , n10766 , n10769 );
xor ( n10771 , n10763 , n10770 );
xor ( n10772 , n10771 , n10198 );
buf ( n10773 , n5706 );
xor ( n10774 , n10772 , n10773 );
buf ( n10775 , n5707 );
xor ( n10776 , n10774 , n10775 );
xor ( n10777 , n10756 , n10776 );
not ( n10778 , n6583 );
buf ( n10779 , n5708 );
and ( n10780 , n10778 , n10779 );
buf ( n10781 , n5709 );
xor ( n10782 , n10781 , n10779 );
and ( n10783 , n10782 , n6583 );
or ( n10784 , n10780 , n10783 );
not ( n10785 , n6583 );
buf ( n10786 , n5710 );
and ( n10787 , n10785 , n10786 );
buf ( n10788 , n5711 );
xor ( n10789 , n10788 , n10786 );
and ( n10790 , n10789 , n6583 );
or ( n10791 , n10787 , n10790 );
xor ( n10792 , n10784 , n10791 );
buf ( n10793 , n5712 );
xor ( n10794 , n10792 , n10793 );
buf ( n10795 , n5713 );
xor ( n10796 , n10794 , n10795 );
xor ( n10797 , n10796 , n9702 );
xor ( n10798 , n10777 , n10797 );
not ( n10799 , n10798 );
and ( n10800 , n10799 , n8106 );
xor ( n10801 , n10755 , n10800 );
not ( n10802 , n6583 );
buf ( n10803 , n5714 );
and ( n10804 , n10802 , n10803 );
buf ( n10805 , n5715 );
xor ( n10806 , n10805 , n10803 );
and ( n10807 , n10806 , n6583 );
or ( n10808 , n10804 , n10807 );
not ( n10809 , n6583 );
buf ( n10810 , n5716 );
and ( n10811 , n10809 , n10810 );
buf ( n10812 , n5717 );
xor ( n10813 , n10812 , n10810 );
and ( n10814 , n10813 , n6583 );
or ( n10815 , n10811 , n10814 );
xor ( n10816 , n10808 , n10815 );
buf ( n10817 , n5718 );
xor ( n10818 , n10816 , n10817 );
buf ( n10819 , n5719 );
xor ( n10820 , n10818 , n10819 );
buf ( n10821 , n5720 );
xor ( n10822 , n10820 , n10821 );
xor ( n10823 , n7122 , n10822 );
xor ( n10824 , n10823 , n10603 );
not ( n10825 , n6583 );
buf ( n10826 , n5721 );
and ( n10827 , n10825 , n10826 );
buf ( n10828 , n5722 );
xor ( n10829 , n10828 , n10826 );
and ( n10830 , n10829 , n6583 );
or ( n10831 , n10827 , n10830 );
not ( n10832 , n6583 );
buf ( n10833 , n5723 );
and ( n10834 , n10832 , n10833 );
buf ( n10835 , n5724 );
xor ( n10836 , n10835 , n10833 );
and ( n10837 , n10836 , n6583 );
or ( n10838 , n10834 , n10837 );
xor ( n10839 , n10831 , n10838 );
buf ( n10840 , n5725 );
xor ( n10841 , n10839 , n10840 );
buf ( n10842 , n5726 );
xor ( n10843 , n10841 , n10842 );
buf ( n10844 , n5727 );
xor ( n10845 , n10843 , n10844 );
xor ( n10846 , n7451 , n10845 );
not ( n10847 , n6583 );
buf ( n10848 , n5728 );
and ( n10849 , n10847 , n10848 );
buf ( n10850 , n5729 );
xor ( n10851 , n10850 , n10848 );
and ( n10852 , n10851 , n6583 );
or ( n10853 , n10849 , n10852 );
not ( n10854 , n6583 );
buf ( n10855 , n5730 );
and ( n10856 , n10854 , n10855 );
buf ( n10857 , n5731 );
xor ( n10858 , n10857 , n10855 );
and ( n10859 , n10858 , n6583 );
or ( n10860 , n10856 , n10859 );
xor ( n10861 , n10853 , n10860 );
buf ( n10862 , n5732 );
xor ( n10863 , n10861 , n10862 );
buf ( n10864 , n5733 );
xor ( n10865 , n10863 , n10864 );
buf ( n10866 , n6586 );
xor ( n10867 , n10865 , n10866 );
xor ( n10868 , n10846 , n10867 );
not ( n10869 , n10868 );
and ( n10870 , n10869 , n8251 );
xor ( n10871 , n10824 , n10870 );
xor ( n10872 , n10801 , n10871 );
not ( n10873 , n6583 );
buf ( n10874 , n5734 );
and ( n10875 , n10873 , n10874 );
buf ( n10876 , n5735 );
xor ( n10877 , n10876 , n10874 );
and ( n10878 , n10877 , n6583 );
or ( n10879 , n10875 , n10878 );
not ( n10880 , n6583 );
buf ( n10881 , n5736 );
and ( n10882 , n10880 , n10881 );
buf ( n10883 , n5737 );
xor ( n10884 , n10883 , n10881 );
and ( n10885 , n10884 , n6583 );
or ( n10886 , n10882 , n10885 );
xor ( n10887 , n10879 , n10886 );
buf ( n10888 , n5738 );
xor ( n10889 , n10887 , n10888 );
buf ( n10890 , n5739 );
xor ( n10891 , n10889 , n10890 );
buf ( n10892 , n5740 );
xor ( n10893 , n10891 , n10892 );
xor ( n10894 , n10527 , n10893 );
not ( n10895 , n6583 );
buf ( n10896 , n5741 );
and ( n10897 , n10895 , n10896 );
buf ( n10898 , n5742 );
xor ( n10899 , n10898 , n10896 );
and ( n10900 , n10899 , n6583 );
or ( n10901 , n10897 , n10900 );
not ( n10902 , n6583 );
buf ( n10903 , n5743 );
and ( n10904 , n10902 , n10903 );
buf ( n10905 , n5744 );
xor ( n10906 , n10905 , n10903 );
and ( n10907 , n10906 , n6583 );
or ( n10908 , n10904 , n10907 );
xor ( n10909 , n10901 , n10908 );
buf ( n10910 , n5745 );
xor ( n10911 , n10909 , n10910 );
buf ( n10912 , n5746 );
xor ( n10913 , n10911 , n10912 );
buf ( n10914 , n5747 );
xor ( n10915 , n10913 , n10914 );
xor ( n10916 , n10894 , n10915 );
xor ( n10917 , n10641 , n9085 );
xor ( n10918 , n10917 , n7406 );
not ( n10919 , n10918 );
and ( n10920 , n10919 , n8341 );
xor ( n10921 , n10916 , n10920 );
xor ( n10922 , n10872 , n10921 );
buf ( n10923 , n5748 );
not ( n10924 , n6583 );
buf ( n10925 , n5749 );
and ( n10926 , n10924 , n10925 );
buf ( n10927 , n5750 );
xor ( n10928 , n10927 , n10925 );
and ( n10929 , n10928 , n6583 );
or ( n10930 , n10926 , n10929 );
not ( n10931 , n6583 );
buf ( n10932 , n5751 );
and ( n10933 , n10931 , n10932 );
buf ( n10934 , n5752 );
xor ( n10935 , n10934 , n10932 );
and ( n10936 , n10935 , n6583 );
or ( n10937 , n10933 , n10936 );
xor ( n10938 , n10930 , n10937 );
buf ( n10939 , n5753 );
xor ( n10940 , n10938 , n10939 );
buf ( n10941 , n5754 );
xor ( n10942 , n10940 , n10941 );
buf ( n10943 , n5755 );
xor ( n10944 , n10942 , n10943 );
xor ( n10945 , n10923 , n10944 );
xor ( n10946 , n10945 , n9140 );
not ( n10947 , n10749 );
and ( n10948 , n10947 , n8483 );
xor ( n10949 , n10946 , n10948 );
xor ( n10950 , n10922 , n10949 );
not ( n10951 , n6583 );
buf ( n10952 , n5756 );
and ( n10953 , n10951 , n10952 );
buf ( n10954 , n5757 );
xor ( n10955 , n10954 , n10952 );
and ( n10956 , n10955 , n6583 );
or ( n10957 , n10953 , n10956 );
not ( n10958 , n6583 );
buf ( n10959 , n5758 );
and ( n10960 , n10958 , n10959 );
buf ( n10961 , n5759 );
xor ( n10962 , n10961 , n10959 );
and ( n10963 , n10962 , n6583 );
or ( n10964 , n10960 , n10963 );
xor ( n10965 , n10957 , n10964 );
buf ( n10966 , n5760 );
xor ( n10967 , n10965 , n10966 );
buf ( n10968 , n5761 );
xor ( n10969 , n10967 , n10968 );
buf ( n10970 , n5762 );
xor ( n10971 , n10969 , n10970 );
xor ( n10972 , n9228 , n10971 );
xor ( n10973 , n10972 , n6947 );
not ( n10974 , n10973 );
and ( n10975 , n10974 , n8607 );
xor ( n10976 , n8059 , n10975 );
xor ( n10977 , n10950 , n10976 );
xor ( n10978 , n10752 , n10977 );
not ( n10979 , n6583 );
buf ( n10980 , n5763 );
and ( n10981 , n10979 , n10980 );
buf ( n10982 , n5764 );
xor ( n10983 , n10982 , n10980 );
and ( n10984 , n10983 , n6583 );
or ( n10985 , n10981 , n10984 );
buf ( n10986 , n5765 );
xor ( n10987 , n10985 , n10986 );
buf ( n10988 , n5766 );
xor ( n10989 , n10987 , n10988 );
buf ( n10990 , n5767 );
xor ( n10991 , n10989 , n10990 );
buf ( n10992 , n5768 );
xor ( n10993 , n10991 , n10992 );
xor ( n10994 , n8303 , n10993 );
xor ( n10995 , n10994 , n9229 );
xor ( n10996 , n7118 , n10822 );
xor ( n10997 , n10996 , n10603 );
not ( n10998 , n10997 );
and ( n10999 , n10998 , n8636 );
xor ( n11000 , n10995 , n10999 );
not ( n11001 , n6583 );
buf ( n11002 , n5769 );
and ( n11003 , n11001 , n11002 );
buf ( n11004 , n5770 );
xor ( n11005 , n11004 , n11002 );
and ( n11006 , n11005 , n6583 );
or ( n11007 , n11003 , n11006 );
not ( n11008 , n6583 );
buf ( n11009 , n5771 );
and ( n11010 , n11008 , n11009 );
buf ( n11011 , n5772 );
xor ( n11012 , n11011 , n11009 );
and ( n11013 , n11012 , n6583 );
or ( n11014 , n11010 , n11013 );
not ( n11015 , n6583 );
buf ( n11016 , n5773 );
and ( n11017 , n11015 , n11016 );
buf ( n11018 , n5774 );
xor ( n11019 , n11018 , n11016 );
and ( n11020 , n11019 , n6583 );
or ( n11021 , n11017 , n11020 );
xor ( n11022 , n11014 , n11021 );
buf ( n11023 , n5775 );
xor ( n11024 , n11022 , n11023 );
buf ( n11025 , n5776 );
xor ( n11026 , n11024 , n11025 );
buf ( n11027 , n5777 );
xor ( n11028 , n11026 , n11027 );
xor ( n11029 , n11007 , n11028 );
xor ( n11030 , n11029 , n10366 );
buf ( n11031 , n5778 );
not ( n11032 , n6583 );
buf ( n11033 , n5779 );
and ( n11034 , n11032 , n11033 );
buf ( n11035 , n5780 );
xor ( n11036 , n11035 , n11033 );
and ( n11037 , n11036 , n6583 );
or ( n11038 , n11034 , n11037 );
not ( n11039 , n6583 );
buf ( n11040 , n5781 );
and ( n11041 , n11039 , n11040 );
buf ( n11042 , n5782 );
xor ( n11043 , n11042 , n11040 );
and ( n11044 , n11043 , n6583 );
or ( n11045 , n11041 , n11044 );
xor ( n11046 , n11038 , n11045 );
xor ( n11047 , n11046 , n9246 );
xor ( n11048 , n11047 , n10753 );
buf ( n11049 , n5783 );
xor ( n11050 , n11048 , n11049 );
xor ( n11051 , n11031 , n11050 );
not ( n11052 , n6583 );
buf ( n11053 , n5784 );
and ( n11054 , n11052 , n11053 );
buf ( n11055 , n5785 );
xor ( n11056 , n11055 , n11053 );
and ( n11057 , n11056 , n6583 );
or ( n11058 , n11054 , n11057 );
not ( n11059 , n6583 );
buf ( n11060 , n5786 );
and ( n11061 , n11059 , n11060 );
buf ( n11062 , n5787 );
xor ( n11063 , n11062 , n11060 );
and ( n11064 , n11063 , n6583 );
or ( n11065 , n11061 , n11064 );
xor ( n11066 , n11058 , n11065 );
buf ( n11067 , n5788 );
xor ( n11068 , n11066 , n11067 );
buf ( n11069 , n5789 );
xor ( n11070 , n11068 , n11069 );
buf ( n11071 , n5790 );
xor ( n11072 , n11070 , n11071 );
xor ( n11073 , n11051 , n11072 );
not ( n11074 , n11073 );
and ( n11075 , n11074 , n8684 );
xor ( n11076 , n11030 , n11075 );
xor ( n11077 , n11000 , n11076 );
xor ( n11078 , n9215 , n10971 );
xor ( n11079 , n11078 , n6947 );
not ( n11080 , n6583 );
buf ( n11081 , n5791 );
and ( n11082 , n11080 , n11081 );
buf ( n11083 , n5792 );
xor ( n11084 , n11083 , n11081 );
and ( n11085 , n11084 , n6583 );
or ( n11086 , n11082 , n11085 );
not ( n11087 , n6583 );
buf ( n11088 , n5793 );
and ( n11089 , n11087 , n11088 );
buf ( n11090 , n5794 );
xor ( n11091 , n11090 , n11088 );
and ( n11092 , n11091 , n6583 );
or ( n11093 , n11089 , n11092 );
xor ( n11094 , n11086 , n11093 );
buf ( n11095 , n5795 );
xor ( n11096 , n11094 , n11095 );
buf ( n11097 , n5796 );
xor ( n11098 , n11096 , n11097 );
buf ( n11099 , n5797 );
xor ( n11100 , n11098 , n11099 );
xor ( n11101 , n9377 , n11100 );
xor ( n11102 , n11101 , n10893 );
not ( n11103 , n11102 );
and ( n11104 , n11103 , n8767 );
xor ( n11105 , n11079 , n11104 );
xor ( n11106 , n11077 , n11105 );
not ( n11107 , n6583 );
buf ( n11108 , n5798 );
and ( n11109 , n11107 , n11108 );
buf ( n11110 , n5799 );
xor ( n11111 , n11110 , n11108 );
and ( n11112 , n11111 , n6583 );
or ( n11113 , n11109 , n11112 );
xor ( n11114 , n11113 , n10327 );
xor ( n11115 , n11114 , n10349 );
not ( n11116 , n6583 );
buf ( n11117 , n5800 );
and ( n11118 , n11116 , n11117 );
buf ( n11119 , n5801 );
xor ( n11120 , n11119 , n11117 );
and ( n11121 , n11120 , n6583 );
or ( n11122 , n11118 , n11121 );
xor ( n11123 , n11122 , n9511 );
xor ( n11124 , n11123 , n9533 );
not ( n11125 , n11124 );
and ( n11126 , n11125 , n8864 );
xor ( n11127 , n11115 , n11126 );
xor ( n11128 , n11106 , n11127 );
not ( n11129 , n6583 );
buf ( n11130 , n5802 );
and ( n11131 , n11129 , n11130 );
buf ( n11132 , n5803 );
xor ( n11133 , n11132 , n11130 );
and ( n11134 , n11133 , n6583 );
or ( n11135 , n11131 , n11134 );
not ( n11136 , n6583 );
buf ( n11137 , n5804 );
and ( n11138 , n11136 , n11137 );
buf ( n11139 , n5805 );
xor ( n11140 , n11139 , n11137 );
and ( n11141 , n11140 , n6583 );
or ( n11142 , n11138 , n11141 );
xor ( n11143 , n11135 , n11142 );
xor ( n11144 , n11143 , n10287 );
buf ( n11145 , n5806 );
xor ( n11146 , n11144 , n11145 );
xor ( n11147 , n11146 , n9900 );
xor ( n11148 , n9747 , n11147 );
not ( n11149 , n6583 );
buf ( n11150 , n5807 );
and ( n11151 , n11149 , n11150 );
buf ( n11152 , n5808 );
xor ( n11153 , n11152 , n11150 );
and ( n11154 , n11153 , n6583 );
or ( n11155 , n11151 , n11154 );
not ( n11156 , n6583 );
buf ( n11157 , n5809 );
and ( n11158 , n11156 , n11157 );
buf ( n11159 , n5810 );
xor ( n11160 , n11159 , n11157 );
and ( n11161 , n11160 , n6583 );
or ( n11162 , n11158 , n11161 );
xor ( n11163 , n11155 , n11162 );
buf ( n11164 , n5811 );
xor ( n11165 , n11163 , n11164 );
buf ( n11166 , n5812 );
xor ( n11167 , n11165 , n11166 );
buf ( n11168 , n5813 );
xor ( n11169 , n11167 , n11168 );
xor ( n11170 , n11148 , n11169 );
xor ( n11171 , n7843 , n10433 );
xor ( n11172 , n11171 , n7029 );
not ( n11173 , n11172 );
and ( n11174 , n11173 , n8976 );
xor ( n11175 , n11170 , n11174 );
xor ( n11176 , n11128 , n11175 );
xor ( n11177 , n10978 , n11176 );
not ( n11178 , n6583 );
buf ( n11179 , n5814 );
and ( n11180 , n11178 , n11179 );
buf ( n11181 , n5815 );
xor ( n11182 , n11181 , n11179 );
and ( n11183 , n11182 , n6583 );
or ( n11184 , n11180 , n11183 );
xor ( n11185 , n11184 , n10282 );
xor ( n11186 , n11185 , n8789 );
not ( n11187 , n6583 );
buf ( n11188 , n5816 );
and ( n11189 , n11187 , n11188 );
buf ( n11190 , n5817 );
xor ( n11191 , n11190 , n11188 );
and ( n11192 , n11191 , n6583 );
or ( n11193 , n11189 , n11192 );
xor ( n11194 , n11193 , n7677 );
xor ( n11195 , n11194 , n7686 );
not ( n11196 , n11195 );
buf ( n11197 , n5818 );
not ( n11198 , n6583 );
buf ( n11199 , n5819 );
and ( n11200 , n11198 , n11199 );
buf ( n11201 , n5820 );
xor ( n11202 , n11201 , n11199 );
and ( n11203 , n11202 , n6583 );
or ( n11204 , n11200 , n11203 );
not ( n11205 , n6583 );
buf ( n11206 , n5821 );
and ( n11207 , n11205 , n11206 );
buf ( n11208 , n5822 );
xor ( n11209 , n11208 , n11206 );
and ( n11210 , n11209 , n6583 );
or ( n11211 , n11207 , n11210 );
xor ( n11212 , n11204 , n11211 );
buf ( n11213 , n5823 );
xor ( n11214 , n11212 , n11213 );
buf ( n11215 , n5824 );
xor ( n11216 , n11214 , n11215 );
buf ( n11217 , n5825 );
xor ( n11218 , n11216 , n11217 );
xor ( n11219 , n11197 , n11218 );
xor ( n11220 , n11219 , n7782 );
and ( n11221 , n11196 , n11220 );
xor ( n11222 , n11186 , n11221 );
buf ( n11223 , n5826 );
xor ( n11224 , n11223 , n9855 );
xor ( n11225 , n11224 , n9877 );
not ( n11226 , n6583 );
buf ( n11227 , n5827 );
and ( n11228 , n11226 , n11227 );
buf ( n11229 , n5828 );
xor ( n11230 , n11229 , n11227 );
and ( n11231 , n11230 , n6583 );
or ( n11232 , n11228 , n11231 );
xor ( n11233 , n11232 , n10509 );
buf ( n11234 , n5829 );
xor ( n11235 , n11233 , n11234 );
buf ( n11236 , n5830 );
xor ( n11237 , n11235 , n11236 );
xor ( n11238 , n11237 , n9088 );
xor ( n11239 , n8516 , n11238 );
xor ( n11240 , n11239 , n9406 );
not ( n11241 , n11240 );
not ( n11242 , n6583 );
buf ( n11243 , n5831 );
and ( n11244 , n11242 , n11243 );
buf ( n11245 , n5832 );
xor ( n11246 , n11245 , n11243 );
and ( n11247 , n11246 , n6583 );
or ( n11248 , n11244 , n11247 );
xor ( n11249 , n11248 , n6774 );
xor ( n11250 , n11249 , n7980 );
and ( n11251 , n11241 , n11250 );
xor ( n11252 , n11225 , n11251 );
xor ( n11253 , n9383 , n11100 );
xor ( n11254 , n11253 , n10893 );
not ( n11255 , n6583 );
buf ( n11256 , n5833 );
and ( n11257 , n11255 , n11256 );
buf ( n11258 , n5834 );
xor ( n11259 , n11258 , n11256 );
and ( n11260 , n11259 , n6583 );
or ( n11261 , n11257 , n11260 );
not ( n11262 , n6583 );
buf ( n11263 , n5835 );
and ( n11264 , n11262 , n11263 );
buf ( n11265 , n5836 );
xor ( n11266 , n11265 , n11263 );
and ( n11267 , n11266 , n6583 );
or ( n11268 , n11264 , n11267 );
xor ( n11269 , n11261 , n11268 );
buf ( n11270 , n5837 );
xor ( n11271 , n11269 , n11270 );
buf ( n11272 , n5838 );
xor ( n11273 , n11271 , n11272 );
buf ( n11274 , n5839 );
xor ( n11275 , n11273 , n11274 );
xor ( n11276 , n7275 , n11275 );
xor ( n11277 , n11276 , n6797 );
not ( n11278 , n11277 );
not ( n11279 , n6583 );
buf ( n11280 , n5840 );
and ( n11281 , n11279 , n11280 );
buf ( n11282 , n5841 );
xor ( n11283 , n11282 , n11280 );
and ( n11284 , n11283 , n6583 );
or ( n11285 , n11281 , n11284 );
xor ( n11286 , n11285 , n7298 );
buf ( n11287 , n5842 );
xor ( n11288 , n11286 , n11287 );
buf ( n11289 , n5843 );
xor ( n11290 , n11288 , n11289 );
buf ( n11291 , n5844 );
xor ( n11292 , n11290 , n11291 );
xor ( n11293 , n10359 , n11292 );
not ( n11294 , n6583 );
buf ( n11295 , n5845 );
and ( n11296 , n11294 , n11295 );
buf ( n11297 , n5846 );
xor ( n11298 , n11297 , n11295 );
and ( n11299 , n11298 , n6583 );
or ( n11300 , n11296 , n11299 );
not ( n11301 , n6583 );
buf ( n11302 , n5847 );
and ( n11303 , n11301 , n11302 );
buf ( n11304 , n5848 );
xor ( n11305 , n11304 , n11302 );
and ( n11306 , n11305 , n6583 );
or ( n11307 , n11303 , n11306 );
xor ( n11308 , n11300 , n11307 );
buf ( n11309 , n5849 );
xor ( n11310 , n11308 , n11309 );
buf ( n11311 , n5850 );
xor ( n11312 , n11310 , n11311 );
buf ( n11313 , n5851 );
xor ( n11314 , n11312 , n11313 );
xor ( n11315 , n11293 , n11314 );
and ( n11316 , n11278 , n11315 );
xor ( n11317 , n11254 , n11316 );
xor ( n11318 , n11252 , n11317 );
buf ( n11319 , n5852 );
xor ( n11320 , n11113 , n11319 );
xor ( n11321 , n11320 , n10313 );
buf ( n11322 , n5853 );
xor ( n11323 , n11321 , n11322 );
buf ( n11324 , n5854 );
xor ( n11325 , n11323 , n11324 );
xor ( n11326 , n8481 , n11325 );
not ( n11327 , n6583 );
buf ( n11328 , n5855 );
and ( n11329 , n11327 , n11328 );
buf ( n11330 , n5856 );
xor ( n11331 , n11330 , n11328 );
and ( n11332 , n11331 , n6583 );
or ( n11333 , n11329 , n11332 );
not ( n11334 , n6583 );
buf ( n11335 , n5857 );
and ( n11336 , n11334 , n11335 );
buf ( n11337 , n5858 );
xor ( n11338 , n11337 , n11335 );
and ( n11339 , n11338 , n6583 );
or ( n11340 , n11336 , n11339 );
xor ( n11341 , n11333 , n11340 );
buf ( n11342 , n5859 );
xor ( n11343 , n11341 , n11342 );
buf ( n11344 , n5860 );
xor ( n11345 , n11343 , n11344 );
buf ( n11346 , n5861 );
xor ( n11347 , n11345 , n11346 );
xor ( n11348 , n11326 , n11347 );
xor ( n11349 , n9393 , n8841 );
xor ( n11350 , n11349 , n8863 );
not ( n11351 , n11350 );
not ( n11352 , n6583 );
buf ( n11353 , n5862 );
and ( n11354 , n11352 , n11353 );
buf ( n11355 , n5863 );
xor ( n11356 , n11355 , n11353 );
and ( n11357 , n11356 , n6583 );
or ( n11358 , n11354 , n11357 );
xor ( n11359 , n11358 , n8886 );
xor ( n11360 , n11359 , n8908 );
and ( n11361 , n11351 , n11360 );
xor ( n11362 , n11348 , n11361 );
xor ( n11363 , n11318 , n11362 );
xor ( n11364 , n6614 , n8340 );
xor ( n11365 , n11364 , n8270 );
xor ( n11366 , n9503 , n6918 );
not ( n11367 , n6583 );
buf ( n11368 , n5864 );
and ( n11369 , n11367 , n11368 );
buf ( n11370 , n5865 );
xor ( n11371 , n11370 , n11368 );
and ( n11372 , n11371 , n6583 );
or ( n11373 , n11369 , n11372 );
not ( n11374 , n6583 );
buf ( n11375 , n5866 );
and ( n11376 , n11374 , n11375 );
buf ( n11377 , n5867 );
xor ( n11378 , n11377 , n11375 );
and ( n11379 , n11378 , n6583 );
or ( n11380 , n11376 , n11379 );
xor ( n11381 , n11373 , n11380 );
buf ( n11382 , n5868 );
xor ( n11383 , n11381 , n11382 );
xor ( n11384 , n11383 , n9882 );
buf ( n11385 , n5869 );
xor ( n11386 , n11384 , n11385 );
xor ( n11387 , n11366 , n11386 );
not ( n11388 , n11387 );
xor ( n11389 , n8698 , n10308 );
not ( n11390 , n6583 );
buf ( n11391 , n5870 );
and ( n11392 , n11390 , n11391 );
buf ( n11393 , n5871 );
xor ( n11394 , n11393 , n11391 );
and ( n11395 , n11394 , n6583 );
or ( n11396 , n11392 , n11395 );
not ( n11397 , n6583 );
buf ( n11398 , n5872 );
and ( n11399 , n11397 , n11398 );
buf ( n11400 , n5873 );
xor ( n11401 , n11400 , n11398 );
and ( n11402 , n11401 , n6583 );
or ( n11403 , n11399 , n11402 );
xor ( n11404 , n11396 , n11403 );
buf ( n11405 , n5874 );
xor ( n11406 , n11404 , n11405 );
buf ( n11407 , n5875 );
xor ( n11408 , n11406 , n11407 );
buf ( n11409 , n5876 );
xor ( n11410 , n11408 , n11409 );
xor ( n11411 , n11389 , n11410 );
and ( n11412 , n11388 , n11411 );
xor ( n11413 , n11365 , n11412 );
xor ( n11414 , n11363 , n11413 );
xor ( n11415 , n6680 , n9598 );
not ( n11416 , n6583 );
buf ( n11417 , n5877 );
and ( n11418 , n11416 , n11417 );
buf ( n11419 , n5878 );
xor ( n11420 , n11419 , n11417 );
and ( n11421 , n11420 , n6583 );
or ( n11422 , n11418 , n11421 );
not ( n11423 , n6583 );
buf ( n11424 , n5879 );
and ( n11425 , n11423 , n11424 );
buf ( n11426 , n5880 );
xor ( n11427 , n11426 , n11424 );
and ( n11428 , n11427 , n6583 );
or ( n11429 , n11425 , n11428 );
xor ( n11430 , n11422 , n11429 );
buf ( n11431 , n5881 );
xor ( n11432 , n11430 , n11431 );
buf ( n11433 , n5882 );
xor ( n11434 , n11432 , n11433 );
buf ( n11435 , n5883 );
xor ( n11436 , n11434 , n11435 );
xor ( n11437 , n11415 , n11436 );
not ( n11438 , n11186 );
and ( n11439 , n11438 , n11195 );
xor ( n11440 , n11437 , n11439 );
xor ( n11441 , n11414 , n11440 );
xor ( n11442 , n11222 , n11441 );
xor ( n11443 , n7821 , n10411 );
xor ( n11444 , n11443 , n10433 );
buf ( n11445 , n5884 );
not ( n11446 , n6583 );
buf ( n11447 , n5885 );
and ( n11448 , n11446 , n11447 );
buf ( n11449 , n5886 );
xor ( n11450 , n11449 , n11447 );
and ( n11451 , n11450 , n6583 );
or ( n11452 , n11448 , n11451 );
xor ( n11453 , n11452 , n11248 );
buf ( n11454 , n5887 );
xor ( n11455 , n11453 , n11454 );
buf ( n11456 , n5888 );
xor ( n11457 , n11455 , n11456 );
buf ( n11458 , n5889 );
xor ( n11459 , n11457 , n11458 );
xor ( n11460 , n11445 , n11459 );
not ( n11461 , n6583 );
buf ( n11462 , n5890 );
and ( n11463 , n11461 , n11462 );
buf ( n11464 , n5891 );
xor ( n11465 , n11464 , n11462 );
and ( n11466 , n11465 , n6583 );
or ( n11467 , n11463 , n11466 );
xor ( n11468 , n11467 , n7960 );
buf ( n11469 , n5892 );
xor ( n11470 , n11468 , n11469 );
buf ( n11471 , n5893 );
xor ( n11472 , n11470 , n11471 );
buf ( n11473 , n5894 );
xor ( n11474 , n11472 , n11473 );
xor ( n11475 , n11460 , n11474 );
not ( n11476 , n11475 );
buf ( n11477 , n5895 );
not ( n11478 , n6583 );
buf ( n11479 , n5896 );
and ( n11480 , n11478 , n11479 );
buf ( n11481 , n5897 );
xor ( n11482 , n11481 , n11479 );
and ( n11483 , n11482 , n6583 );
or ( n11484 , n11480 , n11483 );
not ( n11485 , n6583 );
buf ( n11486 , n5898 );
and ( n11487 , n11485 , n11486 );
buf ( n11488 , n5899 );
xor ( n11489 , n11488 , n11486 );
and ( n11490 , n11489 , n6583 );
or ( n11491 , n11487 , n11490 );
xor ( n11492 , n11484 , n11491 );
xor ( n11493 , n11492 , n10077 );
buf ( n11494 , n5900 );
xor ( n11495 , n11493 , n11494 );
buf ( n11496 , n5901 );
xor ( n11497 , n11495 , n11496 );
xor ( n11498 , n11477 , n11497 );
not ( n11499 , n6583 );
buf ( n11500 , n5902 );
and ( n11501 , n11499 , n11500 );
buf ( n11502 , n5903 );
xor ( n11503 , n11502 , n11500 );
and ( n11504 , n11503 , n6583 );
or ( n11505 , n11501 , n11504 );
buf ( n11506 , n5904 );
xor ( n11507 , n11505 , n11506 );
buf ( n11508 , n5905 );
xor ( n11509 , n11507 , n11508 );
buf ( n11510 , n5906 );
xor ( n11511 , n11509 , n11510 );
buf ( n11512 , n5907 );
xor ( n11513 , n11511 , n11512 );
xor ( n11514 , n11498 , n11513 );
and ( n11515 , n11476 , n11514 );
xor ( n11516 , n11444 , n11515 );
not ( n11517 , n6583 );
buf ( n11518 , n5908 );
and ( n11519 , n11517 , n11518 );
buf ( n11520 , n5909 );
xor ( n11521 , n11520 , n11518 );
and ( n11522 , n11521 , n6583 );
or ( n11523 , n11519 , n11522 );
xor ( n11524 , n11523 , n7862 );
buf ( n11525 , n5910 );
xor ( n11526 , n11524 , n11525 );
buf ( n11527 , n5911 );
xor ( n11528 , n11526 , n11527 );
xor ( n11529 , n11528 , n7152 );
xor ( n11530 , n7328 , n11529 );
not ( n11531 , n6583 );
buf ( n11532 , n5912 );
and ( n11533 , n11531 , n11532 );
buf ( n11534 , n5913 );
xor ( n11535 , n11534 , n11532 );
and ( n11536 , n11535 , n6583 );
or ( n11537 , n11533 , n11536 );
xor ( n11538 , n11537 , n9318 );
buf ( n11539 , n5914 );
xor ( n11540 , n11538 , n11539 );
buf ( n11541 , n5915 );
xor ( n11542 , n11540 , n11541 );
buf ( n11543 , n5916 );
xor ( n11544 , n11542 , n11543 );
xor ( n11545 , n11530 , n11544 );
buf ( n11546 , n5917 );
not ( n11547 , n6583 );
buf ( n11548 , n5918 );
and ( n11549 , n11547 , n11548 );
buf ( n11550 , n5919 );
xor ( n11551 , n11550 , n11548 );
and ( n11552 , n11551 , n6583 );
or ( n11553 , n11549 , n11552 );
buf ( n11554 , n5920 );
xor ( n11555 , n11553 , n11554 );
buf ( n11556 , n5921 );
xor ( n11557 , n11555 , n11556 );
buf ( n11558 , n5922 );
xor ( n11559 , n11557 , n11558 );
xor ( n11560 , n11559 , n10756 );
xor ( n11561 , n11546 , n11560 );
xor ( n11562 , n11561 , n10944 );
not ( n11563 , n11562 );
buf ( n11564 , n5923 );
xor ( n11565 , n11564 , n10698 );
xor ( n11566 , n11565 , n8932 );
and ( n11567 , n11563 , n11566 );
xor ( n11568 , n11545 , n11567 );
xor ( n11569 , n11516 , n11568 );
not ( n11570 , n6583 );
buf ( n11571 , n5924 );
and ( n11572 , n11570 , n11571 );
buf ( n11573 , n5925 );
xor ( n11574 , n11573 , n11571 );
and ( n11575 , n11574 , n6583 );
or ( n11576 , n11572 , n11575 );
not ( n11577 , n6583 );
buf ( n11578 , n5926 );
and ( n11579 , n11577 , n11578 );
buf ( n11580 , n5927 );
xor ( n11581 , n11580 , n11578 );
and ( n11582 , n11581 , n6583 );
or ( n11583 , n11579 , n11582 );
xor ( n11584 , n11576 , n11583 );
buf ( n11585 , n5928 );
xor ( n11586 , n11584 , n11585 );
buf ( n11587 , n5929 );
xor ( n11588 , n11586 , n11587 );
buf ( n11589 , n5930 );
xor ( n11590 , n11588 , n11589 );
xor ( n11591 , n9062 , n11590 );
not ( n11592 , n6583 );
buf ( n11593 , n5931 );
and ( n11594 , n11592 , n11593 );
buf ( n11595 , n5932 );
xor ( n11596 , n11595 , n11593 );
and ( n11597 , n11596 , n6583 );
or ( n11598 , n11594 , n11597 );
xor ( n11599 , n10505 , n11598 );
buf ( n11600 , n5933 );
xor ( n11601 , n11599 , n11600 );
xor ( n11602 , n11601 , n9539 );
buf ( n11603 , n5934 );
xor ( n11604 , n11602 , n11603 );
xor ( n11605 , n11591 , n11604 );
buf ( n11606 , n5935 );
not ( n11607 , n6583 );
buf ( n11608 , n5936 );
and ( n11609 , n11607 , n11608 );
buf ( n11610 , n5937 );
xor ( n11611 , n11610 , n11608 );
and ( n11612 , n11611 , n6583 );
or ( n11613 , n11609 , n11612 );
not ( n11614 , n6583 );
buf ( n11615 , n5938 );
and ( n11616 , n11614 , n11615 );
buf ( n11617 , n5939 );
xor ( n11618 , n11617 , n11615 );
and ( n11619 , n11618 , n6583 );
or ( n11620 , n11616 , n11619 );
xor ( n11621 , n11613 , n11620 );
buf ( n11622 , n5940 );
xor ( n11623 , n11621 , n11622 );
buf ( n11624 , n5941 );
xor ( n11625 , n11623 , n11624 );
xor ( n11626 , n11625 , n6875 );
xor ( n11627 , n11606 , n11626 );
xor ( n11628 , n11627 , n9511 );
not ( n11629 , n11628 );
not ( n11630 , n6583 );
buf ( n11631 , n5942 );
and ( n11632 , n11630 , n11631 );
buf ( n11633 , n5943 );
xor ( n11634 , n11633 , n11631 );
and ( n11635 , n11634 , n6583 );
or ( n11636 , n11632 , n11635 );
not ( n11637 , n6583 );
buf ( n11638 , n5944 );
and ( n11639 , n11637 , n11638 );
buf ( n11640 , n5945 );
xor ( n11641 , n11640 , n11638 );
and ( n11642 , n11641 , n6583 );
or ( n11643 , n11639 , n11642 );
xor ( n11644 , n11636 , n11643 );
buf ( n11645 , n5946 );
xor ( n11646 , n11644 , n11645 );
buf ( n11647 , n5947 );
xor ( n11648 , n11646 , n11647 );
buf ( n11649 , n5948 );
xor ( n11650 , n11648 , n11649 );
xor ( n11651 , n8804 , n11650 );
xor ( n11652 , n11651 , n7368 );
and ( n11653 , n11629 , n11652 );
xor ( n11654 , n11605 , n11653 );
xor ( n11655 , n11569 , n11654 );
not ( n11656 , n6583 );
buf ( n11657 , n5949 );
and ( n11658 , n11656 , n11657 );
buf ( n11659 , n5950 );
xor ( n11660 , n11659 , n11657 );
and ( n11661 , n11660 , n6583 );
or ( n11662 , n11658 , n11661 );
xor ( n11663 , n11662 , n10619 );
not ( n11664 , n6583 );
buf ( n11665 , n5951 );
and ( n11666 , n11664 , n11665 );
buf ( n11667 , n5952 );
xor ( n11668 , n11667 , n11665 );
and ( n11669 , n11668 , n6583 );
or ( n11670 , n11666 , n11669 );
not ( n11671 , n6583 );
buf ( n11672 , n5953 );
and ( n11673 , n11671 , n11672 );
buf ( n11674 , n5954 );
xor ( n11675 , n11674 , n11672 );
and ( n11676 , n11675 , n6583 );
or ( n11677 , n11673 , n11676 );
xor ( n11678 , n11670 , n11677 );
buf ( n11679 , n5955 );
xor ( n11680 , n11678 , n11679 );
buf ( n11681 , n5956 );
xor ( n11682 , n11680 , n11681 );
buf ( n11683 , n5957 );
xor ( n11684 , n11682 , n11683 );
xor ( n11685 , n11663 , n11684 );
buf ( n11686 , n5958 );
xor ( n11687 , n11686 , n7579 );
xor ( n11688 , n11687 , n7600 );
not ( n11689 , n11688 );
not ( n11690 , n6583 );
buf ( n11691 , n5959 );
and ( n11692 , n11690 , n11691 );
buf ( n11693 , n5960 );
xor ( n11694 , n11693 , n11691 );
and ( n11695 , n11694 , n6583 );
or ( n11696 , n11692 , n11695 );
not ( n11697 , n6583 );
buf ( n11698 , n5961 );
and ( n11699 , n11697 , n11698 );
buf ( n11700 , n5962 );
xor ( n11701 , n11700 , n11698 );
and ( n11702 , n11701 , n6583 );
or ( n11703 , n11699 , n11702 );
xor ( n11704 , n11696 , n11703 );
buf ( n11705 , n5963 );
xor ( n11706 , n11704 , n11705 );
buf ( n11707 , n5964 );
xor ( n11708 , n11706 , n11707 );
buf ( n11709 , n5965 );
xor ( n11710 , n11708 , n11709 );
xor ( n11711 , n8754 , n11710 );
xor ( n11712 , n11711 , n8460 );
and ( n11713 , n11689 , n11712 );
xor ( n11714 , n11685 , n11713 );
xor ( n11715 , n11655 , n11714 );
xor ( n11716 , n6608 , n8340 );
xor ( n11717 , n11716 , n8270 );
buf ( n11718 , n5966 );
not ( n11719 , n6583 );
buf ( n11720 , n5967 );
and ( n11721 , n11719 , n11720 );
buf ( n11722 , n5968 );
xor ( n11723 , n11722 , n11720 );
and ( n11724 , n11723 , n6583 );
or ( n11725 , n11721 , n11724 );
not ( n11726 , n6583 );
buf ( n11727 , n5969 );
and ( n11728 , n11726 , n11727 );
buf ( n11729 , n5970 );
xor ( n11730 , n11729 , n11727 );
and ( n11731 , n11730 , n6583 );
or ( n11732 , n11728 , n11731 );
xor ( n11733 , n11725 , n11732 );
buf ( n11734 , n5971 );
xor ( n11735 , n11733 , n11734 );
buf ( n11736 , n5972 );
xor ( n11737 , n11735 , n11736 );
buf ( n11738 , n5973 );
xor ( n11739 , n11737 , n11738 );
xor ( n11740 , n11718 , n11739 );
not ( n11741 , n6583 );
buf ( n11742 , n5974 );
and ( n11743 , n11741 , n11742 );
buf ( n11744 , n5975 );
xor ( n11745 , n11744 , n11742 );
and ( n11746 , n11745 , n6583 );
or ( n11747 , n11743 , n11746 );
not ( n11748 , n6583 );
buf ( n11749 , n5976 );
and ( n11750 , n11748 , n11749 );
buf ( n11751 , n5977 );
xor ( n11752 , n11751 , n11749 );
and ( n11753 , n11752 , n6583 );
or ( n11754 , n11750 , n11753 );
xor ( n11755 , n11747 , n11754 );
buf ( n11756 , n5978 );
xor ( n11757 , n11755 , n11756 );
buf ( n11758 , n5979 );
xor ( n11759 , n11757 , n11758 );
buf ( n11760 , n5980 );
xor ( n11761 , n11759 , n11760 );
xor ( n11762 , n11740 , n11761 );
not ( n11763 , n11762 );
buf ( n11764 , n5981 );
xor ( n11765 , n11764 , n9455 );
not ( n11766 , n6583 );
buf ( n11767 , n5982 );
and ( n11768 , n11766 , n11767 );
buf ( n11769 , n5983 );
xor ( n11770 , n11769 , n11767 );
and ( n11771 , n11770 , n6583 );
or ( n11772 , n11768 , n11771 );
not ( n11773 , n6583 );
buf ( n11774 , n5984 );
and ( n11775 , n11773 , n11774 );
buf ( n11776 , n5985 );
xor ( n11777 , n11776 , n11774 );
and ( n11778 , n11777 , n6583 );
or ( n11779 , n11775 , n11778 );
xor ( n11780 , n11772 , n11779 );
buf ( n11781 , n5986 );
xor ( n11782 , n11780 , n11781 );
buf ( n11783 , n5987 );
xor ( n11784 , n11782 , n11783 );
buf ( n11785 , n5988 );
xor ( n11786 , n11784 , n11785 );
xor ( n11787 , n11765 , n11786 );
and ( n11788 , n11763 , n11787 );
xor ( n11789 , n11717 , n11788 );
xor ( n11790 , n11715 , n11789 );
xor ( n11791 , n11442 , n11790 );
not ( n11792 , n11791 );
not ( n11793 , n6583 );
buf ( n11794 , n5989 );
and ( n11795 , n11793 , n11794 );
buf ( n11796 , n5990 );
xor ( n11797 , n11796 , n11794 );
and ( n11798 , n11797 , n6583 );
or ( n11799 , n11795 , n11798 );
xor ( n11800 , n11799 , n11122 );
buf ( n11801 , n5991 );
xor ( n11802 , n11800 , n11801 );
xor ( n11803 , n11802 , n9496 );
buf ( n11804 , n5992 );
xor ( n11805 , n11803 , n11804 );
xor ( n11806 , n7260 , n11805 );
xor ( n11807 , n11806 , n11275 );
xor ( n11808 , n11622 , n6896 );
xor ( n11809 , n11808 , n6918 );
not ( n11810 , n11809 );
xor ( n11811 , n10773 , n10219 );
xor ( n11812 , n11811 , n9715 );
and ( n11813 , n11810 , n11812 );
xor ( n11814 , n11807 , n11813 );
not ( n11815 , n6583 );
buf ( n11816 , n5993 );
and ( n11817 , n11815 , n11816 );
buf ( n11818 , n5994 );
xor ( n11819 , n11818 , n11816 );
and ( n11820 , n11819 , n6583 );
or ( n11821 , n11817 , n11820 );
xor ( n11822 , n11821 , n7029 );
xor ( n11823 , n11822 , n7051 );
not ( n11824 , n11807 );
and ( n11825 , n11824 , n11809 );
xor ( n11826 , n11823 , n11825 );
xor ( n11827 , n11038 , n7390 );
xor ( n11828 , n11827 , n9262 );
buf ( n11829 , n5995 );
xor ( n11830 , n11829 , n9787 );
not ( n11831 , n6583 );
buf ( n11832 , n5996 );
and ( n11833 , n11831 , n11832 );
buf ( n11834 , n5997 );
xor ( n11835 , n11834 , n11832 );
and ( n11836 , n11835 , n6583 );
or ( n11837 , n11833 , n11836 );
not ( n11838 , n6583 );
buf ( n11839 , n5998 );
and ( n11840 , n11838 , n11839 );
buf ( n11841 , n5999 );
xor ( n11842 , n11841 , n11839 );
and ( n11843 , n11842 , n6583 );
or ( n11844 , n11840 , n11843 );
xor ( n11845 , n11837 , n11844 );
xor ( n11846 , n11845 , n11546 );
buf ( n11847 , n6000 );
xor ( n11848 , n11846 , n11847 );
buf ( n11849 , n6001 );
xor ( n11850 , n11848 , n11849 );
xor ( n11851 , n11830 , n11850 );
not ( n11852 , n11851 );
not ( n11853 , n6583 );
buf ( n11854 , n6002 );
and ( n11855 , n11853 , n11854 );
buf ( n11856 , n6003 );
xor ( n11857 , n11856 , n11854 );
and ( n11858 , n11857 , n6583 );
or ( n11859 , n11855 , n11858 );
xor ( n11860 , n11859 , n7473 );
buf ( n11861 , n6004 );
xor ( n11862 , n11860 , n11861 );
buf ( n11863 , n6005 );
xor ( n11864 , n11862 , n11863 );
buf ( n11865 , n6006 );
xor ( n11866 , n11864 , n11865 );
xor ( n11867 , n7004 , n11866 );
xor ( n11868 , n11867 , n10845 );
and ( n11869 , n11852 , n11868 );
xor ( n11870 , n11828 , n11869 );
xor ( n11871 , n11826 , n11870 );
not ( n11872 , n6583 );
buf ( n11873 , n6007 );
and ( n11874 , n11872 , n11873 );
buf ( n11875 , n6008 );
xor ( n11876 , n11875 , n11873 );
and ( n11877 , n11876 , n6583 );
or ( n11878 , n11874 , n11877 );
not ( n11879 , n6583 );
buf ( n11880 , n6009 );
and ( n11881 , n11879 , n11880 );
buf ( n11882 , n6010 );
xor ( n11883 , n11882 , n11880 );
and ( n11884 , n11883 , n6583 );
or ( n11885 , n11881 , n11884 );
xor ( n11886 , n11878 , n11885 );
buf ( n11887 , n6011 );
xor ( n11888 , n11886 , n11887 );
buf ( n11889 , n6012 );
xor ( n11890 , n11888 , n11889 );
buf ( n11891 , n6013 );
xor ( n11892 , n11890 , n11891 );
xor ( n11893 , n7037 , n11892 );
not ( n11894 , n6583 );
buf ( n11895 , n6014 );
and ( n11896 , n11894 , n11895 );
buf ( n11897 , n6015 );
xor ( n11898 , n11897 , n11895 );
and ( n11899 , n11898 , n6583 );
or ( n11900 , n11896 , n11899 );
xor ( n11901 , n9951 , n11900 );
buf ( n11902 , n6016 );
xor ( n11903 , n11901 , n11902 );
buf ( n11904 , n6017 );
xor ( n11905 , n11903 , n11904 );
buf ( n11906 , n6018 );
xor ( n11907 , n11905 , n11906 );
xor ( n11908 , n11893 , n11907 );
xor ( n11909 , n9754 , n11147 );
xor ( n11910 , n11909 , n11169 );
not ( n11911 , n11910 );
xor ( n11912 , n11600 , n9560 );
xor ( n11913 , n11912 , n8807 );
and ( n11914 , n11911 , n11913 );
xor ( n11915 , n11908 , n11914 );
xor ( n11916 , n11871 , n11915 );
not ( n11917 , n6583 );
buf ( n11918 , n6019 );
and ( n11919 , n11917 , n11918 );
buf ( n11920 , n6020 );
xor ( n11921 , n11920 , n11918 );
and ( n11922 , n11921 , n6583 );
or ( n11923 , n11919 , n11922 );
xor ( n11924 , n11923 , n7428 );
xor ( n11925 , n11924 , n7579 );
xor ( n11926 , n10342 , n8250 );
not ( n11927 , n6583 );
buf ( n11928 , n6021 );
and ( n11929 , n11927 , n11928 );
buf ( n11930 , n6022 );
xor ( n11931 , n11930 , n11928 );
and ( n11932 , n11931 , n6583 );
or ( n11933 , n11929 , n11932 );
not ( n11934 , n6583 );
buf ( n11935 , n6023 );
and ( n11936 , n11934 , n11935 );
buf ( n11937 , n6024 );
xor ( n11938 , n11937 , n11935 );
and ( n11939 , n11938 , n6583 );
or ( n11940 , n11936 , n11939 );
xor ( n11941 , n11933 , n11940 );
buf ( n11942 , n6025 );
xor ( n11943 , n11941 , n11942 );
buf ( n11944 , n6026 );
xor ( n11945 , n11943 , n11944 );
buf ( n11946 , n6027 );
xor ( n11947 , n11945 , n11946 );
xor ( n11948 , n11926 , n11947 );
not ( n11949 , n11948 );
buf ( n11950 , n6028 );
xor ( n11951 , n11950 , n6636 );
xor ( n11952 , n11951 , n9018 );
and ( n11953 , n11949 , n11952 );
xor ( n11954 , n11925 , n11953 );
xor ( n11955 , n11916 , n11954 );
xor ( n11956 , n7967 , n7828 );
xor ( n11957 , n11956 , n7851 );
not ( n11958 , n6583 );
buf ( n11959 , n6029 );
and ( n11960 , n11958 , n11959 );
buf ( n11961 , n6030 );
xor ( n11962 , n11961 , n11959 );
and ( n11963 , n11962 , n6583 );
or ( n11964 , n11960 , n11963 );
not ( n11965 , n6583 );
buf ( n11966 , n6031 );
and ( n11967 , n11965 , n11966 );
buf ( n11968 , n6032 );
xor ( n11969 , n11968 , n11966 );
and ( n11970 , n11969 , n6583 );
or ( n11971 , n11967 , n11970 );
xor ( n11972 , n11964 , n11971 );
buf ( n11973 , n6033 );
xor ( n11974 , n11972 , n11973 );
buf ( n11975 , n6034 );
xor ( n11976 , n11974 , n11975 );
buf ( n11977 , n6035 );
xor ( n11978 , n11976 , n11977 );
xor ( n11979 , n7703 , n11978 );
not ( n11980 , n6583 );
buf ( n11981 , n6036 );
and ( n11982 , n11980 , n11981 );
buf ( n11983 , n6037 );
xor ( n11984 , n11983 , n11981 );
and ( n11985 , n11984 , n6583 );
or ( n11986 , n11982 , n11985 );
buf ( n11987 , n6038 );
xor ( n11988 , n11986 , n11987 );
xor ( n11989 , n11988 , n11197 );
buf ( n11990 , n6039 );
xor ( n11991 , n11989 , n11990 );
buf ( n11992 , n6040 );
xor ( n11993 , n11991 , n11992 );
xor ( n11994 , n11979 , n11993 );
not ( n11995 , n11994 );
not ( n11996 , n6583 );
buf ( n11997 , n6041 );
and ( n11998 , n11996 , n11997 );
buf ( n11999 , n6042 );
xor ( n12000 , n11999 , n11997 );
and ( n12001 , n12000 , n6583 );
or ( n12002 , n11998 , n12001 );
not ( n12003 , n6583 );
buf ( n12004 , n6043 );
and ( n12005 , n12003 , n12004 );
buf ( n12006 , n6044 );
xor ( n12007 , n12006 , n12004 );
and ( n12008 , n12007 , n6583 );
or ( n12009 , n12005 , n12008 );
xor ( n12010 , n12002 , n12009 );
buf ( n12011 , n6045 );
xor ( n12012 , n12010 , n12011 );
xor ( n12013 , n12012 , n11477 );
buf ( n12014 , n6046 );
xor ( n12015 , n12013 , n12014 );
xor ( n12016 , n7184 , n12015 );
not ( n12017 , n6583 );
buf ( n12018 , n6047 );
and ( n12019 , n12017 , n12018 );
buf ( n12020 , n6048 );
xor ( n12021 , n12020 , n12018 );
and ( n12022 , n12021 , n6583 );
or ( n12023 , n12019 , n12022 );
not ( n12024 , n6583 );
buf ( n12025 , n6049 );
and ( n12026 , n12024 , n12025 );
buf ( n12027 , n6050 );
xor ( n12028 , n12027 , n12025 );
and ( n12029 , n12028 , n6583 );
or ( n12030 , n12026 , n12029 );
xor ( n12031 , n12023 , n12030 );
buf ( n12032 , n6051 );
xor ( n12033 , n12031 , n12032 );
buf ( n12034 , n6052 );
xor ( n12035 , n12033 , n12034 );
buf ( n12036 , n6053 );
xor ( n12037 , n12035 , n12036 );
xor ( n12038 , n12016 , n12037 );
and ( n12039 , n11995 , n12038 );
xor ( n12040 , n11957 , n12039 );
xor ( n12041 , n11955 , n12040 );
xor ( n12042 , n11814 , n12041 );
buf ( n12043 , n6054 );
xor ( n12044 , n12043 , n7267 );
xor ( n12045 , n12044 , n7289 );
not ( n12046 , n6583 );
buf ( n12047 , n6055 );
and ( n12048 , n12046 , n12047 );
buf ( n12049 , n6056 );
xor ( n12050 , n12049 , n12047 );
and ( n12051 , n12050 , n6583 );
or ( n12052 , n12048 , n12051 );
not ( n12053 , n6583 );
buf ( n12054 , n6057 );
and ( n12055 , n12053 , n12054 );
buf ( n12056 , n6058 );
xor ( n12057 , n12056 , n12054 );
and ( n12058 , n12057 , n6583 );
or ( n12059 , n12055 , n12058 );
xor ( n12060 , n12052 , n12059 );
buf ( n12061 , n6059 );
xor ( n12062 , n12060 , n12061 );
xor ( n12063 , n12062 , n10923 );
buf ( n12064 , n6060 );
xor ( n12065 , n12063 , n12064 );
xor ( n12066 , n7883 , n12065 );
not ( n12067 , n6583 );
buf ( n12068 , n6061 );
and ( n12069 , n12067 , n12068 );
buf ( n12070 , n6062 );
xor ( n12071 , n12070 , n12068 );
and ( n12072 , n12071 , n6583 );
or ( n12073 , n12069 , n12072 );
xor ( n12074 , n12073 , n9119 );
buf ( n12075 , n6063 );
xor ( n12076 , n12074 , n12075 );
buf ( n12077 , n6064 );
xor ( n12078 , n12076 , n12077 );
buf ( n12079 , n6065 );
xor ( n12080 , n12078 , n12079 );
xor ( n12081 , n12066 , n12080 );
not ( n12082 , n12081 );
xor ( n12083 , n10529 , n10893 );
xor ( n12084 , n12083 , n10915 );
and ( n12085 , n12082 , n12084 );
xor ( n12086 , n12045 , n12085 );
xor ( n12087 , n7511 , n9615 );
xor ( n12088 , n12087 , n8584 );
not ( n12089 , n6583 );
buf ( n12090 , n6066 );
and ( n12091 , n12089 , n12090 );
buf ( n12092 , n6067 );
xor ( n12093 , n12092 , n12090 );
and ( n12094 , n12093 , n6583 );
or ( n12095 , n12091 , n12094 );
xor ( n12096 , n6782 , n12095 );
buf ( n12097 , n6068 );
xor ( n12098 , n12096 , n12097 );
buf ( n12099 , n6069 );
xor ( n12100 , n12098 , n12099 );
buf ( n12101 , n6070 );
xor ( n12102 , n12100 , n12101 );
xor ( n12103 , n9043 , n12102 );
not ( n12104 , n6583 );
buf ( n12105 , n6071 );
and ( n12106 , n12104 , n12105 );
buf ( n12107 , n6072 );
xor ( n12108 , n12107 , n12105 );
and ( n12109 , n12108 , n6583 );
or ( n12110 , n12106 , n12109 );
not ( n12111 , n6583 );
buf ( n12112 , n6073 );
and ( n12113 , n12111 , n12112 );
buf ( n12114 , n6074 );
xor ( n12115 , n12114 , n12112 );
and ( n12116 , n12115 , n6583 );
or ( n12117 , n12113 , n12116 );
xor ( n12118 , n12110 , n12117 );
buf ( n12119 , n6075 );
buf ( n12120 , n12119 );
xor ( n12121 , n12118 , n12120 );
buf ( n12122 , n6076 );
xor ( n12123 , n12121 , n12122 );
buf ( n12124 , n6077 );
xor ( n12125 , n12123 , n12124 );
xor ( n12126 , n12103 , n12125 );
not ( n12127 , n12126 );
xor ( n12128 , n7979 , n7828 );
xor ( n12129 , n12128 , n7851 );
and ( n12130 , n12127 , n12129 );
xor ( n12131 , n12088 , n12130 );
xor ( n12132 , n12086 , n12131 );
not ( n12133 , n6583 );
buf ( n12134 , n6078 );
and ( n12135 , n12133 , n12134 );
buf ( n12136 , n6079 );
xor ( n12137 , n12136 , n12134 );
and ( n12138 , n12137 , n6583 );
or ( n12139 , n12135 , n12138 );
not ( n12140 , n6583 );
buf ( n12141 , n6080 );
and ( n12142 , n12140 , n12141 );
buf ( n12143 , n6081 );
xor ( n12144 , n12143 , n12141 );
and ( n12145 , n12144 , n6583 );
or ( n12146 , n12142 , n12145 );
xor ( n12147 , n12139 , n12146 );
xor ( n12148 , n12147 , n7392 );
buf ( n12149 , n6082 );
xor ( n12150 , n12148 , n12149 );
buf ( n12151 , n6083 );
xor ( n12152 , n12150 , n12151 );
xor ( n12153 , n11645 , n12152 );
xor ( n12154 , n11923 , n8252 );
buf ( n12155 , n6084 );
xor ( n12156 , n12154 , n12155 );
buf ( n12157 , n6085 );
xor ( n12158 , n12156 , n12157 );
buf ( n12159 , n6086 );
xor ( n12160 , n12158 , n12159 );
xor ( n12161 , n12153 , n12160 );
xor ( n12162 , n7683 , n6615 );
xor ( n12163 , n12162 , n6636 );
not ( n12164 , n12163 );
xor ( n12165 , n9597 , n7737 );
xor ( n12166 , n12165 , n7759 );
and ( n12167 , n12164 , n12166 );
xor ( n12168 , n12161 , n12167 );
xor ( n12169 , n12132 , n12168 );
xor ( n12170 , n8287 , n10166 );
not ( n12171 , n6583 );
buf ( n12172 , n6087 );
and ( n12173 , n12171 , n12172 );
buf ( n12174 , n6088 );
xor ( n12175 , n12174 , n12172 );
and ( n12176 , n12175 , n6583 );
or ( n12177 , n12173 , n12176 );
not ( n12178 , n6583 );
buf ( n12179 , n6089 );
and ( n12180 , n12178 , n12179 );
buf ( n12181 , n6090 );
xor ( n12182 , n12181 , n12179 );
and ( n12183 , n12182 , n6583 );
or ( n12184 , n12180 , n12183 );
xor ( n12185 , n12177 , n12184 );
buf ( n12186 , n6091 );
xor ( n12187 , n12185 , n12186 );
buf ( n12188 , n6092 );
xor ( n12189 , n12187 , n12188 );
buf ( n12190 , n6093 );
xor ( n12191 , n12189 , n12190 );
xor ( n12192 , n12170 , n12191 );
buf ( n12193 , n6094 );
buf ( n12194 , n12193 );
xor ( n12195 , n12194 , n10552 );
xor ( n12196 , n12195 , n9109 );
not ( n12197 , n12196 );
xor ( n12198 , n11738 , n6727 );
not ( n12199 , n6583 );
buf ( n12200 , n6095 );
and ( n12201 , n12199 , n12200 );
buf ( n12202 , n6096 );
xor ( n12203 , n12202 , n12200 );
and ( n12204 , n12203 , n6583 );
or ( n12205 , n12201 , n12204 );
buf ( n12206 , n6097 );
xor ( n12207 , n12205 , n12206 );
buf ( n12208 , n6098 );
xor ( n12209 , n12207 , n12208 );
buf ( n12210 , n6099 );
xor ( n12211 , n12209 , n12210 );
buf ( n12212 , n6100 );
xor ( n12213 , n12211 , n12212 );
xor ( n12214 , n12198 , n12213 );
and ( n12215 , n12197 , n12214 );
xor ( n12216 , n12192 , n12215 );
xor ( n12217 , n12169 , n12216 );
xor ( n12218 , n11508 , n10120 );
xor ( n12219 , n12218 , n10012 );
buf ( n12220 , n6101 );
not ( n12221 , n6583 );
buf ( n12222 , n6102 );
and ( n12223 , n12221 , n12222 );
buf ( n12224 , n6103 );
xor ( n12225 , n12224 , n12222 );
and ( n12226 , n12225 , n6583 );
or ( n12227 , n12223 , n12226 );
buf ( n12228 , n6104 );
xor ( n12229 , n12227 , n12228 );
xor ( n12230 , n12229 , n9457 );
buf ( n12231 , n6105 );
xor ( n12232 , n12230 , n12231 );
buf ( n12233 , n6106 );
xor ( n12234 , n12232 , n12233 );
xor ( n12235 , n12220 , n12234 );
xor ( n12236 , n12235 , n6896 );
not ( n12237 , n12236 );
xor ( n12238 , n10583 , n7009 );
xor ( n12239 , n12238 , n7452 );
and ( n12240 , n12237 , n12239 );
xor ( n12241 , n12219 , n12240 );
xor ( n12242 , n12217 , n12241 );
xor ( n12243 , n12042 , n12242 );
and ( n12244 , n11792 , n12243 );
xor ( n12245 , n11177 , n12244 );
and ( n12246 , n12245 , n6584 );
or ( n12247 , n10747 , n12246 );
and ( n12248 , n10745 , n12247 );
buf ( n12249 , n12248 );
buf ( n12250 , n12249 );
not ( n12251 , n6578 );
not ( n12252 , n6584 );
buf ( n12253 , n6107 );
and ( n12254 , n12252 , n12253 );
not ( n12255 , n6583 );
buf ( n12256 , n6108 );
and ( n12257 , n12255 , n12256 );
buf ( n12258 , n6109 );
xor ( n12259 , n12258 , n12256 );
and ( n12260 , n12259 , n6583 );
or ( n12261 , n12257 , n12260 );
xor ( n12262 , n12261 , n8482 );
xor ( n12263 , n12262 , n11028 );
not ( n12264 , n6583 );
buf ( n12265 , n6110 );
and ( n12266 , n12264 , n12265 );
buf ( n12267 , n6111 );
xor ( n12268 , n12267 , n12265 );
and ( n12269 , n12268 , n6583 );
or ( n12270 , n12266 , n12269 );
xor ( n12271 , n12270 , n9340 );
not ( n12272 , n6583 );
buf ( n12273 , n6112 );
and ( n12274 , n12272 , n12273 );
buf ( n12275 , n6113 );
xor ( n12276 , n12275 , n12273 );
and ( n12277 , n12276 , n6583 );
or ( n12278 , n12274 , n12277 );
not ( n12279 , n6583 );
buf ( n12280 , n6114 );
and ( n12281 , n12279 , n12280 );
buf ( n12282 , n6115 );
xor ( n12283 , n12282 , n12280 );
and ( n12284 , n12283 , n6583 );
or ( n12285 , n12281 , n12284 );
xor ( n12286 , n12278 , n12285 );
buf ( n12287 , n6116 );
xor ( n12288 , n12286 , n12287 );
buf ( n12289 , n6117 );
xor ( n12290 , n12288 , n12289 );
buf ( n12291 , n6118 );
xor ( n12292 , n12290 , n12291 );
xor ( n12293 , n12271 , n12292 );
not ( n12294 , n12293 );
not ( n12295 , n6583 );
buf ( n12296 , n6119 );
and ( n12297 , n12295 , n12296 );
buf ( n12298 , n6120 );
xor ( n12299 , n12298 , n12296 );
and ( n12300 , n12299 , n6583 );
or ( n12301 , n12297 , n12300 );
xor ( n12302 , n10707 , n12301 );
buf ( n12303 , n6121 );
xor ( n12304 , n12302 , n12303 );
buf ( n12305 , n6122 );
xor ( n12306 , n12304 , n12305 );
buf ( n12307 , n6123 );
xor ( n12308 , n12306 , n12307 );
xor ( n12309 , n10492 , n12308 );
not ( n12310 , n6583 );
buf ( n12311 , n6124 );
and ( n12312 , n12310 , n12311 );
buf ( n12313 , n6125 );
xor ( n12314 , n12313 , n12311 );
and ( n12315 , n12314 , n6583 );
or ( n12316 , n12312 , n12315 );
buf ( n12317 , n6126 );
xor ( n12318 , n12316 , n12317 );
buf ( n12319 , n6127 );
xor ( n12320 , n12318 , n12319 );
buf ( n12321 , n6128 );
xor ( n12322 , n12320 , n12321 );
xor ( n12323 , n12322 , n6731 );
xor ( n12324 , n12309 , n12323 );
and ( n12325 , n12294 , n12324 );
xor ( n12326 , n12263 , n12325 );
not ( n12327 , n6583 );
buf ( n12328 , n6129 );
and ( n12329 , n12327 , n12328 );
buf ( n12330 , n6130 );
xor ( n12331 , n12330 , n12328 );
and ( n12332 , n12331 , n6583 );
or ( n12333 , n12329 , n12332 );
not ( n12334 , n6583 );
buf ( n12335 , n6131 );
and ( n12336 , n12334 , n12335 );
buf ( n12337 , n6132 );
xor ( n12338 , n12337 , n12335 );
and ( n12339 , n12338 , n6583 );
or ( n12340 , n12336 , n12339 );
xor ( n12341 , n12333 , n12340 );
buf ( n12342 , n6133 );
xor ( n12343 , n12341 , n12342 );
buf ( n12344 , n6134 );
xor ( n12345 , n12343 , n12344 );
buf ( n12346 , n6135 );
xor ( n12347 , n12345 , n12346 );
xor ( n12348 , n8035 , n12347 );
xor ( n12349 , n12348 , n9639 );
not ( n12350 , n6583 );
buf ( n12351 , n6136 );
and ( n12352 , n12350 , n12351 );
buf ( n12353 , n6137 );
xor ( n12354 , n12353 , n12351 );
and ( n12355 , n12354 , n6583 );
or ( n12356 , n12352 , n12355 );
xor ( n12357 , n12356 , n8766 );
not ( n12358 , n6583 );
buf ( n12359 , n6138 );
and ( n12360 , n12358 , n12359 );
buf ( n12361 , n6139 );
xor ( n12362 , n12361 , n12359 );
and ( n12363 , n12362 , n6583 );
or ( n12364 , n12360 , n12363 );
xor ( n12365 , n12261 , n12364 );
buf ( n12366 , n6140 );
xor ( n12367 , n12365 , n12366 );
buf ( n12368 , n6141 );
xor ( n12369 , n12367 , n12368 );
buf ( n12370 , n6142 );
xor ( n12371 , n12369 , n12370 );
xor ( n12372 , n12357 , n12371 );
not ( n12373 , n12372 );
not ( n12374 , n6583 );
buf ( n12375 , n6143 );
and ( n12376 , n12374 , n12375 );
buf ( n12377 , n6144 );
xor ( n12378 , n12377 , n12375 );
and ( n12379 , n12378 , n6583 );
or ( n12380 , n12376 , n12379 );
not ( n12381 , n6583 );
buf ( n12382 , n6145 );
and ( n12383 , n12381 , n12382 );
buf ( n12384 , n6146 );
xor ( n12385 , n12384 , n12382 );
and ( n12386 , n12385 , n6583 );
or ( n12387 , n12383 , n12386 );
xor ( n12388 , n12380 , n12387 );
buf ( n12389 , n6147 );
xor ( n12390 , n12388 , n12389 );
buf ( n12391 , n6148 );
xor ( n12392 , n12390 , n12391 );
xor ( n12393 , n12392 , n10245 );
xor ( n12394 , n11093 , n12393 );
not ( n12395 , n6583 );
buf ( n12396 , n6149 );
and ( n12397 , n12395 , n12396 );
buf ( n12398 , n6150 );
xor ( n12399 , n12398 , n12396 );
and ( n12400 , n12399 , n6583 );
or ( n12401 , n12397 , n12400 );
xor ( n12402 , n11184 , n12401 );
buf ( n12403 , n6151 );
xor ( n12404 , n12402 , n12403 );
buf ( n12405 , n6152 );
xor ( n12406 , n12404 , n12405 );
buf ( n12407 , n6153 );
xor ( n12408 , n12406 , n12407 );
xor ( n12409 , n12394 , n12408 );
and ( n12410 , n12373 , n12409 );
xor ( n12411 , n12349 , n12410 );
buf ( n12412 , n6154 );
not ( n12413 , n6583 );
buf ( n12414 , n6155 );
and ( n12415 , n12413 , n12414 );
buf ( n12416 , n6156 );
xor ( n12417 , n12416 , n12414 );
and ( n12418 , n12417 , n6583 );
or ( n12419 , n12415 , n12418 );
not ( n12420 , n6583 );
buf ( n12421 , n6157 );
and ( n12422 , n12420 , n12421 );
buf ( n12423 , n6158 );
xor ( n12424 , n12423 , n12421 );
and ( n12425 , n12424 , n6583 );
or ( n12426 , n12422 , n12425 );
xor ( n12427 , n12419 , n12426 );
buf ( n12428 , n6159 );
xor ( n12429 , n12427 , n12428 );
buf ( n12430 , n6160 );
xor ( n12431 , n12429 , n12430 );
buf ( n12432 , n6161 );
xor ( n12433 , n12431 , n12432 );
xor ( n12434 , n12412 , n12433 );
not ( n12435 , n6583 );
buf ( n12436 , n6162 );
and ( n12437 , n12435 , n12436 );
buf ( n12438 , n6163 );
xor ( n12439 , n12438 , n12436 );
and ( n12440 , n12439 , n6583 );
or ( n12441 , n12437 , n12440 );
xor ( n12442 , n9672 , n12441 );
xor ( n12443 , n12442 , n8391 );
buf ( n12444 , n6164 );
xor ( n12445 , n12443 , n12444 );
buf ( n12446 , n6165 );
xor ( n12447 , n12445 , n12446 );
xor ( n12448 , n12434 , n12447 );
xor ( n12449 , n11467 , n7980 );
xor ( n12450 , n12449 , n7996 );
not ( n12451 , n12450 );
xor ( n12452 , n10612 , n7654 );
not ( n12453 , n6583 );
buf ( n12454 , n6166 );
and ( n12455 , n12453 , n12454 );
buf ( n12456 , n6167 );
xor ( n12457 , n12456 , n12454 );
and ( n12458 , n12457 , n6583 );
or ( n12459 , n12455 , n12458 );
not ( n12460 , n6583 );
buf ( n12461 , n6168 );
and ( n12462 , n12460 , n12461 );
buf ( n12463 , n6169 );
xor ( n12464 , n12463 , n12461 );
and ( n12465 , n12464 , n6583 );
or ( n12466 , n12462 , n12465 );
xor ( n12467 , n12459 , n12466 );
buf ( n12468 , n6170 );
xor ( n12469 , n12467 , n12468 );
buf ( n12470 , n6171 );
xor ( n12471 , n12469 , n12470 );
buf ( n12472 , n6172 );
xor ( n12473 , n12471 , n12472 );
xor ( n12474 , n12452 , n12473 );
and ( n12475 , n12451 , n12474 );
xor ( n12476 , n12448 , n12475 );
xor ( n12477 , n12411 , n12476 );
not ( n12478 , n6583 );
buf ( n12479 , n6173 );
and ( n12480 , n12478 , n12479 );
buf ( n12481 , n6174 );
xor ( n12482 , n12481 , n12479 );
and ( n12483 , n12482 , n6583 );
or ( n12484 , n12480 , n12483 );
buf ( n12485 , n6175 );
xor ( n12486 , n12484 , n12485 );
buf ( n12487 , n6176 );
xor ( n12488 , n12486 , n12487 );
buf ( n12489 , n6177 );
xor ( n12490 , n12488 , n12489 );
buf ( n12491 , n6178 );
xor ( n12492 , n12490 , n12491 );
xor ( n12493 , n10821 , n12492 );
xor ( n12494 , n12493 , n7632 );
not ( n12495 , n12263 );
and ( n12496 , n12495 , n12293 );
xor ( n12497 , n12494 , n12496 );
xor ( n12498 , n12477 , n12497 );
xor ( n12499 , n11649 , n12152 );
xor ( n12500 , n12499 , n12160 );
not ( n12501 , n6583 );
buf ( n12502 , n6179 );
and ( n12503 , n12501 , n12502 );
buf ( n12504 , n6180 );
xor ( n12505 , n12504 , n12502 );
and ( n12506 , n12505 , n6583 );
or ( n12507 , n12503 , n12506 );
not ( n12508 , n6583 );
buf ( n12509 , n6181 );
and ( n12510 , n12508 , n12509 );
buf ( n12511 , n6182 );
xor ( n12512 , n12511 , n12509 );
and ( n12513 , n12512 , n6583 );
or ( n12514 , n12510 , n12513 );
xor ( n12515 , n12507 , n12514 );
buf ( n12516 , n6183 );
xor ( n12517 , n12515 , n12516 );
buf ( n12518 , n6184 );
xor ( n12519 , n12517 , n12518 );
buf ( n12520 , n6185 );
xor ( n12521 , n12519 , n12520 );
xor ( n12522 , n9817 , n12521 );
xor ( n12523 , n12522 , n10411 );
not ( n12524 , n12523 );
xor ( n12525 , n9914 , n9178 );
xor ( n12526 , n12525 , n9200 );
and ( n12527 , n12524 , n12526 );
xor ( n12528 , n12500 , n12527 );
xor ( n12529 , n12498 , n12528 );
xor ( n12530 , n11346 , n10349 );
xor ( n12531 , n12530 , n7319 );
not ( n12532 , n6583 );
buf ( n12533 , n6186 );
and ( n12534 , n12532 , n12533 );
buf ( n12535 , n6187 );
xor ( n12536 , n12535 , n12533 );
and ( n12537 , n12536 , n6583 );
or ( n12538 , n12534 , n12537 );
not ( n12539 , n6583 );
buf ( n12540 , n6188 );
and ( n12541 , n12539 , n12540 );
buf ( n12542 , n6189 );
xor ( n12543 , n12542 , n12540 );
and ( n12544 , n12543 , n6583 );
or ( n12545 , n12541 , n12544 );
xor ( n12546 , n12538 , n12545 );
buf ( n12547 , n6190 );
xor ( n12548 , n12546 , n12547 );
buf ( n12549 , n6191 );
xor ( n12550 , n12548 , n12549 );
buf ( n12551 , n6192 );
xor ( n12552 , n12550 , n12551 );
xor ( n12553 , n8398 , n12552 );
not ( n12554 , n6583 );
buf ( n12555 , n6193 );
and ( n12556 , n12554 , n12555 );
buf ( n12557 , n6194 );
xor ( n12558 , n12557 , n12555 );
and ( n12559 , n12558 , n6583 );
or ( n12560 , n12556 , n12559 );
not ( n12561 , n6583 );
buf ( n12562 , n6195 );
and ( n12563 , n12561 , n12562 );
buf ( n12564 , n6196 );
xor ( n12565 , n12564 , n12562 );
and ( n12566 , n12565 , n6583 );
or ( n12567 , n12563 , n12566 );
xor ( n12568 , n12560 , n12567 );
xor ( n12569 , n12568 , n8736 );
buf ( n12570 , n6197 );
xor ( n12571 , n12569 , n12570 );
buf ( n12572 , n6198 );
xor ( n12573 , n12571 , n12572 );
xor ( n12574 , n12553 , n12573 );
not ( n12575 , n12574 );
xor ( n12576 , n11598 , n9560 );
xor ( n12577 , n12576 , n8807 );
and ( n12578 , n12575 , n12577 );
xor ( n12579 , n12531 , n12578 );
xor ( n12580 , n12529 , n12579 );
xor ( n12581 , n12326 , n12580 );
not ( n12582 , n6583 );
buf ( n12583 , n6199 );
and ( n12584 , n12582 , n12583 );
buf ( n12585 , n6200 );
xor ( n12586 , n12585 , n12583 );
and ( n12587 , n12586 , n6583 );
or ( n12588 , n12584 , n12587 );
not ( n12589 , n6583 );
buf ( n12590 , n6201 );
and ( n12591 , n12589 , n12590 );
buf ( n12592 , n6202 );
xor ( n12593 , n12592 , n12590 );
and ( n12594 , n12593 , n6583 );
or ( n12595 , n12591 , n12594 );
xor ( n12596 , n12588 , n12595 );
buf ( n12597 , n6203 );
xor ( n12598 , n12596 , n12597 );
buf ( n12599 , n6204 );
xor ( n12600 , n12598 , n12599 );
xor ( n12601 , n12600 , n10515 );
xor ( n12602 , n10275 , n12601 );
not ( n12603 , n6583 );
buf ( n12604 , n6205 );
and ( n12605 , n12603 , n12604 );
buf ( n12606 , n6206 );
xor ( n12607 , n12606 , n12604 );
and ( n12608 , n12607 , n6583 );
or ( n12609 , n12605 , n12608 );
not ( n12610 , n6583 );
buf ( n12611 , n6207 );
and ( n12612 , n12610 , n12611 );
buf ( n12613 , n6208 );
xor ( n12614 , n12613 , n12611 );
and ( n12615 , n12614 , n6583 );
or ( n12616 , n12612 , n12615 );
xor ( n12617 , n12609 , n12616 );
buf ( n12618 , n6209 );
xor ( n12619 , n12617 , n12618 );
xor ( n12620 , n12619 , n12194 );
buf ( n12621 , n6210 );
xor ( n12622 , n12620 , n12621 );
xor ( n12623 , n12602 , n12622 );
xor ( n12624 , n9379 , n11100 );
xor ( n12625 , n12624 , n10893 );
not ( n12626 , n12625 );
not ( n12627 , n6583 );
buf ( n12628 , n6211 );
and ( n12629 , n12627 , n12628 );
buf ( n12630 , n6212 );
xor ( n12631 , n12630 , n12628 );
and ( n12632 , n12631 , n6583 );
or ( n12633 , n12629 , n12632 );
not ( n12634 , n6583 );
buf ( n12635 , n6213 );
and ( n12636 , n12634 , n12635 );
buf ( n12637 , n6214 );
xor ( n12638 , n12637 , n12635 );
and ( n12639 , n12638 , n6583 );
or ( n12640 , n12636 , n12639 );
xor ( n12641 , n12633 , n12640 );
buf ( n12642 , n6215 );
xor ( n12643 , n12641 , n12642 );
buf ( n12644 , n6216 );
xor ( n12645 , n12643 , n12644 );
buf ( n12646 , n6217 );
xor ( n12647 , n12645 , n12646 );
xor ( n12648 , n11215 , n12647 );
not ( n12649 , n6583 );
buf ( n12650 , n6218 );
and ( n12651 , n12649 , n12650 );
buf ( n12652 , n6219 );
xor ( n12653 , n12652 , n12650 );
and ( n12654 , n12653 , n6583 );
or ( n12655 , n12651 , n12654 );
buf ( n12656 , n6220 );
xor ( n12657 , n12655 , n12656 );
xor ( n12658 , n12657 , n11718 );
buf ( n12659 , n6221 );
xor ( n12660 , n12658 , n12659 );
buf ( n12661 , n6222 );
xor ( n12662 , n12660 , n12661 );
xor ( n12663 , n12648 , n12662 );
and ( n12664 , n12626 , n12663 );
xor ( n12665 , n12623 , n12664 );
buf ( n12666 , n6223 );
xor ( n12667 , n12666 , n7710 );
xor ( n12668 , n12667 , n6705 );
xor ( n12669 , n11309 , n7335 );
xor ( n12670 , n12669 , n10098 );
not ( n12671 , n12670 );
xor ( n12672 , n10549 , n10915 );
xor ( n12673 , n12672 , n10142 );
and ( n12674 , n12671 , n12673 );
xor ( n12675 , n12668 , n12674 );
xor ( n12676 , n12665 , n12675 );
not ( n12677 , n6583 );
buf ( n12678 , n6224 );
and ( n12679 , n12677 , n12678 );
buf ( n12680 , n6225 );
xor ( n12681 , n12680 , n12678 );
and ( n12682 , n12681 , n6583 );
or ( n12683 , n12679 , n12682 );
not ( n12684 , n6583 );
buf ( n12685 , n6226 );
and ( n12686 , n12684 , n12685 );
buf ( n12687 , n6227 );
xor ( n12688 , n12687 , n12685 );
and ( n12689 , n12688 , n6583 );
or ( n12690 , n12686 , n12689 );
xor ( n12691 , n12690 , n10450 );
buf ( n12692 , n6228 );
xor ( n12693 , n12691 , n12692 );
xor ( n12694 , n12693 , n9991 );
buf ( n12695 , n6229 );
xor ( n12696 , n12694 , n12695 );
xor ( n12697 , n12683 , n12696 );
xor ( n12698 , n12697 , n9478 );
xor ( n12699 , n6747 , n9809 );
xor ( n12700 , n12699 , n9825 );
not ( n12701 , n12700 );
not ( n12702 , n6583 );
buf ( n12703 , n6230 );
and ( n12704 , n12702 , n12703 );
buf ( n12705 , n6231 );
xor ( n12706 , n12705 , n12703 );
and ( n12707 , n12706 , n6583 );
or ( n12708 , n12704 , n12707 );
not ( n12709 , n6583 );
buf ( n12710 , n6232 );
and ( n12711 , n12709 , n12710 );
buf ( n12712 , n6233 );
xor ( n12713 , n12712 , n12710 );
and ( n12714 , n12713 , n6583 );
or ( n12715 , n12711 , n12714 );
xor ( n12716 , n12708 , n12715 );
xor ( n12717 , n12716 , n11606 );
buf ( n12718 , n6234 );
xor ( n12719 , n12717 , n12718 );
buf ( n12720 , n6235 );
xor ( n12721 , n12719 , n12720 );
xor ( n12722 , n8502 , n12721 );
xor ( n12723 , n12722 , n11805 );
and ( n12724 , n12701 , n12723 );
xor ( n12725 , n12698 , n12724 );
xor ( n12726 , n12676 , n12725 );
not ( n12727 , n6583 );
buf ( n12728 , n6236 );
and ( n12729 , n12727 , n12728 );
buf ( n12730 , n6237 );
xor ( n12731 , n12730 , n12728 );
and ( n12732 , n12731 , n6583 );
or ( n12733 , n12729 , n12732 );
xor ( n12734 , n12733 , n8083 );
xor ( n12735 , n12734 , n8105 );
xor ( n12736 , n9528 , n11386 );
not ( n12737 , n6583 );
buf ( n12738 , n6238 );
and ( n12739 , n12737 , n12738 );
buf ( n12740 , n6239 );
xor ( n12741 , n12740 , n12738 );
and ( n12742 , n12741 , n6583 );
or ( n12743 , n12739 , n12742 );
not ( n12744 , n6583 );
buf ( n12745 , n6240 );
and ( n12746 , n12744 , n12745 );
buf ( n12747 , n6241 );
xor ( n12748 , n12747 , n12745 );
and ( n12749 , n12748 , n6583 );
or ( n12750 , n12746 , n12749 );
xor ( n12751 , n12743 , n12750 );
xor ( n12752 , n12751 , n9025 );
buf ( n12753 , n6242 );
xor ( n12754 , n12752 , n12753 );
buf ( n12755 , n6243 );
xor ( n12756 , n12754 , n12755 );
xor ( n12757 , n12736 , n12756 );
not ( n12758 , n12757 );
xor ( n12759 , n9657 , n8167 );
xor ( n12760 , n12759 , n8189 );
and ( n12761 , n12758 , n12760 );
xor ( n12762 , n12735 , n12761 );
xor ( n12763 , n12726 , n12762 );
xor ( n12764 , n11643 , n12152 );
xor ( n12765 , n12764 , n12160 );
xor ( n12766 , n8265 , n9244 );
xor ( n12767 , n12766 , n10166 );
not ( n12768 , n12767 );
not ( n12769 , n6583 );
buf ( n12770 , n6244 );
and ( n12771 , n12769 , n12770 );
buf ( n12772 , n6245 );
xor ( n12773 , n12772 , n12770 );
and ( n12774 , n12773 , n6583 );
or ( n12775 , n12771 , n12774 );
buf ( n12776 , n6246 );
xor ( n12777 , n12775 , n12776 );
buf ( n12778 , n6247 );
xor ( n12779 , n12777 , n12778 );
xor ( n12780 , n12779 , n9678 );
buf ( n12781 , n6248 );
xor ( n12782 , n12780 , n12781 );
xor ( n12783 , n9304 , n12782 );
xor ( n12784 , n12783 , n8369 );
and ( n12785 , n12768 , n12784 );
xor ( n12786 , n12765 , n12785 );
xor ( n12787 , n12763 , n12786 );
xor ( n12788 , n12581 , n12787 );
xor ( n12789 , n7209 , n8036 );
xor ( n12790 , n12789 , n8058 );
xor ( n12791 , n10939 , n10797 );
not ( n12792 , n6583 );
buf ( n12793 , n6249 );
and ( n12794 , n12792 , n12793 );
buf ( n12795 , n6250 );
xor ( n12796 , n12795 , n12793 );
and ( n12797 , n12796 , n6583 );
or ( n12798 , n12794 , n12797 );
xor ( n12799 , n12798 , n11358 );
buf ( n12800 , n6251 );
xor ( n12801 , n12799 , n12800 );
xor ( n12802 , n12801 , n8865 );
buf ( n12803 , n6252 );
xor ( n12804 , n12802 , n12803 );
xor ( n12805 , n12791 , n12804 );
not ( n12806 , n12805 );
xor ( n12807 , n6868 , n8822 );
xor ( n12808 , n12807 , n11050 );
and ( n12809 , n12806 , n12808 );
xor ( n12810 , n12790 , n12809 );
xor ( n12811 , n9293 , n12782 );
xor ( n12812 , n12811 , n8369 );
not ( n12813 , n6583 );
buf ( n12814 , n6253 );
and ( n12815 , n12813 , n12814 );
buf ( n12816 , n6254 );
xor ( n12817 , n12816 , n12814 );
and ( n12818 , n12817 , n6583 );
or ( n12819 , n12815 , n12818 );
xor ( n12820 , n12819 , n6705 );
xor ( n12821 , n12820 , n6727 );
not ( n12822 , n12821 );
xor ( n12823 , n11973 , n11684 );
xor ( n12824 , n12823 , n11218 );
and ( n12825 , n12822 , n12824 );
xor ( n12826 , n12812 , n12825 );
not ( n12827 , n6583 );
buf ( n12828 , n6255 );
and ( n12829 , n12827 , n12828 );
buf ( n12830 , n6256 );
xor ( n12831 , n12830 , n12828 );
and ( n12832 , n12831 , n6583 );
or ( n12833 , n12829 , n12832 );
xor ( n12834 , n12833 , n12270 );
buf ( n12835 , n6257 );
xor ( n12836 , n12834 , n12835 );
buf ( n12837 , n6258 );
xor ( n12838 , n12836 , n12837 );
buf ( n12839 , n6259 );
xor ( n12840 , n12838 , n12839 );
xor ( n12841 , n10106 , n12840 );
not ( n12842 , n6583 );
buf ( n12843 , n6260 );
and ( n12844 , n12842 , n12843 );
buf ( n12845 , n6261 );
xor ( n12846 , n12845 , n12843 );
and ( n12847 , n12846 , n6583 );
or ( n12848 , n12844 , n12847 );
buf ( n12849 , n6262 );
xor ( n12850 , n12848 , n12849 );
buf ( n12851 , n6263 );
xor ( n12852 , n12850 , n12851 );
buf ( n12853 , n6264 );
xor ( n12854 , n12852 , n12853 );
buf ( n12855 , n6265 );
xor ( n12856 , n12854 , n12855 );
xor ( n12857 , n12841 , n12856 );
buf ( n12858 , n6266 );
xor ( n12859 , n12858 , n12447 );
not ( n12860 , n6583 );
buf ( n12861 , n6267 );
and ( n12862 , n12860 , n12861 );
buf ( n12863 , n6268 );
xor ( n12864 , n12863 , n12861 );
and ( n12865 , n12864 , n6583 );
or ( n12866 , n12862 , n12865 );
xor ( n12867 , n12866 , n10651 );
buf ( n12868 , n6269 );
xor ( n12869 , n12867 , n12868 );
buf ( n12870 , n6270 );
xor ( n12871 , n12869 , n12870 );
buf ( n12872 , n6271 );
xor ( n12873 , n12871 , n12872 );
xor ( n12874 , n12859 , n12873 );
not ( n12875 , n12874 );
xor ( n12876 , n12597 , n10530 );
xor ( n12877 , n12876 , n10552 );
and ( n12878 , n12875 , n12877 );
xor ( n12879 , n12857 , n12878 );
xor ( n12880 , n12826 , n12879 );
xor ( n12881 , n8355 , n9362 );
xor ( n12882 , n12881 , n9384 );
xor ( n12883 , n8545 , n9406 );
xor ( n12884 , n12883 , n9428 );
not ( n12885 , n12884 );
xor ( n12886 , n11287 , n7319 );
xor ( n12887 , n12886 , n7335 );
and ( n12888 , n12885 , n12887 );
xor ( n12889 , n12882 , n12888 );
xor ( n12890 , n12880 , n12889 );
xor ( n12891 , n7181 , n12015 );
xor ( n12892 , n12891 , n12037 );
not ( n12893 , n12790 );
and ( n12894 , n12893 , n12805 );
xor ( n12895 , n12892 , n12894 );
xor ( n12896 , n12890 , n12895 );
not ( n12897 , n6583 );
buf ( n12898 , n6272 );
and ( n12899 , n12897 , n12898 );
buf ( n12900 , n6273 );
xor ( n12901 , n12900 , n12898 );
and ( n12902 , n12901 , n6583 );
or ( n12903 , n12899 , n12902 );
not ( n12904 , n6583 );
buf ( n12905 , n6274 );
and ( n12906 , n12904 , n12905 );
buf ( n12907 , n6275 );
xor ( n12908 , n12907 , n12905 );
and ( n12909 , n12908 , n6583 );
or ( n12910 , n12906 , n12909 );
xor ( n12911 , n12903 , n12910 );
xor ( n12912 , n12911 , n11950 );
buf ( n12913 , n6276 );
xor ( n12914 , n12912 , n12913 );
xor ( n12915 , n12914 , n8996 );
xor ( n12916 , n6933 , n12915 );
xor ( n12917 , n12916 , n9285 );
not ( n12918 , n6583 );
buf ( n12919 , n6277 );
and ( n12920 , n12918 , n12919 );
buf ( n12921 , n6278 );
xor ( n12922 , n12921 , n12919 );
and ( n12923 , n12922 , n6583 );
or ( n12924 , n12920 , n12923 );
xor ( n12925 , n12924 , n10563 );
buf ( n12926 , n6279 );
xor ( n12927 , n12925 , n12926 );
buf ( n12928 , n6280 );
xor ( n12929 , n12927 , n12928 );
buf ( n12930 , n6281 );
xor ( n12931 , n12929 , n12930 );
xor ( n12932 , n7487 , n12931 );
xor ( n12933 , n12932 , n9615 );
not ( n12934 , n12933 );
buf ( n12935 , n6282 );
xor ( n12936 , n12935 , n8189 );
xor ( n12937 , n12936 , n10822 );
and ( n12938 , n12934 , n12937 );
xor ( n12939 , n12917 , n12938 );
xor ( n12940 , n12896 , n12939 );
xor ( n12941 , n12810 , n12940 );
not ( n12942 , n6583 );
buf ( n12943 , n6283 );
and ( n12944 , n12942 , n12943 );
buf ( n12945 , n6284 );
xor ( n12946 , n12945 , n12943 );
and ( n12947 , n12946 , n6583 );
or ( n12948 , n12944 , n12947 );
xor ( n12949 , n12948 , n12819 );
xor ( n12950 , n12949 , n6684 );
buf ( n12951 , n6285 );
xor ( n12952 , n12950 , n12951 );
buf ( n12953 , n6286 );
xor ( n12954 , n12952 , n12953 );
xor ( n12955 , n12642 , n12954 );
xor ( n12956 , n12955 , n11739 );
not ( n12957 , n6583 );
buf ( n12958 , n6287 );
and ( n12959 , n12957 , n12958 );
buf ( n12960 , n6288 );
xor ( n12961 , n12960 , n12958 );
and ( n12962 , n12961 , n6583 );
or ( n12963 , n12959 , n12962 );
not ( n12964 , n6583 );
buf ( n12965 , n6289 );
and ( n12966 , n12964 , n12965 );
buf ( n12967 , n6290 );
xor ( n12968 , n12967 , n12965 );
and ( n12969 , n12968 , n6583 );
or ( n12970 , n12966 , n12969 );
xor ( n12971 , n12963 , n12970 );
buf ( n12972 , n6291 );
xor ( n12973 , n12971 , n12972 );
buf ( n12974 , n6292 );
buf ( n12975 , n12974 );
xor ( n12976 , n12973 , n12975 );
buf ( n12977 , n6293 );
xor ( n12978 , n12976 , n12977 );
xor ( n12979 , n8457 , n12978 );
xor ( n12980 , n12979 , n11325 );
not ( n12981 , n12980 );
xor ( n12982 , n12159 , n7428 );
xor ( n12983 , n12982 , n7579 );
and ( n12984 , n12981 , n12983 );
xor ( n12985 , n12956 , n12984 );
not ( n12986 , n6583 );
buf ( n12987 , n6294 );
and ( n12988 , n12986 , n12987 );
buf ( n12989 , n6295 );
xor ( n12990 , n12989 , n12987 );
and ( n12991 , n12990 , n6583 );
or ( n12992 , n12988 , n12991 );
buf ( n12993 , n6296 );
xor ( n12994 , n12992 , n12993 );
buf ( n12995 , n6297 );
xor ( n12996 , n12994 , n12995 );
xor ( n12997 , n12996 , n8768 );
buf ( n12998 , n6298 );
xor ( n12999 , n12997 , n12998 );
xor ( n13000 , n10910 , n12999 );
not ( n13001 , n6583 );
buf ( n13002 , n6299 );
and ( n13003 , n13001 , n13002 );
buf ( n13004 , n6300 );
xor ( n13005 , n13004 , n13002 );
and ( n13006 , n13005 , n6583 );
or ( n13007 , n13003 , n13006 );
not ( n13008 , n6583 );
buf ( n13009 , n6301 );
and ( n13010 , n13008 , n13009 );
buf ( n13011 , n6302 );
xor ( n13012 , n13011 , n13009 );
and ( n13013 , n13012 , n6583 );
or ( n13014 , n13010 , n13013 );
xor ( n13015 , n13007 , n13014 );
xor ( n13016 , n13015 , n8509 );
buf ( n13017 , n6303 );
xor ( n13018 , n13016 , n13017 );
buf ( n13019 , n6304 );
xor ( n13020 , n13018 , n13019 );
xor ( n13021 , n13000 , n13020 );
xor ( n13022 , n10472 , n11761 );
xor ( n13023 , n13022 , n12308 );
not ( n13024 , n13023 );
xor ( n13025 , n6946 , n12915 );
xor ( n13026 , n13025 , n9285 );
and ( n13027 , n13024 , n13026 );
xor ( n13028 , n13021 , n13027 );
xor ( n13029 , n12985 , n13028 );
xor ( n13030 , n11525 , n7173 );
xor ( n13031 , n13030 , n7189 );
xor ( n13032 , n11558 , n10776 );
xor ( n13033 , n13032 , n10797 );
not ( n13034 , n13033 );
buf ( n13035 , n6305 );
buf ( n13036 , n6306 );
xor ( n13037 , n9834 , n13036 );
buf ( n13038 , n6307 );
xor ( n13039 , n13037 , n13038 );
buf ( n13040 , n6308 );
xor ( n13041 , n13039 , n13040 );
xor ( n13042 , n13041 , n11223 );
xor ( n13043 , n13035 , n13042 );
xor ( n13044 , n13043 , n12552 );
and ( n13045 , n13034 , n13044 );
xor ( n13046 , n13031 , n13045 );
xor ( n13047 , n13029 , n13046 );
xor ( n13048 , n8881 , n7908 );
xor ( n13049 , n13048 , n9069 );
not ( n13050 , n6583 );
buf ( n13051 , n6309 );
and ( n13052 , n13050 , n13051 );
buf ( n13053 , n6310 );
xor ( n13054 , n13053 , n13051 );
and ( n13055 , n13054 , n6583 );
or ( n13056 , n13052 , n13055 );
not ( n13057 , n6583 );
buf ( n13058 , n6311 );
and ( n13059 , n13057 , n13058 );
buf ( n13060 , n6312 );
xor ( n13061 , n13060 , n13058 );
and ( n13062 , n13061 , n6583 );
or ( n13063 , n13059 , n13062 );
xor ( n13064 , n13056 , n13063 );
xor ( n13065 , n13064 , n11686 );
xor ( n13066 , n13065 , n7558 );
buf ( n13067 , n6313 );
xor ( n13068 , n13066 , n13067 );
xor ( n13069 , n7387 , n13068 );
not ( n13070 , n6583 );
buf ( n13071 , n6314 );
and ( n13072 , n13070 , n13071 );
buf ( n13073 , n6315 );
xor ( n13074 , n13073 , n13071 );
and ( n13075 , n13074 , n6583 );
or ( n13076 , n13072 , n13075 );
not ( n13077 , n6583 );
buf ( n13078 , n6316 );
and ( n13079 , n13077 , n13078 );
buf ( n13080 , n6317 );
xor ( n13081 , n13080 , n13078 );
and ( n13082 , n13081 , n6583 );
or ( n13083 , n13079 , n13082 );
xor ( n13084 , n13076 , n13083 );
buf ( n13085 , n6318 );
xor ( n13086 , n13084 , n13085 );
xor ( n13087 , n13086 , n8637 );
buf ( n13088 , n6319 );
xor ( n13089 , n13087 , n13088 );
xor ( n13090 , n13069 , n13089 );
not ( n13091 , n13090 );
not ( n13092 , n6583 );
buf ( n13093 , n6320 );
and ( n13094 , n13092 , n13093 );
buf ( n13095 , n6321 );
xor ( n13096 , n13095 , n13093 );
and ( n13097 , n13096 , n6583 );
or ( n13098 , n13094 , n13097 );
xor ( n13099 , n8563 , n13098 );
buf ( n13100 , n6322 );
xor ( n13101 , n13099 , n13100 );
buf ( n13102 , n6323 );
xor ( n13103 , n13101 , n13102 );
xor ( n13104 , n13103 , n8730 );
xor ( n13105 , n10866 , n13104 );
xor ( n13106 , n13105 , n9178 );
and ( n13107 , n13091 , n13106 );
xor ( n13108 , n13049 , n13107 );
xor ( n13109 , n13047 , n13108 );
xor ( n13110 , n12487 , n8635 );
xor ( n13111 , n13110 , n8705 );
buf ( n13112 , n6324 );
xor ( n13113 , n13112 , n10619 );
xor ( n13114 , n13113 , n11684 );
not ( n13115 , n13114 );
xor ( n13116 , n10281 , n12601 );
xor ( n13117 , n13116 , n12622 );
and ( n13118 , n13115 , n13117 );
xor ( n13119 , n13111 , n13118 );
xor ( n13120 , n13109 , n13119 );
xor ( n13121 , n12941 , n13120 );
not ( n13122 , n13121 );
xor ( n13123 , n11861 , n7494 );
xor ( n13124 , n13123 , n7516 );
xor ( n13125 , n9736 , n7469 );
xor ( n13126 , n13125 , n11147 );
not ( n13127 , n13126 );
buf ( n13128 , n6325 );
not ( n13129 , n6583 );
buf ( n13130 , n6326 );
and ( n13131 , n13129 , n13130 );
buf ( n13132 , n6327 );
xor ( n13133 , n13132 , n13130 );
and ( n13134 , n13133 , n6583 );
or ( n13135 , n13131 , n13134 );
not ( n13136 , n6583 );
buf ( n13137 , n6328 );
and ( n13138 , n13136 , n13137 );
buf ( n13139 , n6329 );
xor ( n13140 , n13139 , n13137 );
and ( n13141 , n13140 , n6583 );
or ( n13142 , n13138 , n13141 );
xor ( n13143 , n13135 , n13142 );
buf ( n13144 , n6330 );
xor ( n13145 , n13143 , n13144 );
buf ( n13146 , n6331 );
xor ( n13147 , n13145 , n13146 );
buf ( n13148 , n6332 );
xor ( n13149 , n13147 , n13148 );
xor ( n13150 , n13128 , n13149 );
not ( n13151 , n6583 );
buf ( n13152 , n6333 );
and ( n13153 , n13151 , n13152 );
buf ( n13154 , n6334 );
xor ( n13155 , n13154 , n13152 );
and ( n13156 , n13155 , n6583 );
or ( n13157 , n13153 , n13156 );
not ( n13158 , n6583 );
and ( n13159 , n13158 , n12253 );
buf ( n13160 , n6335 );
xor ( n13161 , n13160 , n12253 );
and ( n13162 , n13161 , n6583 );
or ( n13163 , n13159 , n13162 );
xor ( n13164 , n13157 , n13163 );
buf ( n13165 , n6336 );
xor ( n13166 , n13164 , n13165 );
buf ( n13167 , n6337 );
xor ( n13168 , n13166 , n13167 );
xor ( n13169 , n13168 , n12412 );
xor ( n13170 , n13150 , n13169 );
and ( n13171 , n13127 , n13170 );
xor ( n13172 , n13124 , n13171 );
xor ( n13173 , n8098 , n8318 );
xor ( n13174 , n13173 , n8340 );
xor ( n13175 , n9937 , n9200 );
not ( n13176 , n6583 );
buf ( n13177 , n6338 );
and ( n13178 , n13176 , n13177 );
buf ( n13179 , n6339 );
xor ( n13180 , n13179 , n13177 );
and ( n13181 , n13180 , n6583 );
or ( n13182 , n13178 , n13181 );
xor ( n13183 , n13182 , n11193 );
xor ( n13184 , n13183 , n7656 );
buf ( n13185 , n6340 );
xor ( n13186 , n13184 , n13185 );
buf ( n13187 , n6341 );
xor ( n13188 , n13186 , n13187 );
xor ( n13189 , n13175 , n13188 );
not ( n13190 , n13189 );
buf ( n13191 , n6342 );
xor ( n13192 , n13191 , n7238 );
xor ( n13193 , n13192 , n7533 );
and ( n13194 , n13190 , n13193 );
xor ( n13195 , n13174 , n13194 );
xor ( n13196 , n8029 , n12347 );
xor ( n13197 , n13196 , n9639 );
buf ( n13198 , n6343 );
xor ( n13199 , n13198 , n13042 );
xor ( n13200 , n13199 , n12552 );
not ( n13201 , n13200 );
xor ( n13202 , n9226 , n10971 );
xor ( n13203 , n13202 , n6947 );
and ( n13204 , n13201 , n13203 );
xor ( n13205 , n13197 , n13204 );
xor ( n13206 , n13195 , n13205 );
xor ( n13207 , n12970 , n10673 );
xor ( n13208 , n13207 , n10327 );
xor ( n13209 , n7142 , n10603 );
xor ( n13210 , n13209 , n10619 );
not ( n13211 , n13210 );
not ( n13212 , n6583 );
buf ( n13213 , n6344 );
and ( n13214 , n13212 , n13213 );
buf ( n13215 , n6345 );
xor ( n13216 , n13215 , n13213 );
and ( n13217 , n13216 , n6583 );
or ( n13218 , n13214 , n13217 );
xor ( n13219 , n11007 , n13218 );
buf ( n13220 , n6346 );
xor ( n13221 , n13219 , n13220 );
buf ( n13222 , n6347 );
xor ( n13223 , n13221 , n13222 );
buf ( n13224 , n6348 );
xor ( n13225 , n13223 , n13224 );
xor ( n13226 , n8247 , n13225 );
not ( n13227 , n6583 );
buf ( n13228 , n6349 );
and ( n13229 , n13227 , n13228 );
buf ( n13230 , n6350 );
xor ( n13231 , n13230 , n13228 );
and ( n13232 , n13231 , n6583 );
or ( n13233 , n13229 , n13232 );
not ( n13234 , n6583 );
buf ( n13235 , n6351 );
and ( n13236 , n13234 , n13235 );
buf ( n13237 , n6352 );
xor ( n13238 , n13237 , n13235 );
and ( n13239 , n13238 , n6583 );
or ( n13240 , n13236 , n13239 );
xor ( n13241 , n13233 , n13240 );
buf ( n13242 , n6353 );
xor ( n13243 , n13241 , n13242 );
xor ( n13244 , n13243 , n10351 );
buf ( n13245 , n6354 );
xor ( n13246 , n13244 , n13245 );
xor ( n13247 , n13226 , n13246 );
and ( n13248 , n13211 , n13247 );
xor ( n13249 , n13208 , n13248 );
xor ( n13250 , n13206 , n13249 );
not ( n13251 , n6583 );
buf ( n13252 , n6355 );
and ( n13253 , n13251 , n13252 );
buf ( n13254 , n6356 );
xor ( n13255 , n13254 , n13252 );
and ( n13256 , n13255 , n6583 );
or ( n13257 , n13253 , n13256 );
xor ( n13258 , n13257 , n7029 );
xor ( n13259 , n13258 , n7051 );
xor ( n13260 , n10383 , n11314 );
xor ( n13261 , n13260 , n11497 );
not ( n13262 , n13261 );
xor ( n13263 , n11624 , n6896 );
xor ( n13264 , n13263 , n6918 );
and ( n13265 , n13262 , n13264 );
xor ( n13266 , n13259 , n13265 );
xor ( n13267 , n13250 , n13266 );
xor ( n13268 , n9421 , n8863 );
not ( n13269 , n6583 );
buf ( n13270 , n6357 );
and ( n13271 , n13269 , n13270 );
buf ( n13272 , n6358 );
xor ( n13273 , n13272 , n13270 );
and ( n13274 , n13273 , n6583 );
or ( n13275 , n13271 , n13274 );
xor ( n13276 , n13275 , n11829 );
buf ( n13277 , n6359 );
xor ( n13278 , n13276 , n13277 );
buf ( n13279 , n6360 );
xor ( n13280 , n13278 , n13279 );
buf ( n13281 , n6361 );
xor ( n13282 , n13280 , n13281 );
xor ( n13283 , n13268 , n13282 );
not ( n13284 , n13124 );
and ( n13285 , n13284 , n13126 );
xor ( n13286 , n13283 , n13285 );
xor ( n13287 , n13267 , n13286 );
xor ( n13288 , n13172 , n13287 );
buf ( n13289 , n6362 );
xor ( n13290 , n13289 , n9660 );
not ( n13291 , n6583 );
buf ( n13292 , n6363 );
and ( n13293 , n13291 , n13292 );
buf ( n13294 , n6364 );
xor ( n13295 , n13294 , n13292 );
and ( n13296 , n13295 , n6583 );
or ( n13297 , n13293 , n13296 );
buf ( n13298 , n6365 );
xor ( n13299 , n13297 , n13298 );
xor ( n13300 , n13299 , n12935 );
buf ( n13301 , n6366 );
xor ( n13302 , n13300 , n13301 );
buf ( n13303 , n6367 );
xor ( n13304 , n13302 , n13303 );
xor ( n13305 , n13290 , n13304 );
xor ( n13306 , n8504 , n12721 );
xor ( n13307 , n13306 , n11805 );
not ( n13308 , n13307 );
xor ( n13309 , n11058 , n9262 );
not ( n13310 , n6583 );
buf ( n13311 , n6368 );
and ( n13312 , n13310 , n13311 );
buf ( n13313 , n6369 );
xor ( n13314 , n13313 , n13311 );
and ( n13315 , n13314 , n6583 );
or ( n13316 , n13312 , n13315 );
not ( n13317 , n6583 );
buf ( n13318 , n6370 );
and ( n13319 , n13317 , n13318 );
buf ( n13320 , n6371 );
xor ( n13321 , n13320 , n13318 );
and ( n13322 , n13321 , n6583 );
or ( n13323 , n13319 , n13322 );
xor ( n13324 , n13316 , n13323 );
buf ( n13325 , n6372 );
xor ( n13326 , n13324 , n13325 );
buf ( n13327 , n6373 );
xor ( n13328 , n13326 , n13327 );
xor ( n13329 , n13328 , n13128 );
xor ( n13330 , n13309 , n13329 );
and ( n13331 , n13308 , n13330 );
xor ( n13332 , n13305 , n13331 );
xor ( n13333 , n12913 , n6636 );
xor ( n13334 , n13333 , n9018 );
xor ( n13335 , n12151 , n7406 );
xor ( n13336 , n13335 , n7428 );
not ( n13337 , n13336 );
xor ( n13338 , n11725 , n6727 );
xor ( n13339 , n13338 , n12213 );
and ( n13340 , n13337 , n13339 );
xor ( n13341 , n13334 , n13340 );
xor ( n13342 , n13332 , n13341 );
xor ( n13343 , n10363 , n11292 );
xor ( n13344 , n13343 , n11314 );
not ( n13345 , n6583 );
buf ( n13346 , n6374 );
and ( n13347 , n13345 , n13346 );
buf ( n13348 , n6375 );
xor ( n13349 , n13348 , n13346 );
and ( n13350 , n13349 , n6583 );
or ( n13351 , n13347 , n13350 );
buf ( n13352 , n6376 );
xor ( n13353 , n13351 , n13352 );
xor ( n13354 , n13353 , n8953 );
buf ( n13355 , n6377 );
xor ( n13356 , n13354 , n13355 );
buf ( n13357 , n6378 );
xor ( n13358 , n13356 , n13357 );
xor ( n13359 , n7072 , n13358 );
not ( n13360 , n6583 );
buf ( n13361 , n6379 );
and ( n13362 , n13360 , n13361 );
buf ( n13363 , n6380 );
xor ( n13364 , n13363 , n13361 );
and ( n13365 , n13364 , n6583 );
or ( n13366 , n13362 , n13365 );
not ( n13367 , n6583 );
buf ( n13368 , n6381 );
and ( n13369 , n13367 , n13368 );
buf ( n13370 , n6382 );
xor ( n13371 , n13370 , n13368 );
and ( n13372 , n13371 , n6583 );
or ( n13373 , n13369 , n13372 );
xor ( n13374 , n13366 , n13373 );
buf ( n13375 , n6383 );
xor ( n13376 , n13374 , n13375 );
xor ( n13377 , n13376 , n9203 );
xor ( n13378 , n13377 , n7195 );
xor ( n13379 , n13359 , n13378 );
not ( n13380 , n13379 );
xor ( n13381 , n13316 , n13149 );
xor ( n13382 , n13381 , n13169 );
and ( n13383 , n13380 , n13382 );
xor ( n13384 , n13344 , n13383 );
xor ( n13385 , n13342 , n13384 );
buf ( n13386 , n6384 );
xor ( n13387 , n13386 , n7267 );
xor ( n13388 , n13387 , n7289 );
xor ( n13389 , n10775 , n10219 );
xor ( n13390 , n13389 , n9715 );
not ( n13391 , n13390 );
xor ( n13392 , n11986 , n11218 );
xor ( n13393 , n13392 , n7782 );
and ( n13394 , n13391 , n13393 );
xor ( n13395 , n13388 , n13394 );
xor ( n13396 , n13385 , n13395 );
xor ( n13397 , n9917 , n9178 );
xor ( n13398 , n13397 , n9200 );
not ( n13399 , n6583 );
buf ( n13400 , n6385 );
and ( n13401 , n13399 , n13400 );
buf ( n13402 , n6386 );
xor ( n13403 , n13402 , n13400 );
and ( n13404 , n13403 , n6583 );
or ( n13405 , n13401 , n13404 );
not ( n13406 , n6583 );
buf ( n13407 , n6387 );
and ( n13408 , n13406 , n13407 );
buf ( n13409 , n6388 );
xor ( n13410 , n13409 , n13407 );
and ( n13411 , n13410 , n6583 );
or ( n13412 , n13408 , n13411 );
xor ( n13413 , n13405 , n13412 );
xor ( n13414 , n13413 , n13198 );
buf ( n13415 , n6389 );
xor ( n13416 , n13414 , n13415 );
xor ( n13417 , n13416 , n13035 );
xor ( n13418 , n12432 , n13417 );
xor ( n13419 , n13418 , n8412 );
not ( n13420 , n13419 );
xor ( n13421 , n6857 , n8822 );
xor ( n13422 , n13421 , n11050 );
and ( n13423 , n13420 , n13422 );
xor ( n13424 , n13398 , n13423 );
xor ( n13425 , n13396 , n13424 );
xor ( n13426 , n13288 , n13425 );
and ( n13427 , n13122 , n13426 );
xor ( n13428 , n12788 , n13427 );
and ( n13429 , n13428 , n6584 );
or ( n13430 , n12254 , n13429 );
and ( n13431 , n12251 , n13430 );
buf ( n13432 , n13431 );
buf ( n13433 , n13432 );
not ( n13434 , n6578 );
not ( n13435 , n6584 );
and ( n13436 , n13435 , n9621 );
xor ( n13437 , n9626 , n8992 );
xor ( n13438 , n13437 , n8167 );
not ( n13439 , n6583 );
buf ( n13440 , n6390 );
and ( n13441 , n13439 , n13440 );
buf ( n13442 , n6391 );
xor ( n13443 , n13442 , n13440 );
and ( n13444 , n13443 , n6583 );
or ( n13445 , n13441 , n13444 );
xor ( n13446 , n13445 , n11072 );
not ( n13447 , n6583 );
buf ( n13448 , n6392 );
and ( n13449 , n13447 , n13448 );
buf ( n13450 , n6393 );
xor ( n13451 , n13450 , n13448 );
and ( n13452 , n13451 , n6583 );
or ( n13453 , n13449 , n13452 );
not ( n13454 , n6583 );
buf ( n13455 , n6394 );
and ( n13456 , n13454 , n13455 );
buf ( n13457 , n6395 );
xor ( n13458 , n13457 , n13455 );
and ( n13459 , n13458 , n6583 );
or ( n13460 , n13456 , n13459 );
xor ( n13461 , n13453 , n13460 );
buf ( n13462 , n6396 );
xor ( n13463 , n13461 , n13462 );
buf ( n13464 , n6397 );
xor ( n13465 , n13463 , n13464 );
buf ( n13466 , n6398 );
xor ( n13467 , n13465 , n13466 );
xor ( n13468 , n13446 , n13467 );
not ( n13469 , n13468 );
xor ( n13470 , n7385 , n13068 );
xor ( n13471 , n13470 , n13089 );
and ( n13472 , n13469 , n13471 );
xor ( n13473 , n13438 , n13472 );
xor ( n13474 , n7995 , n7851 );
xor ( n13475 , n11821 , n13257 );
buf ( n13476 , n6399 );
xor ( n13477 , n13475 , n13476 );
buf ( n13478 , n6400 );
xor ( n13479 , n13477 , n13478 );
xor ( n13480 , n13479 , n7014 );
xor ( n13481 , n13474 , n13480 );
not ( n13482 , n13438 );
and ( n13483 , n13482 , n13468 );
xor ( n13484 , n13481 , n13483 );
xor ( n13485 , n12755 , n9046 );
xor ( n13486 , n13485 , n8974 );
not ( n13487 , n6583 );
buf ( n13488 , n6401 );
and ( n13489 , n13487 , n13488 );
buf ( n13490 , n6402 );
xor ( n13491 , n13490 , n13488 );
and ( n13492 , n13491 , n6583 );
or ( n13493 , n13489 , n13492 );
not ( n13494 , n6583 );
buf ( n13495 , n6403 );
and ( n13496 , n13494 , n13495 );
buf ( n13497 , n6404 );
xor ( n13498 , n13497 , n13495 );
and ( n13499 , n13498 , n6583 );
or ( n13500 , n13496 , n13499 );
xor ( n13501 , n13500 , n8348 );
buf ( n13502 , n6405 );
xor ( n13503 , n13501 , n13502 );
buf ( n13504 , n6406 );
xor ( n13505 , n13503 , n13504 );
buf ( n13506 , n6407 );
xor ( n13507 , n13505 , n13506 );
xor ( n13508 , n13493 , n13507 );
xor ( n13509 , n13508 , n10260 );
not ( n13510 , n13509 );
xor ( n13511 , n7461 , n10867 );
xor ( n13512 , n13511 , n9920 );
and ( n13513 , n13510 , n13512 );
xor ( n13514 , n13486 , n13513 );
xor ( n13515 , n13484 , n13514 );
xor ( n13516 , n7008 , n11866 );
xor ( n13517 , n13516 , n10845 );
not ( n13518 , n6583 );
buf ( n13519 , n6408 );
and ( n13520 , n13518 , n13519 );
buf ( n13521 , n6409 );
xor ( n13522 , n13521 , n13519 );
and ( n13523 , n13522 , n6583 );
or ( n13524 , n13520 , n13523 );
not ( n13525 , n6583 );
buf ( n13526 , n6410 );
and ( n13527 , n13525 , n13526 );
buf ( n13528 , n6411 );
xor ( n13529 , n13528 , n13526 );
and ( n13530 , n13529 , n6583 );
or ( n13531 , n13527 , n13530 );
xor ( n13532 , n13524 , n13531 );
xor ( n13533 , n13532 , n7518 );
buf ( n13534 , n6412 );
xor ( n13535 , n13533 , n13534 );
buf ( n13536 , n6413 );
xor ( n13537 , n13535 , n13536 );
xor ( n13538 , n8152 , n13537 );
not ( n13539 , n6583 );
buf ( n13540 , n6414 );
and ( n13541 , n13539 , n13540 );
buf ( n13542 , n6415 );
xor ( n13543 , n13542 , n13540 );
and ( n13544 , n13543 , n6583 );
or ( n13545 , n13541 , n13544 );
not ( n13546 , n6583 );
buf ( n13547 , n6416 );
and ( n13548 , n13546 , n13547 );
buf ( n13549 , n6417 );
xor ( n13550 , n13549 , n13547 );
and ( n13551 , n13550 , n6583 );
or ( n13552 , n13548 , n13551 );
xor ( n13553 , n13545 , n13552 );
xor ( n13554 , n13553 , n8613 );
buf ( n13555 , n6418 );
xor ( n13556 , n13554 , n13555 );
buf ( n13557 , n6419 );
xor ( n13558 , n13556 , n13557 );
xor ( n13559 , n13538 , n13558 );
not ( n13560 , n13559 );
xor ( n13561 , n11971 , n11684 );
xor ( n13562 , n13561 , n11218 );
and ( n13563 , n13560 , n13562 );
xor ( n13564 , n13517 , n13563 );
xor ( n13565 , n13515 , n13564 );
not ( n13566 , n6583 );
buf ( n13567 , n6420 );
and ( n13568 , n13566 , n13567 );
buf ( n13569 , n6421 );
xor ( n13570 , n13569 , n13567 );
and ( n13571 , n13570 , n6583 );
or ( n13572 , n13568 , n13571 );
xor ( n13573 , n13572 , n12683 );
buf ( n13574 , n6422 );
xor ( n13575 , n13573 , n13574 );
buf ( n13576 , n6423 );
xor ( n13577 , n13575 , n13576 );
buf ( n13578 , n6424 );
xor ( n13579 , n13577 , n13578 );
xor ( n13580 , n12291 , n13579 );
xor ( n13581 , n13580 , n12234 );
xor ( n13582 , n12775 , n9699 );
xor ( n13583 , n13582 , n9362 );
not ( n13584 , n13583 );
xor ( n13585 , n11844 , n11560 );
xor ( n13586 , n13585 , n10944 );
and ( n13587 , n13584 , n13586 );
xor ( n13588 , n13581 , n13587 );
xor ( n13589 , n13565 , n13588 );
xor ( n13590 , n7554 , n8127 );
xor ( n13591 , n13590 , n8142 );
xor ( n13592 , n12110 , n6819 );
xor ( n13593 , n13592 , n12347 );
not ( n13594 , n13593 );
xor ( n13595 , n10113 , n12840 );
xor ( n13596 , n13595 , n12856 );
and ( n13597 , n13594 , n13596 );
xor ( n13598 , n13591 , n13597 );
xor ( n13599 , n13589 , n13598 );
xor ( n13600 , n13473 , n13599 );
xor ( n13601 , n13323 , n13149 );
xor ( n13602 , n13601 , n13169 );
not ( n13603 , n6583 );
buf ( n13604 , n6425 );
and ( n13605 , n13603 , n13604 );
buf ( n13606 , n6426 );
xor ( n13607 , n13606 , n13604 );
and ( n13608 , n13607 , n6583 );
or ( n13609 , n13605 , n13608 );
xor ( n13610 , n13609 , n13445 );
buf ( n13611 , n6427 );
xor ( n13612 , n13610 , n13611 );
buf ( n13613 , n6428 );
xor ( n13614 , n13612 , n13613 );
buf ( n13615 , n6429 );
xor ( n13616 , n13614 , n13615 );
buf ( n13617 , n13616 );
not ( n13618 , n6583 );
buf ( n13619 , n6430 );
and ( n13620 , n13618 , n13619 );
buf ( n13621 , n6431 );
xor ( n13622 , n13621 , n13619 );
and ( n13623 , n13622 , n6583 );
or ( n13624 , n13620 , n13623 );
not ( n13625 , n6583 );
buf ( n13626 , n6432 );
and ( n13627 , n13625 , n13626 );
buf ( n13628 , n6433 );
xor ( n13629 , n13628 , n13626 );
and ( n13630 , n13629 , n6583 );
or ( n13631 , n13627 , n13630 );
xor ( n13632 , n13624 , n13631 );
buf ( n13633 , n6434 );
xor ( n13634 , n13632 , n13633 );
buf ( n13635 , n6435 );
xor ( n13636 , n13634 , n13635 );
buf ( n13637 , n6436 );
xor ( n13638 , n13636 , n13637 );
xor ( n13639 , n13617 , n13638 );
not ( n13640 , n13639 );
xor ( n13641 , n11166 , n9942 );
xor ( n13642 , n13641 , n10993 );
and ( n13643 , n13640 , n13642 );
xor ( n13644 , n13602 , n13643 );
xor ( n13645 , n9171 , n8606 );
xor ( n13646 , n8068 , n12733 );
buf ( n13647 , n6437 );
xor ( n13648 , n13646 , n13647 );
buf ( n13649 , n6438 );
xor ( n13650 , n13648 , n13649 );
buf ( n13651 , n6439 );
xor ( n13652 , n13650 , n13651 );
xor ( n13653 , n13645 , n13652 );
xor ( n13654 , n8700 , n10308 );
xor ( n13655 , n13654 , n11410 );
not ( n13656 , n13655 );
xor ( n13657 , n12430 , n13417 );
xor ( n13658 , n13657 , n8412 );
and ( n13659 , n13656 , n13658 );
xor ( n13660 , n13653 , n13659 );
xor ( n13661 , n13644 , n13660 );
xor ( n13662 , n12640 , n12954 );
xor ( n13663 , n13662 , n11739 );
xor ( n13664 , n9280 , n9018 );
xor ( n13665 , n13664 , n12782 );
not ( n13666 , n13665 );
xor ( n13667 , n12210 , n10070 );
not ( n13668 , n6583 );
buf ( n13669 , n6440 );
and ( n13670 , n13668 , n13669 );
buf ( n13671 , n6441 );
xor ( n13672 , n13671 , n13669 );
and ( n13673 , n13672 , n6583 );
or ( n13674 , n13670 , n13673 );
not ( n13675 , n6583 );
buf ( n13676 , n6442 );
and ( n13677 , n13675 , n13676 );
buf ( n13678 , n6443 );
xor ( n13679 , n13678 , n13676 );
and ( n13680 , n13679 , n6583 );
or ( n13681 , n13677 , n13680 );
xor ( n13682 , n13674 , n13681 );
buf ( n13683 , n6444 );
xor ( n13684 , n13682 , n13683 );
xor ( n13685 , n13684 , n11764 );
buf ( n13686 , n6445 );
xor ( n13687 , n13685 , n13686 );
xor ( n13688 , n13667 , n13687 );
and ( n13689 , n13666 , n13688 );
xor ( n13690 , n13663 , n13689 );
xor ( n13691 , n13661 , n13690 );
xor ( n13692 , n10791 , n9715 );
xor ( n13693 , n13692 , n8886 );
not ( n13694 , n6583 );
buf ( n13695 , n6446 );
and ( n13696 , n13694 , n13695 );
buf ( n13697 , n6447 );
xor ( n13698 , n13697 , n13695 );
and ( n13699 , n13698 , n6583 );
or ( n13700 , n13696 , n13699 );
not ( n13701 , n6583 );
buf ( n13702 , n6448 );
and ( n13703 , n13701 , n13702 );
buf ( n13704 , n6449 );
xor ( n13705 , n13704 , n13702 );
and ( n13706 , n13705 , n6583 );
or ( n13707 , n13703 , n13706 );
xor ( n13708 , n13700 , n13707 );
buf ( n13709 , n6450 );
xor ( n13710 , n13708 , n13709 );
buf ( n13711 , n6451 );
xor ( n13712 , n13710 , n13711 );
buf ( n13713 , n6452 );
xor ( n13714 , n13712 , n13713 );
xor ( n13715 , n11781 , n13714 );
not ( n13716 , n6583 );
buf ( n13717 , n6453 );
and ( n13718 , n13716 , n13717 );
buf ( n13719 , n6454 );
xor ( n13720 , n13719 , n13717 );
and ( n13721 , n13720 , n6583 );
or ( n13722 , n13718 , n13721 );
not ( n13723 , n6583 );
buf ( n13724 , n6455 );
and ( n13725 , n13723 , n13724 );
buf ( n13726 , n6456 );
xor ( n13727 , n13726 , n13724 );
and ( n13728 , n13727 , n6583 );
or ( n13729 , n13725 , n13728 );
xor ( n13730 , n13722 , n13729 );
xor ( n13731 , n13730 , n11445 );
buf ( n13732 , n6457 );
xor ( n13733 , n13731 , n13732 );
buf ( n13734 , n6458 );
xor ( n13735 , n13733 , n13734 );
xor ( n13736 , n13715 , n13735 );
not ( n13737 , n13736 );
buf ( n13738 , n6459 );
xor ( n13739 , n13738 , n7051 );
xor ( n13740 , n13739 , n6987 );
and ( n13741 , n13737 , n13740 );
xor ( n13742 , n13693 , n13741 );
xor ( n13743 , n13691 , n13742 );
xor ( n13744 , n12285 , n13579 );
xor ( n13745 , n13744 , n12234 );
xor ( n13746 , n9080 , n11604 );
xor ( n13747 , n13746 , n6849 );
not ( n13748 , n13747 );
xor ( n13749 , n7365 , n12160 );
xor ( n13750 , n13749 , n13068 );
and ( n13751 , n13748 , n13750 );
xor ( n13752 , n13745 , n13751 );
xor ( n13753 , n13743 , n13752 );
xor ( n13754 , n13600 , n13753 );
not ( n13755 , n6583 );
buf ( n13756 , n6460 );
and ( n13757 , n13755 , n13756 );
buf ( n13758 , n6461 );
xor ( n13759 , n13758 , n13756 );
and ( n13760 , n13759 , n6583 );
or ( n13761 , n13757 , n13760 );
not ( n13762 , n6583 );
buf ( n13763 , n6462 );
and ( n13764 , n13762 , n13763 );
buf ( n13765 , n6463 );
xor ( n13766 , n13765 , n13763 );
and ( n13767 , n13766 , n6583 );
or ( n13768 , n13764 , n13767 );
xor ( n13769 , n13761 , n13768 );
buf ( n13770 , n6464 );
xor ( n13771 , n13769 , n13770 );
xor ( n13772 , n13771 , n13191 );
buf ( n13773 , n6465 );
xor ( n13774 , n13772 , n13773 );
xor ( n13775 , n8985 , n13774 );
xor ( n13776 , n13775 , n13537 );
not ( n13777 , n6583 );
buf ( n13778 , n6466 );
and ( n13779 , n13777 , n13778 );
buf ( n13780 , n6467 );
xor ( n13781 , n13780 , n13778 );
and ( n13782 , n13781 , n6583 );
or ( n13783 , n13779 , n13782 );
xor ( n13784 , n13783 , n12858 );
buf ( n13785 , n6468 );
xor ( n13786 , n13784 , n13785 );
buf ( n13787 , n6469 );
xor ( n13788 , n13786 , n13787 );
buf ( n13789 , n6470 );
xor ( n13790 , n13788 , n13789 );
xor ( n13791 , n9872 , n13790 );
xor ( n13792 , n13791 , n11710 );
not ( n13793 , n13792 );
and ( n13794 , n13793 , n13334 );
xor ( n13795 , n13776 , n13794 );
xor ( n13796 , n9222 , n10971 );
xor ( n13797 , n13796 , n6947 );
not ( n13798 , n13797 );
xor ( n13799 , n7672 , n8105 );
xor ( n13800 , n13799 , n6615 );
and ( n13801 , n13798 , n13800 );
xor ( n13802 , n13330 , n13801 );
not ( n13803 , n13776 );
and ( n13804 , n13803 , n13792 );
xor ( n13805 , n13339 , n13804 );
xor ( n13806 , n13802 , n13805 );
xor ( n13807 , n8227 , n12371 );
xor ( n13808 , n13807 , n13225 );
not ( n13809 , n13808 );
xor ( n13810 , n7649 , n8727 );
not ( n13811 , n6583 );
buf ( n13812 , n6471 );
and ( n13813 , n13811 , n13812 );
buf ( n13814 , n6472 );
xor ( n13815 , n13814 , n13812 );
and ( n13816 , n13815 , n6583 );
or ( n13817 , n13813 , n13816 );
xor ( n13818 , n13817 , n12666 );
buf ( n13819 , n6473 );
xor ( n13820 , n13818 , n13819 );
xor ( n13821 , n13820 , n7689 );
buf ( n13822 , n6474 );
xor ( n13823 , n13821 , n13822 );
xor ( n13824 , n13810 , n13823 );
and ( n13825 , n13809 , n13824 );
xor ( n13826 , n13382 , n13825 );
xor ( n13827 , n13806 , n13826 );
xor ( n13828 , n11885 , n8948 );
xor ( n13829 , n13828 , n9972 );
not ( n13830 , n13829 );
xor ( n13831 , n10093 , n11544 );
xor ( n13832 , n13831 , n12840 );
and ( n13833 , n13830 , n13832 );
xor ( n13834 , n13393 , n13833 );
xor ( n13835 , n13827 , n13834 );
xor ( n13836 , n9780 , n11436 );
xor ( n13837 , n13836 , n11560 );
not ( n13838 , n13837 );
xor ( n13839 , n9610 , n10241 );
xor ( n13840 , n13839 , n9739 );
and ( n13841 , n13838 , n13840 );
xor ( n13842 , n13422 , n13841 );
xor ( n13843 , n13835 , n13842 );
xor ( n13844 , n13795 , n13843 );
xor ( n13845 , n8335 , n9229 );
xor ( n13846 , n13845 , n9244 );
xor ( n13847 , n8186 , n13558 );
xor ( n13848 , n13847 , n12492 );
not ( n13849 , n13848 );
xor ( n13850 , n9510 , n6918 );
xor ( n13851 , n13850 , n11386 );
and ( n13852 , n13849 , n13851 );
xor ( n13853 , n13846 , n13852 );
xor ( n13854 , n12868 , n8428 );
xor ( n13855 , n13854 , n10673 );
xor ( n13856 , n8289 , n10166 );
xor ( n13857 , n13856 , n12191 );
not ( n13858 , n13857 );
xor ( n13859 , n6870 , n8822 );
xor ( n13860 , n13859 , n11050 );
and ( n13861 , n13858 , n13860 );
xor ( n13862 , n13855 , n13861 );
xor ( n13863 , n13853 , n13862 );
xor ( n13864 , n7705 , n11978 );
xor ( n13865 , n13864 , n11993 );
xor ( n13866 , n7332 , n11529 );
xor ( n13867 , n13866 , n11544 );
not ( n13868 , n13867 );
xor ( n13869 , n7215 , n8036 );
xor ( n13870 , n13869 , n8058 );
and ( n13871 , n13868 , n13870 );
xor ( n13872 , n13865 , n13871 );
xor ( n13873 , n13863 , n13872 );
xor ( n13874 , n9335 , n12037 );
xor ( n13875 , n13874 , n13579 );
xor ( n13876 , n11272 , n9533 );
xor ( n13877 , n13876 , n8018 );
not ( n13878 , n13877 );
xor ( n13879 , n7885 , n12065 );
xor ( n13880 , n13879 , n12080 );
and ( n13881 , n13878 , n13880 );
xor ( n13882 , n13875 , n13881 );
xor ( n13883 , n13873 , n13882 );
xor ( n13884 , n7463 , n10867 );
xor ( n13885 , n13884 , n9920 );
xor ( n13886 , n13649 , n8083 );
xor ( n13887 , n13886 , n8105 );
not ( n13888 , n13887 );
xor ( n13889 , n12551 , n9877 );
xor ( n13890 , n13889 , n8757 );
and ( n13891 , n13888 , n13890 );
xor ( n13892 , n13885 , n13891 );
xor ( n13893 , n13883 , n13892 );
xor ( n13894 , n13844 , n13893 );
not ( n13895 , n13894 );
not ( n13896 , n13247 );
xor ( n13897 , n12101 , n6797 );
xor ( n13898 , n13897 , n6819 );
and ( n13899 , n13896 , n13898 );
xor ( n13900 , n13210 , n13899 );
xor ( n13901 , n13900 , n13287 );
xor ( n13902 , n13901 , n13425 );
and ( n13903 , n13895 , n13902 );
xor ( n13904 , n13754 , n13903 );
and ( n13905 , n13904 , n6584 );
or ( n13906 , n13436 , n13905 );
and ( n13907 , n13434 , n13906 );
buf ( n13908 , n13907 );
buf ( n13909 , n13908 );
not ( n13910 , n6578 );
not ( n13911 , n6584 );
and ( n13912 , n13911 , n12193 );
xor ( n13913 , n8405 , n12552 );
xor ( n13914 , n13913 , n12573 );
xor ( n13915 , n8184 , n13558 );
xor ( n13916 , n13915 , n12492 );
not ( n13917 , n13916 );
xor ( n13918 , n8763 , n8460 );
xor ( n13919 , n13918 , n8482 );
and ( n13920 , n13917 , n13919 );
xor ( n13921 , n13914 , n13920 );
xor ( n13922 , n6835 , n8807 );
xor ( n13923 , n13922 , n8822 );
xor ( n13924 , n11142 , n9920 );
xor ( n13925 , n13924 , n9942 );
not ( n13926 , n13925 );
xor ( n13927 , n13100 , n8584 );
xor ( n13928 , n13927 , n8606 );
and ( n13929 , n13926 , n13928 );
xor ( n13930 , n13923 , n13929 );
xor ( n13931 , n7640 , n8727 );
xor ( n13932 , n13931 , n13823 );
xor ( n13933 , n6790 , n8018 );
xor ( n13934 , n13933 , n7073 );
not ( n13935 , n13934 );
xor ( n13936 , n11067 , n9262 );
xor ( n13937 , n13936 , n13329 );
and ( n13938 , n13935 , n13937 );
xor ( n13939 , n13932 , n13938 );
xor ( n13940 , n13930 , n13939 );
xor ( n13941 , n8815 , n7368 );
xor ( n13942 , n13941 , n7390 );
not ( n13943 , n13914 );
and ( n13944 , n13943 , n13916 );
xor ( n13945 , n13942 , n13944 );
xor ( n13946 , n13940 , n13945 );
xor ( n13947 , n10300 , n7147 );
not ( n13948 , n6583 );
buf ( n13949 , n6475 );
and ( n13950 , n13948 , n13949 );
buf ( n13951 , n6476 );
xor ( n13952 , n13951 , n13949 );
and ( n13953 , n13952 , n6583 );
or ( n13954 , n13950 , n13953 );
xor ( n13955 , n13954 , n11662 );
buf ( n13956 , n6477 );
xor ( n13957 , n13955 , n13956 );
xor ( n13958 , n13957 , n13112 );
buf ( n13959 , n6478 );
xor ( n13960 , n13958 , n13959 );
xor ( n13961 , n13947 , n13960 );
not ( n13962 , n6583 );
buf ( n13963 , n6479 );
and ( n13964 , n13962 , n13963 );
buf ( n13965 , n6480 );
xor ( n13966 , n13965 , n13963 );
and ( n13967 , n13966 , n6583 );
or ( n13968 , n13964 , n13967 );
buf ( n13969 , n6481 );
xor ( n13970 , n13968 , n13969 );
buf ( n13971 , n6482 );
xor ( n13972 , n13970 , n13971 );
buf ( n13973 , n6483 );
xor ( n13974 , n13972 , n13973 );
buf ( n13975 , n6484 );
xor ( n13976 , n13974 , n13975 );
xor ( n13977 , n10404 , n13976 );
not ( n13978 , n6583 );
buf ( n13979 , n6485 );
and ( n13980 , n13978 , n13979 );
buf ( n13981 , n6486 );
xor ( n13982 , n13981 , n13979 );
and ( n13983 , n13982 , n6583 );
or ( n13984 , n13980 , n13983 );
not ( n13985 , n6583 );
buf ( n13986 , n6487 );
and ( n13987 , n13985 , n13986 );
buf ( n13988 , n6488 );
xor ( n13989 , n13988 , n13986 );
and ( n13990 , n13989 , n6583 );
or ( n13991 , n13987 , n13990 );
xor ( n13992 , n13984 , n13991 );
buf ( n13993 , n6489 );
xor ( n13994 , n13992 , n13993 );
xor ( n13995 , n13994 , n11564 );
xor ( n13996 , n13995 , n10678 );
xor ( n13997 , n13977 , n13996 );
not ( n13998 , n13997 );
xor ( n13999 , n11342 , n10349 );
xor ( n14000 , n13999 , n7319 );
and ( n14001 , n13998 , n14000 );
xor ( n14002 , n13961 , n14001 );
xor ( n14003 , n13946 , n14002 );
xor ( n14004 , n9055 , n11590 );
xor ( n14005 , n14004 , n11604 );
xor ( n14006 , n9102 , n10142 );
xor ( n14007 , n14006 , n6659 );
not ( n14008 , n14007 );
not ( n14009 , n6583 );
buf ( n14010 , n6490 );
and ( n14011 , n14009 , n14010 );
buf ( n14012 , n6491 );
xor ( n14013 , n14012 , n14010 );
and ( n14014 , n14013 , n6583 );
or ( n14015 , n14011 , n14014 );
not ( n14016 , n6583 );
buf ( n14017 , n6492 );
and ( n14018 , n14016 , n14017 );
buf ( n14019 , n6493 );
xor ( n14020 , n14019 , n14017 );
and ( n14021 , n14020 , n6583 );
or ( n14022 , n14018 , n14021 );
xor ( n14023 , n14015 , n14022 );
buf ( n14024 , n6494 );
xor ( n14025 , n14023 , n14024 );
buf ( n14026 , n6495 );
xor ( n14027 , n14025 , n14026 );
buf ( n14028 , n6496 );
xor ( n14029 , n14027 , n14028 );
xor ( n14030 , n8943 , n14029 );
not ( n14031 , n6583 );
buf ( n14032 , n6497 );
and ( n14033 , n14031 , n14032 );
buf ( n14034 , n6498 );
xor ( n14035 , n14034 , n14032 );
and ( n14036 , n14035 , n6583 );
or ( n14037 , n14033 , n14036 );
not ( n14038 , n6583 );
buf ( n14039 , n6499 );
and ( n14040 , n14038 , n14039 );
buf ( n14041 , n6500 );
xor ( n14042 , n14041 , n14039 );
and ( n14043 , n14042 , n6583 );
or ( n14044 , n14040 , n14043 );
xor ( n14045 , n14037 , n14044 );
buf ( n14046 , n6501 );
xor ( n14047 , n14045 , n14046 );
buf ( n14048 , n6502 );
xor ( n14049 , n14047 , n14048 );
buf ( n14050 , n6503 );
xor ( n14051 , n14049 , n14050 );
xor ( n14052 , n14030 , n14051 );
and ( n14053 , n14008 , n14052 );
xor ( n14054 , n14005 , n14053 );
xor ( n14055 , n14003 , n14054 );
xor ( n14056 , n13921 , n14055 );
xor ( n14057 , n9756 , n11147 );
xor ( n14058 , n14057 , n11169 );
xor ( n14059 , n12344 , n7095 );
xor ( n14060 , n14059 , n8992 );
not ( n14061 , n14060 );
xor ( n14062 , n12855 , n12292 );
not ( n14063 , n6583 );
buf ( n14064 , n6504 );
and ( n14065 , n14063 , n14064 );
buf ( n14066 , n6505 );
xor ( n14067 , n14066 , n14064 );
and ( n14068 , n14067 , n6583 );
or ( n14069 , n14065 , n14068 );
not ( n14070 , n6583 );
buf ( n14071 , n6506 );
and ( n14072 , n14070 , n14071 );
buf ( n14073 , n6507 );
xor ( n14074 , n14073 , n14071 );
and ( n14075 , n14074 , n6583 );
or ( n14076 , n14072 , n14075 );
xor ( n14077 , n14069 , n14076 );
buf ( n14078 , n6508 );
xor ( n14079 , n14077 , n14078 );
xor ( n14080 , n14079 , n12220 );
buf ( n14081 , n6509 );
xor ( n14082 , n14080 , n14081 );
xor ( n14083 , n14062 , n14082 );
and ( n14084 , n14061 , n14083 );
xor ( n14085 , n14058 , n14084 );
xor ( n14086 , n13144 , n8653 );
xor ( n14087 , n14086 , n12433 );
xor ( n14088 , n8102 , n8318 );
xor ( n14089 , n14088 , n8340 );
not ( n14090 , n14089 );
xor ( n14091 , n9068 , n11590 );
xor ( n14092 , n14091 , n11604 );
and ( n14093 , n14090 , n14092 );
xor ( n14094 , n14087 , n14093 );
xor ( n14095 , n14085 , n14094 );
xor ( n14096 , n8630 , n8142 );
xor ( n14097 , n14096 , n10308 );
xor ( n14098 , n11322 , n10327 );
xor ( n14099 , n14098 , n10349 );
not ( n14100 , n14099 );
xor ( n14101 , n11385 , n9897 );
xor ( n14102 , n14101 , n9046 );
and ( n14103 , n14100 , n14102 );
xor ( n14104 , n14097 , n14103 );
xor ( n14105 , n14095 , n14104 );
xor ( n14106 , n11942 , n13246 );
xor ( n14107 , n14106 , n7173 );
not ( n14108 , n6583 );
buf ( n14109 , n6510 );
and ( n14110 , n14108 , n14109 );
buf ( n14111 , n6511 );
xor ( n14112 , n14111 , n14109 );
and ( n14113 , n14112 , n6583 );
or ( n14114 , n14110 , n14113 );
not ( n14115 , n6583 );
buf ( n14116 , n6512 );
and ( n14117 , n14115 , n14116 );
buf ( n14118 , n6513 );
xor ( n14119 , n14118 , n14116 );
and ( n14120 , n14119 , n6583 );
or ( n14121 , n14117 , n14120 );
xor ( n14122 , n14114 , n14121 );
buf ( n14123 , n6514 );
xor ( n14124 , n14122 , n14123 );
buf ( n14125 , n6515 );
xor ( n14126 , n14124 , n14125 );
buf ( n14127 , n6516 );
xor ( n14128 , n14126 , n14127 );
xor ( n14129 , n10031 , n14128 );
xor ( n14130 , n14129 , n12721 );
not ( n14131 , n14130 );
xor ( n14132 , n9427 , n8863 );
xor ( n14133 , n14132 , n13282 );
and ( n14134 , n14131 , n14133 );
xor ( n14135 , n14107 , n14134 );
xor ( n14136 , n14105 , n14135 );
buf ( n14137 , n6517 );
xor ( n14138 , n14137 , n6987 );
xor ( n14139 , n14138 , n7009 );
xor ( n14140 , n7513 , n9615 );
xor ( n14141 , n14140 , n8584 );
not ( n14142 , n14141 );
xor ( n14143 , n13615 , n11072 );
xor ( n14144 , n14143 , n13467 );
and ( n14145 , n14142 , n14144 );
xor ( n14146 , n14139 , n14145 );
xor ( n14147 , n14136 , n14146 );
xor ( n14148 , n14056 , n14147 );
xor ( n14149 , n12692 , n10012 );
xor ( n14150 , n14149 , n10034 );
xor ( n14151 , n12753 , n9046 );
xor ( n14152 , n14151 , n8974 );
not ( n14153 , n14152 );
xor ( n14154 , n9139 , n12804 );
xor ( n14155 , n14154 , n7926 );
and ( n14156 , n14153 , n14155 );
xor ( n14157 , n14150 , n14156 );
xor ( n14158 , n8285 , n10166 );
xor ( n14159 , n14158 , n12191 );
xor ( n14160 , n6942 , n12915 );
xor ( n14161 , n14160 , n9285 );
not ( n14162 , n14161 );
xor ( n14163 , n8632 , n8142 );
xor ( n14164 , n14163 , n10308 );
and ( n14165 , n14162 , n14164 );
xor ( n14166 , n14159 , n14165 );
xor ( n14167 , n13298 , n8189 );
xor ( n14168 , n14167 , n10822 );
buf ( n14169 , n6518 );
xor ( n14170 , n14169 , n8766 );
xor ( n14171 , n14170 , n12371 );
not ( n14172 , n14171 );
xor ( n14173 , n8680 , n9307 );
xor ( n14174 , n14173 , n13507 );
and ( n14175 , n14172 , n14174 );
xor ( n14176 , n14168 , n14175 );
xor ( n14177 , n14166 , n14176 );
xor ( n14178 , n7312 , n11947 );
xor ( n14179 , n14178 , n11529 );
xor ( n14180 , n11213 , n12647 );
xor ( n14181 , n14180 , n12662 );
not ( n14182 , n14181 );
xor ( n14183 , n7186 , n12015 );
xor ( n14184 , n14183 , n12037 );
and ( n14185 , n14182 , n14184 );
xor ( n14186 , n14179 , n14185 );
xor ( n14187 , n14177 , n14186 );
xor ( n14188 , n7002 , n11866 );
xor ( n14189 , n14188 , n10845 );
not ( n14190 , n14150 );
and ( n14191 , n14190 , n14152 );
xor ( n14192 , n14189 , n14191 );
xor ( n14193 , n14187 , n14192 );
xor ( n14194 , n7879 , n12065 );
xor ( n14195 , n14194 , n12080 );
xor ( n14196 , n9173 , n8606 );
xor ( n14197 , n14196 , n13652 );
not ( n14198 , n14197 );
xor ( n14199 , n8314 , n10993 );
xor ( n14200 , n14199 , n9229 );
and ( n14201 , n14198 , n14200 );
xor ( n14202 , n14195 , n14201 );
xor ( n14203 , n14193 , n14202 );
xor ( n14204 , n14157 , n14203 );
xor ( n14205 , n7144 , n10603 );
xor ( n14206 , n14205 , n10619 );
xor ( n14207 , n6796 , n8018 );
xor ( n14208 , n14207 , n7073 );
not ( n14209 , n14208 );
xor ( n14210 , n9863 , n13790 );
xor ( n14211 , n14210 , n11710 );
and ( n14212 , n14209 , n14211 );
xor ( n14213 , n14206 , n14212 );
xor ( n14214 , n8366 , n9362 );
xor ( n14215 , n14214 , n9384 );
xor ( n14216 , n7599 , n13616 );
xor ( n14217 , n14216 , n13638 );
not ( n14218 , n14217 );
xor ( n14219 , n6738 , n9809 );
xor ( n14220 , n14219 , n9825 );
and ( n14221 , n14218 , n14220 );
xor ( n14222 , n14215 , n14221 );
xor ( n14223 , n14213 , n14222 );
xor ( n14224 , n11510 , n10120 );
xor ( n14225 , n14224 , n10012 );
xor ( n14226 , n13536 , n7533 );
xor ( n14227 , n14226 , n7555 );
not ( n14228 , n14227 );
xor ( n14229 , n11696 , n12873 );
xor ( n14230 , n14229 , n12978 );
and ( n14231 , n14228 , n14230 );
xor ( n14232 , n14225 , n14231 );
xor ( n14233 , n14223 , n14232 );
xor ( n14234 , n12122 , n6819 );
xor ( n14235 , n14234 , n12347 );
xor ( n14236 , n8907 , n9069 );
xor ( n14237 , n14236 , n9085 );
not ( n14238 , n14237 );
xor ( n14239 , n9447 , n10497 );
xor ( n14240 , n14239 , n13714 );
and ( n14241 , n14238 , n14240 );
xor ( n14242 , n14235 , n14241 );
xor ( n14243 , n14233 , n14242 );
xor ( n14244 , n10968 , n7686 );
xor ( n14245 , n14244 , n12915 );
not ( n14246 , n6583 );
buf ( n14247 , n6519 );
and ( n14248 , n14246 , n14247 );
buf ( n14249 , n6520 );
xor ( n14250 , n14249 , n14247 );
and ( n14251 , n14250 , n6583 );
or ( n14252 , n14248 , n14251 );
xor ( n14253 , n12356 , n14252 );
xor ( n14254 , n14253 , n14169 );
buf ( n14255 , n6521 );
xor ( n14256 , n14254 , n14255 );
buf ( n14257 , n6522 );
xor ( n14258 , n14256 , n14257 );
xor ( n14259 , n10672 , n14258 );
xor ( n14260 , n14259 , n8234 );
not ( n14261 , n14260 );
xor ( n14262 , n13453 , n13329 );
xor ( n14263 , n14262 , n9855 );
and ( n14264 , n14261 , n14263 );
xor ( n14265 , n14245 , n14264 );
xor ( n14266 , n14243 , n14265 );
xor ( n14267 , n14204 , n14266 );
not ( n14268 , n14267 );
not ( n14269 , n9019 );
and ( n14270 , n14269 , n11170 );
xor ( n14271 , n8994 , n14270 );
xor ( n14272 , n14271 , n9022 );
xor ( n14273 , n12079 , n9140 );
xor ( n14274 , n14273 , n9161 );
xor ( n14275 , n10957 , n7686 );
xor ( n14276 , n14275 , n12915 );
not ( n14277 , n14276 );
xor ( n14278 , n7625 , n8705 );
xor ( n14279 , n14278 , n8727 );
and ( n14280 , n14277 , n14279 );
xor ( n14281 , n14274 , n14280 );
xor ( n14282 , n9760 , n11147 );
xor ( n14283 , n14282 , n11169 );
xor ( n14284 , n11285 , n7319 );
xor ( n14285 , n14284 , n7335 );
not ( n14286 , n14285 );
xor ( n14287 , n9255 , n13089 );
xor ( n14288 , n14287 , n13149 );
and ( n14289 , n14286 , n14288 );
xor ( n14290 , n14283 , n14289 );
xor ( n14291 , n14281 , n14290 );
xor ( n14292 , n7367 , n12160 );
xor ( n14293 , n14292 , n13068 );
xor ( n14294 , n12903 , n6636 );
xor ( n14295 , n14294 , n9018 );
not ( n14296 , n14295 );
xor ( n14297 , n12401 , n10282 );
xor ( n14298 , n14297 , n8789 );
and ( n14299 , n14296 , n14298 );
xor ( n14300 , n14293 , n14299 );
xor ( n14301 , n14291 , n14300 );
not ( n14302 , n6583 );
buf ( n14303 , n6523 );
and ( n14304 , n14302 , n14303 );
buf ( n14305 , n6524 );
xor ( n14306 , n14305 , n14303 );
and ( n14307 , n14306 , n6583 );
or ( n14308 , n14304 , n14307 );
not ( n14309 , n6583 );
buf ( n14310 , n6525 );
and ( n14311 , n14309 , n14310 );
buf ( n14312 , n6526 );
xor ( n14313 , n14312 , n14310 );
and ( n14314 , n14313 , n6583 );
or ( n14315 , n14311 , n14314 );
xor ( n14316 , n14308 , n14315 );
buf ( n14317 , n6527 );
xor ( n14318 , n14316 , n14317 );
xor ( n14319 , n14318 , n13738 );
xor ( n14320 , n14319 , n9662 );
xor ( n14321 , n14028 , n14320 );
not ( n14322 , n6583 );
buf ( n14323 , n6528 );
and ( n14324 , n14322 , n14323 );
buf ( n14325 , n6529 );
xor ( n14326 , n14325 , n14323 );
and ( n14327 , n14326 , n6583 );
or ( n14328 , n14324 , n14327 );
xor ( n14329 , n14328 , n6966 );
xor ( n14330 , n14329 , n14137 );
buf ( n14331 , n6530 );
xor ( n14332 , n14330 , n14331 );
buf ( n14333 , n6531 );
xor ( n14334 , n14332 , n14333 );
xor ( n14335 , n14321 , n14334 );
xor ( n14336 , n8242 , n13225 );
xor ( n14337 , n14336 , n13246 );
not ( n14338 , n14337 );
xor ( n14339 , n11380 , n9897 );
xor ( n14340 , n14339 , n9046 );
and ( n14341 , n14338 , n14340 );
xor ( n14342 , n14335 , n14341 );
xor ( n14343 , n14301 , n14342 );
xor ( n14344 , n8291 , n10166 );
xor ( n14345 , n14344 , n12191 );
xor ( n14346 , n9928 , n9200 );
xor ( n14347 , n14346 , n13188 );
not ( n14348 , n14347 );
not ( n14349 , n6583 );
buf ( n14350 , n6532 );
and ( n14351 , n14349 , n14350 );
buf ( n14352 , n6533 );
xor ( n14353 , n14352 , n14350 );
and ( n14354 , n14353 , n6583 );
or ( n14355 , n14351 , n14354 );
xor ( n14356 , n14355 , n8932 );
xor ( n14357 , n14356 , n8948 );
and ( n14358 , n14348 , n14357 );
xor ( n14359 , n14345 , n14358 );
xor ( n14360 , n14343 , n14359 );
xor ( n14361 , n14272 , n14360 );
and ( n14362 , n14268 , n14361 );
xor ( n14363 , n14148 , n14362 );
and ( n14364 , n14363 , n6584 );
or ( n14365 , n13912 , n14364 );
and ( n14366 , n13910 , n14365 );
buf ( n14367 , n14366 );
buf ( n14368 , n14367 );
not ( n14369 , n6578 );
not ( n14370 , n6584 );
and ( n14371 , n14370 , n8316 );
xor ( n14372 , n7233 , n8058 );
not ( n14373 , n6583 );
buf ( n14374 , n6534 );
and ( n14375 , n14373 , n14374 );
buf ( n14376 , n6535 );
xor ( n14377 , n14376 , n14374 );
and ( n14378 , n14377 , n6583 );
or ( n14379 , n14375 , n14378 );
not ( n14380 , n6583 );
buf ( n14381 , n6536 );
and ( n14382 , n14380 , n14381 );
buf ( n14383 , n6537 );
xor ( n14384 , n14383 , n14381 );
and ( n14385 , n14384 , n6583 );
or ( n14386 , n14382 , n14385 );
xor ( n14387 , n14379 , n14386 );
buf ( n14388 , n6538 );
xor ( n14389 , n14387 , n14388 );
xor ( n14390 , n14389 , n13289 );
buf ( n14391 , n6539 );
xor ( n14392 , n14390 , n14391 );
xor ( n14393 , n14372 , n14392 );
xor ( n14394 , n7425 , n6871 );
not ( n14395 , n6583 );
buf ( n14396 , n6540 );
and ( n14397 , n14395 , n14396 );
buf ( n14398 , n6541 );
xor ( n14399 , n14398 , n14396 );
and ( n14400 , n14399 , n6583 );
or ( n14401 , n14397 , n14400 );
xor ( n14402 , n14401 , n11031 );
buf ( n14403 , n6542 );
xor ( n14404 , n14402 , n14403 );
buf ( n14405 , n6543 );
xor ( n14406 , n14404 , n14405 );
buf ( n14407 , n6544 );
xor ( n14408 , n14406 , n14407 );
xor ( n14409 , n14394 , n14408 );
not ( n14410 , n14409 );
xor ( n14411 , n13281 , n9787 );
xor ( n14412 , n14411 , n11850 );
and ( n14413 , n14410 , n14412 );
xor ( n14414 , n14393 , n14413 );
xor ( n14415 , n8159 , n13537 );
xor ( n14416 , n14415 , n13558 );
not ( n14417 , n14393 );
and ( n14418 , n14417 , n14409 );
xor ( n14419 , n14416 , n14418 );
xor ( n14420 , n8800 , n11650 );
xor ( n14421 , n14420 , n7368 );
xor ( n14422 , n10966 , n7686 );
xor ( n14423 , n14422 , n12915 );
not ( n14424 , n14423 );
xor ( n14425 , n7552 , n8127 );
xor ( n14426 , n14425 , n8142 );
and ( n14427 , n14424 , n14426 );
xor ( n14428 , n14421 , n14427 );
xor ( n14429 , n14419 , n14428 );
xor ( n14430 , n12184 , n8683 );
not ( n14431 , n6583 );
buf ( n14432 , n6545 );
and ( n14433 , n14431 , n14432 );
buf ( n14434 , n6546 );
xor ( n14435 , n14434 , n14432 );
and ( n14436 , n14435 , n6583 );
or ( n14437 , n14433 , n14436 );
xor ( n14438 , n13493 , n14437 );
buf ( n14439 , n6547 );
xor ( n14440 , n14438 , n14439 );
buf ( n14441 , n6548 );
xor ( n14442 , n14440 , n14441 );
buf ( n14443 , n6549 );
xor ( n14444 , n14442 , n14443 );
xor ( n14445 , n14430 , n14444 );
xor ( n14446 , n9850 , n13169 );
xor ( n14447 , n14446 , n13790 );
not ( n14448 , n14447 );
xor ( n14449 , n10257 , n8388 );
xor ( n14450 , n14449 , n12601 );
and ( n14451 , n14448 , n14450 );
xor ( n14452 , n14445 , n14451 );
xor ( n14453 , n14429 , n14452 );
xor ( n14454 , n14076 , n12234 );
xor ( n14455 , n14454 , n6896 );
xor ( n14456 , n10547 , n10915 );
xor ( n14457 , n14456 , n10142 );
not ( n14458 , n14457 );
not ( n14459 , n6583 );
buf ( n14460 , n6550 );
and ( n14461 , n14459 , n14460 );
buf ( n14462 , n6551 );
xor ( n14463 , n14462 , n14460 );
and ( n14464 , n14463 , n6583 );
or ( n14465 , n14461 , n14464 );
not ( n14466 , n6583 );
buf ( n14467 , n6552 );
and ( n14468 , n14466 , n14467 );
buf ( n14469 , n6553 );
xor ( n14470 , n14469 , n14467 );
and ( n14471 , n14470 , n6583 );
or ( n14472 , n14468 , n14471 );
xor ( n14473 , n14465 , n14472 );
buf ( n14474 , n6554 );
xor ( n14475 , n14473 , n14474 );
buf ( n14476 , n6555 );
xor ( n14477 , n14475 , n14476 );
buf ( n14478 , n6556 );
xor ( n14479 , n14477 , n14478 );
xor ( n14480 , n10216 , n14479 );
xor ( n14481 , n14480 , n7886 );
and ( n14482 , n14458 , n14481 );
xor ( n14483 , n14455 , n14482 );
xor ( n14484 , n14453 , n14483 );
xor ( n14485 , n12514 , n13735 );
xor ( n14486 , n14485 , n13976 );
xor ( n14487 , n9892 , n7289 );
xor ( n14488 , n14487 , n12102 );
not ( n14489 , n14488 );
xor ( n14490 , n7070 , n13358 );
xor ( n14491 , n14490 , n13378 );
and ( n14492 , n14489 , n14491 );
xor ( n14493 , n14486 , n14492 );
xor ( n14494 , n14484 , n14493 );
xor ( n14495 , n14414 , n14494 );
xor ( n14496 , n14495 , n10977 );
xor ( n14497 , n7264 , n11805 );
xor ( n14498 , n14497 , n11275 );
xor ( n14499 , n9808 , n11786 );
xor ( n14500 , n14499 , n12521 );
not ( n14501 , n14500 );
xor ( n14502 , n7414 , n6871 );
xor ( n14503 , n14502 , n14408 );
and ( n14504 , n14501 , n14503 );
xor ( n14505 , n14498 , n14504 );
xor ( n14506 , n10029 , n14128 );
xor ( n14507 , n14506 , n12721 );
xor ( n14508 , n9784 , n11436 );
xor ( n14509 , n14508 , n11560 );
not ( n14510 , n14509 );
buf ( n14511 , n6557 );
xor ( n14512 , n14511 , n14444 );
xor ( n14513 , n14512 , n12393 );
and ( n14514 , n14510 , n14513 );
xor ( n14515 , n14507 , n14514 );
xor ( n14516 , n14046 , n14334 );
xor ( n14517 , n14516 , n10584 );
not ( n14518 , n14498 );
and ( n14519 , n14518 , n14500 );
xor ( n14520 , n14517 , n14519 );
xor ( n14521 , n14515 , n14520 );
xor ( n14522 , n8903 , n9069 );
xor ( n14523 , n14522 , n9085 );
xor ( n14524 , n8080 , n11169 );
xor ( n14525 , n14524 , n8318 );
not ( n14526 , n14525 );
xor ( n14527 , n8529 , n11238 );
xor ( n14528 , n14527 , n9406 );
and ( n14529 , n14526 , n14528 );
xor ( n14530 , n14523 , n14529 );
xor ( n14531 , n14521 , n14530 );
xor ( n14532 , n9224 , n10971 );
xor ( n14533 , n14532 , n6947 );
xor ( n14534 , n9381 , n11100 );
xor ( n14535 , n14534 , n10893 );
not ( n14536 , n14535 );
xor ( n14537 , n7709 , n11978 );
xor ( n14538 , n14537 , n11993 );
and ( n14539 , n14536 , n14538 );
xor ( n14540 , n14533 , n14539 );
xor ( n14541 , n14531 , n14540 );
xor ( n14542 , n7330 , n11529 );
xor ( n14543 , n14542 , n11544 );
xor ( n14544 , n12034 , n11513 );
xor ( n14545 , n14544 , n12696 );
not ( n14546 , n14545 );
xor ( n14547 , n7050 , n11892 );
xor ( n14548 , n14547 , n11907 );
and ( n14549 , n14546 , n14548 );
xor ( n14550 , n14543 , n14549 );
xor ( n14551 , n14541 , n14550 );
xor ( n14552 , n14505 , n14551 );
xor ( n14553 , n10259 , n8388 );
xor ( n14554 , n14553 , n12601 );
not ( n14555 , n11823 );
and ( n14556 , n14555 , n11807 );
xor ( n14557 , n14554 , n14556 );
xor ( n14558 , n13734 , n11459 );
xor ( n14559 , n14558 , n11474 );
not ( n14560 , n11828 );
and ( n14561 , n14560 , n11851 );
xor ( n14562 , n14559 , n14561 );
xor ( n14563 , n14557 , n14562 );
xor ( n14564 , n8840 , n6659 );
xor ( n14565 , n14564 , n6681 );
not ( n14566 , n11908 );
and ( n14567 , n14566 , n11910 );
xor ( n14568 , n14565 , n14567 );
xor ( n14569 , n14563 , n14568 );
xor ( n14570 , n11217 , n12647 );
xor ( n14571 , n14570 , n12662 );
not ( n14572 , n11925 );
and ( n14573 , n14572 , n11948 );
xor ( n14574 , n14571 , n14573 );
xor ( n14575 , n14569 , n14574 );
xor ( n14576 , n9971 , n14051 );
xor ( n14577 , n14576 , n12931 );
not ( n14578 , n11957 );
and ( n14579 , n14578 , n11994 );
xor ( n14580 , n14577 , n14579 );
xor ( n14581 , n14575 , n14580 );
xor ( n14582 , n14552 , n14581 );
not ( n14583 , n14582 );
xor ( n14584 , n11891 , n8948 );
xor ( n14585 , n14584 , n9972 );
xor ( n14586 , n13366 , n7216 );
xor ( n14587 , n14586 , n7238 );
not ( n14588 , n14587 );
and ( n14589 , n14588 , n7655 );
xor ( n14590 , n14585 , n14589 );
xor ( n14591 , n9824 , n12521 );
xor ( n14592 , n14591 , n10411 );
not ( n14593 , n14592 );
xor ( n14594 , n7059 , n13358 );
xor ( n14595 , n14594 , n13378 );
and ( n14596 , n14593 , n14595 );
xor ( n14597 , n7470 , n14596 );
buf ( n14598 , n6558 );
xor ( n14599 , n14598 , n7267 );
xor ( n14600 , n14599 , n7289 );
not ( n14601 , n14600 );
xor ( n14602 , n9271 , n9018 );
xor ( n14603 , n14602 , n12782 );
and ( n14604 , n14601 , n14603 );
xor ( n14605 , n7601 , n14604 );
xor ( n14606 , n14597 , n14605 );
not ( n14607 , n14585 );
and ( n14608 , n14607 , n14587 );
xor ( n14609 , n7712 , n14608 );
xor ( n14610 , n14606 , n14609 );
xor ( n14611 , n12014 , n11497 );
xor ( n14612 , n14611 , n11513 );
not ( n14613 , n14612 );
xor ( n14614 , n8262 , n9244 );
xor ( n14615 , n14614 , n10166 );
and ( n14616 , n14613 , n14615 );
xor ( n14617 , n7852 , n14616 );
xor ( n14618 , n14610 , n14617 );
xor ( n14619 , n8057 , n9639 );
xor ( n14620 , n14619 , n9660 );
not ( n14621 , n14620 );
xor ( n14622 , n11261 , n9533 );
xor ( n14623 , n14622 , n8018 );
and ( n14624 , n14621 , n14623 );
xor ( n14625 , n7949 , n14624 );
xor ( n14626 , n14618 , n14625 );
xor ( n14627 , n14590 , n14626 );
xor ( n14628 , n7202 , n8036 );
xor ( n14629 , n14628 , n8058 );
xor ( n14630 , n13063 , n7579 );
xor ( n14631 , n14630 , n7600 );
not ( n14632 , n14631 );
xor ( n14633 , n6866 , n8822 );
xor ( n14634 , n14633 , n11050 );
and ( n14635 , n14632 , n14634 );
xor ( n14636 , n14629 , n14635 );
xor ( n14637 , n9685 , n12191 );
not ( n14638 , n6583 );
buf ( n14639 , n6559 );
and ( n14640 , n14638 , n14639 );
buf ( n14641 , n6560 );
xor ( n14642 , n14641 , n14639 );
and ( n14643 , n14642 , n6583 );
or ( n14644 , n14640 , n14643 );
buf ( n14645 , n6561 );
xor ( n14646 , n14644 , n14645 );
buf ( n14647 , n6562 );
xor ( n14648 , n14646 , n14647 );
buf ( n14649 , n6563 );
xor ( n14650 , n14648 , n14649 );
xor ( n14651 , n14650 , n14511 );
xor ( n14652 , n14637 , n14651 );
xor ( n14653 , n9608 , n10241 );
xor ( n14654 , n14653 , n9739 );
not ( n14655 , n14654 );
xor ( n14656 , n8122 , n13304 );
xor ( n14657 , n14656 , n7125 );
and ( n14658 , n14655 , n14657 );
xor ( n14659 , n14652 , n14658 );
xor ( n14660 , n14636 , n14659 );
xor ( n14661 , n8044 , n9639 );
xor ( n14662 , n14661 , n9660 );
xor ( n14663 , n8720 , n11410 );
xor ( n14664 , n14663 , n7710 );
not ( n14665 , n14664 );
xor ( n14666 , n6610 , n8340 );
xor ( n14667 , n14666 , n8270 );
and ( n14668 , n14665 , n14667 );
xor ( n14669 , n14662 , n14668 );
xor ( n14670 , n14660 , n14669 );
xor ( n14671 , n6955 , n9285 );
xor ( n14672 , n14671 , n9307 );
not ( n14673 , n6583 );
buf ( n14674 , n6564 );
and ( n14675 , n14673 , n14674 );
buf ( n14676 , n6565 );
xor ( n14677 , n14676 , n14674 );
and ( n14678 , n14677 , n6583 );
or ( n14679 , n14675 , n14678 );
xor ( n14680 , n14679 , n13282 );
xor ( n14681 , n14680 , n14479 );
not ( n14682 , n14681 );
xor ( n14683 , n10470 , n11761 );
xor ( n14684 , n14683 , n12308 );
and ( n14685 , n14682 , n14684 );
xor ( n14686 , n14672 , n14685 );
xor ( n14687 , n14670 , n14686 );
xor ( n14688 , n12743 , n9046 );
xor ( n14689 , n14688 , n8974 );
xor ( n14690 , n12009 , n11497 );
xor ( n14691 , n14690 , n11513 );
not ( n14692 , n14691 );
xor ( n14693 , n12075 , n9140 );
xor ( n14694 , n14693 , n9161 );
and ( n14695 , n14692 , n14694 );
xor ( n14696 , n14689 , n14695 );
xor ( n14697 , n14687 , n14696 );
xor ( n14698 , n14627 , n14697 );
and ( n14699 , n14583 , n14698 );
xor ( n14700 , n14496 , n14699 );
and ( n14701 , n14700 , n6584 );
or ( n14702 , n14371 , n14701 );
and ( n14703 , n14369 , n14702 );
buf ( n14704 , n14703 );
buf ( n14705 , n14704 );
not ( n14706 , n6578 );
not ( n14707 , n6584 );
and ( n14708 , n14707 , n12119 );
not ( n14709 , n8823 );
and ( n14710 , n14709 , n11079 );
xor ( n14711 , n8791 , n14710 );
xor ( n14712 , n14711 , n9022 );
xor ( n14713 , n14712 , n14360 );
xor ( n14714 , n8973 , n12125 );
xor ( n14715 , n14714 , n8036 );
xor ( n14716 , n6651 , n9583 );
xor ( n14717 , n14716 , n9598 );
not ( n14718 , n14717 );
xor ( n14719 , n7361 , n12160 );
xor ( n14720 , n14719 , n13068 );
and ( n14721 , n14718 , n14720 );
xor ( n14722 , n14715 , n14721 );
xor ( n14723 , n9696 , n12191 );
xor ( n14724 , n14723 , n14651 );
xor ( n14725 , n7468 , n10867 );
xor ( n14726 , n14725 , n9920 );
not ( n14727 , n14726 );
xor ( n14728 , n12459 , n13823 );
xor ( n14729 , n14728 , n12954 );
and ( n14730 , n14727 , n14729 );
xor ( n14731 , n14724 , n14730 );
xor ( n14732 , n11344 , n10349 );
xor ( n14733 , n14732 , n7319 );
xor ( n14734 , n8141 , n7125 );
xor ( n14735 , n14734 , n7147 );
not ( n14736 , n14735 );
xor ( n14737 , n9414 , n8863 );
xor ( n14738 , n14737 , n13282 );
and ( n14739 , n14736 , n14738 );
xor ( n14740 , n14733 , n14739 );
xor ( n14741 , n14731 , n14740 );
xor ( n14742 , n7993 , n7851 );
xor ( n14743 , n14742 , n13480 );
xor ( n14744 , n10970 , n7686 );
xor ( n14745 , n14744 , n12915 );
not ( n14746 , n14745 );
xor ( n14747 , n12948 , n6705 );
xor ( n14748 , n14747 , n6727 );
and ( n14749 , n14746 , n14748 );
xor ( n14750 , n14743 , n14749 );
xor ( n14751 , n14741 , n14750 );
xor ( n14752 , n9758 , n11147 );
xor ( n14753 , n14752 , n11169 );
not ( n14754 , n14715 );
and ( n14755 , n14754 , n14717 );
xor ( n14756 , n14753 , n14755 );
xor ( n14757 , n14751 , n14756 );
xor ( n14758 , n9874 , n13790 );
xor ( n14759 , n14758 , n11710 );
xor ( n14760 , n10054 , n7782 );
xor ( n14761 , n14760 , n7804 );
not ( n14762 , n14761 );
xor ( n14763 , n10596 , n7632 );
xor ( n14764 , n14763 , n7654 );
and ( n14765 , n14762 , n14764 );
xor ( n14766 , n14759 , n14765 );
xor ( n14767 , n14757 , n14766 );
xor ( n14768 , n14722 , n14767 );
xor ( n14769 , n6691 , n11993 );
xor ( n14770 , n14769 , n10055 );
xor ( n14771 , n11340 , n10349 );
xor ( n14772 , n14771 , n7319 );
not ( n14773 , n14772 );
xor ( n14774 , n8229 , n12371 );
xor ( n14775 , n14774 , n13225 );
and ( n14776 , n14773 , n14775 );
xor ( n14777 , n14770 , n14776 );
xor ( n14778 , n9773 , n11436 );
xor ( n14779 , n14778 , n11560 );
xor ( n14780 , n12776 , n9699 );
xor ( n14781 , n14780 , n9362 );
not ( n14782 , n14781 );
xor ( n14783 , n13683 , n9455 );
xor ( n14784 , n14783 , n11786 );
and ( n14785 , n14782 , n14784 );
xor ( n14786 , n14779 , n14785 );
xor ( n14787 , n14777 , n14786 );
xor ( n14788 , n10042 , n7782 );
xor ( n14789 , n14788 , n7804 );
xor ( n14790 , n7974 , n7828 );
xor ( n14791 , n14790 , n7851 );
not ( n14792 , n14791 );
xor ( n14793 , n9104 , n10142 );
xor ( n14794 , n14793 , n6659 );
and ( n14795 , n14792 , n14794 );
xor ( n14796 , n14789 , n14795 );
xor ( n14797 , n14787 , n14796 );
xor ( n14798 , n7729 , n9428 );
not ( n14799 , n6583 );
buf ( n14800 , n6566 );
and ( n14801 , n14799 , n14800 );
buf ( n14802 , n6567 );
xor ( n14803 , n14802 , n14800 );
and ( n14804 , n14803 , n6583 );
or ( n14805 , n14801 , n14804 );
xor ( n14806 , n14805 , n14679 );
buf ( n14807 , n6568 );
xor ( n14808 , n14806 , n14807 );
buf ( n14809 , n6569 );
xor ( n14810 , n14808 , n14809 );
buf ( n14811 , n6570 );
xor ( n14812 , n14810 , n14811 );
xor ( n14813 , n14798 , n14812 );
xor ( n14814 , n7572 , n14408 );
xor ( n14815 , n14814 , n13616 );
not ( n14816 , n14815 );
xor ( n14817 , n9967 , n14051 );
xor ( n14818 , n14817 , n12931 );
and ( n14819 , n14816 , n14818 );
xor ( n14820 , n14813 , n14819 );
xor ( n14821 , n14797 , n14820 );
xor ( n14822 , n8713 , n11410 );
xor ( n14823 , n14822 , n7710 );
xor ( n14824 , n8967 , n12125 );
xor ( n14825 , n14824 , n8036 );
not ( n14826 , n14825 );
xor ( n14827 , n13038 , n9855 );
xor ( n14828 , n14827 , n9877 );
and ( n14829 , n14826 , n14828 );
xor ( n14830 , n14823 , n14829 );
xor ( n14831 , n14821 , n14830 );
xor ( n14832 , n14768 , n14831 );
not ( n14833 , n14832 );
xor ( n14834 , n10419 , n13996 );
not ( n14835 , n6583 );
buf ( n14836 , n6571 );
and ( n14837 , n14835 , n14836 );
buf ( n14838 , n6572 );
xor ( n14839 , n14838 , n14836 );
and ( n14840 , n14839 , n6583 );
or ( n14841 , n14837 , n14840 );
xor ( n14842 , n14841 , n14355 );
buf ( n14843 , n6573 );
xor ( n14844 , n14842 , n14843 );
buf ( n14845 , n6574 );
xor ( n14846 , n14844 , n14845 );
xor ( n14847 , n14846 , n8911 );
xor ( n14848 , n14834 , n14847 );
xor ( n14849 , n11211 , n12647 );
xor ( n14850 , n14849 , n12662 );
not ( n14851 , n14850 );
and ( n14852 , n14851 , n12219 );
xor ( n14853 , n14848 , n14852 );
xor ( n14854 , n11878 , n8948 );
xor ( n14855 , n14854 , n9972 );
not ( n14856 , n14855 );
xor ( n14857 , n9526 , n11386 );
xor ( n14858 , n14857 , n12756 );
and ( n14859 , n14856 , n14858 );
xor ( n14860 , n12084 , n14859 );
xor ( n14861 , n13076 , n7600 );
xor ( n14862 , n14861 , n8653 );
not ( n14863 , n14862 );
xor ( n14864 , n11554 , n10776 );
xor ( n14865 , n14864 , n10797 );
and ( n14866 , n14863 , n14865 );
xor ( n14867 , n12129 , n14866 );
xor ( n14868 , n14860 , n14867 );
xor ( n14869 , n9958 , n14051 );
xor ( n14870 , n14869 , n12931 );
not ( n14871 , n14870 );
xor ( n14872 , n9935 , n9200 );
xor ( n14873 , n14872 , n13188 );
and ( n14874 , n14871 , n14873 );
xor ( n14875 , n12166 , n14874 );
xor ( n14876 , n14868 , n14875 );
xor ( n14877 , n14401 , n11050 );
xor ( n14878 , n14877 , n11072 );
not ( n14879 , n14878 );
xor ( n14880 , n13240 , n10366 );
xor ( n14881 , n14880 , n10388 );
and ( n14882 , n14879 , n14881 );
xor ( n14883 , n12214 , n14882 );
xor ( n14884 , n14876 , n14883 );
not ( n14885 , n14848 );
and ( n14886 , n14885 , n14850 );
xor ( n14887 , n12239 , n14886 );
xor ( n14888 , n14884 , n14887 );
xor ( n14889 , n14853 , n14888 );
xor ( n14890 , n9039 , n12102 );
xor ( n14891 , n14890 , n12125 );
xor ( n14892 , n11270 , n9533 );
xor ( n14893 , n14892 , n8018 );
not ( n14894 , n14893 );
xor ( n14895 , n9137 , n12804 );
xor ( n14896 , n14895 , n7926 );
and ( n14897 , n14894 , n14896 );
xor ( n14898 , n14891 , n14897 );
xor ( n14899 , n9710 , n7886 );
xor ( n14900 , n14899 , n7908 );
xor ( n14901 , n9734 , n7469 );
xor ( n14902 , n14901 , n11147 );
not ( n14903 , n14902 );
xor ( n14904 , n6816 , n7073 );
xor ( n14905 , n14904 , n7095 );
and ( n14906 , n14903 , n14905 );
xor ( n14907 , n14900 , n14906 );
xor ( n14908 , n14898 , n14907 );
xor ( n14909 , n7670 , n8105 );
xor ( n14910 , n14909 , n6615 );
xor ( n14911 , n7423 , n6871 );
xor ( n14912 , n14911 , n14408 );
not ( n14913 , n14912 );
xor ( n14914 , n8267 , n9244 );
xor ( n14915 , n14914 , n10166 );
and ( n14916 , n14913 , n14915 );
xor ( n14917 , n14910 , n14916 );
xor ( n14918 , n14908 , n14917 );
xor ( n14919 , n11307 , n7335 );
xor ( n14920 , n14919 , n10098 );
xor ( n14921 , n8678 , n9307 );
xor ( n14922 , n14921 , n13507 );
not ( n14923 , n14922 );
xor ( n14924 , n10139 , n13020 );
xor ( n14925 , n14924 , n9583 );
and ( n14926 , n14923 , n14925 );
xor ( n14927 , n14920 , n14926 );
xor ( n14928 , n14918 , n14927 );
xor ( n14929 , n11732 , n6727 );
xor ( n14930 , n14929 , n12213 );
xor ( n14931 , n12851 , n12292 );
xor ( n14932 , n14931 , n14082 );
not ( n14933 , n14932 );
xor ( n14934 , n9490 , n8505 );
xor ( n14935 , n14934 , n7267 );
and ( n14936 , n14933 , n14935 );
xor ( n14937 , n14930 , n14936 );
xor ( n14938 , n14928 , n14937 );
xor ( n14939 , n14889 , n14938 );
and ( n14940 , n14833 , n14939 );
xor ( n14941 , n14713 , n14940 );
and ( n14942 , n14941 , n6584 );
or ( n14943 , n14708 , n14942 );
and ( n14944 , n14706 , n14943 );
buf ( n14945 , n14944 );
buf ( n14946 , n14945 );
not ( n14947 , n6578 );
not ( n14948 , n6584 );
and ( n14949 , n14948 , n12974 );
xor ( n14950 , n9654 , n8167 );
xor ( n14951 , n14950 , n8189 );
xor ( n14952 , n10862 , n13104 );
xor ( n14953 , n14952 , n9178 );
not ( n14954 , n14953 );
xor ( n14955 , n12489 , n8635 );
xor ( n14956 , n14955 , n8705 );
and ( n14957 , n14954 , n14956 );
xor ( n14958 , n14951 , n14957 );
xor ( n14959 , n11799 , n9511 );
xor ( n14960 , n14959 , n9533 );
xor ( n14961 , n11583 , n9161 );
xor ( n14962 , n14961 , n9560 );
not ( n14963 , n14962 );
xor ( n14964 , n12800 , n8886 );
xor ( n14965 , n14964 , n8908 );
and ( n14966 , n14963 , n14965 );
xor ( n14967 , n14960 , n14966 );
xor ( n14968 , n13182 , n7677 );
xor ( n14969 , n14968 , n7686 );
xor ( n14970 , n7022 , n14847 );
xor ( n14971 , n14970 , n11892 );
not ( n14972 , n14971 );
xor ( n14973 , n7068 , n13358 );
xor ( n14974 , n14973 , n13378 );
and ( n14975 , n14972 , n14974 );
xor ( n14976 , n14969 , n14975 );
xor ( n14977 , n14967 , n14976 );
xor ( n14978 , n9519 , n11386 );
xor ( n14979 , n14978 , n12756 );
not ( n14980 , n14951 );
and ( n14981 , n14980 , n14953 );
xor ( n14982 , n14979 , n14981 );
xor ( n14983 , n14977 , n14982 );
xor ( n14984 , n8075 , n11169 );
xor ( n14985 , n14984 , n8318 );
xor ( n14986 , n10908 , n12999 );
xor ( n14987 , n14986 , n13020 );
not ( n14988 , n14987 );
xor ( n14989 , n11405 , n13960 );
xor ( n14990 , n14989 , n11978 );
and ( n14991 , n14988 , n14990 );
xor ( n14992 , n14985 , n14991 );
xor ( n14993 , n14983 , n14992 );
xor ( n14994 , n10020 , n14128 );
xor ( n14995 , n14994 , n12721 );
xor ( n14996 , n10320 , n8234 );
xor ( n14997 , n14996 , n8250 );
not ( n14998 , n14997 );
xor ( n14999 , n7732 , n9428 );
xor ( n15000 , n14999 , n14812 );
and ( n15001 , n14998 , n15000 );
xor ( n15002 , n14995 , n15001 );
xor ( n15003 , n14993 , n15002 );
xor ( n15004 , n14958 , n15003 );
xor ( n15005 , n9064 , n11590 );
xor ( n15006 , n15005 , n11604 );
xor ( n15007 , n6984 , n11907 );
xor ( n15008 , n15007 , n11866 );
not ( n15009 , n15008 );
xor ( n15010 , n9454 , n10497 );
xor ( n15011 , n15010 , n13714 );
and ( n15012 , n15009 , n15011 );
xor ( n15013 , n15006 , n15012 );
xor ( n15014 , n7211 , n8036 );
xor ( n15015 , n15014 , n8058 );
xor ( n15016 , n7403 , n6849 );
xor ( n15017 , n15016 , n6871 );
not ( n15018 , n15017 );
xor ( n15019 , n10033 , n14128 );
xor ( n15020 , n15019 , n12721 );
and ( n15021 , n15018 , n15020 );
xor ( n15022 , n15015 , n15021 );
xor ( n15023 , n15013 , n15022 );
xor ( n15024 , n8601 , n9761 );
xor ( n15025 , n15024 , n8083 );
xor ( n15026 , n10305 , n7147 );
xor ( n15027 , n15026 , n13960 );
not ( n15028 , n15027 );
xor ( n15029 , n10697 , n7996 );
xor ( n15030 , n15029 , n10192 );
and ( n15031 , n15028 , n15030 );
xor ( n15032 , n15025 , n15031 );
xor ( n15033 , n15023 , n15032 );
xor ( n15034 , n11679 , n12473 );
xor ( n15035 , n15034 , n12647 );
xor ( n15036 , n9806 , n11786 );
xor ( n15037 , n15036 , n12521 );
not ( n15038 , n15037 );
xor ( n15039 , n11291 , n7319 );
xor ( n15040 , n15039 , n7335 );
and ( n15041 , n15038 , n15040 );
xor ( n15042 , n15035 , n15041 );
xor ( n15043 , n15033 , n15042 );
xor ( n15044 , n13277 , n9787 );
xor ( n15045 , n15044 , n11850 );
xor ( n15046 , n10795 , n9715 );
xor ( n15047 , n15046 , n8886 );
not ( n15048 , n15047 );
xor ( n15049 , n6818 , n7073 );
xor ( n15050 , n15049 , n7095 );
and ( n15051 , n15048 , n15050 );
xor ( n15052 , n15045 , n15051 );
xor ( n15053 , n15043 , n15052 );
xor ( n15054 , n15004 , n15053 );
xor ( n15055 , n10723 , n13687 );
xor ( n15056 , n15055 , n9809 );
xor ( n15057 , n8929 , n10192 );
xor ( n15058 , n15057 , n14029 );
not ( n15059 , n15058 );
and ( n15060 , n15059 , n13581 );
xor ( n15061 , n15056 , n15060 );
not ( n15062 , n13471 );
xor ( n15063 , n8603 , n9761 );
xor ( n15064 , n15063 , n8083 );
and ( n15065 , n15062 , n15064 );
xor ( n15066 , n13468 , n15065 );
xor ( n15067 , n10817 , n12492 );
xor ( n15068 , n15067 , n7632 );
not ( n15069 , n15068 );
xor ( n15070 , n13327 , n13149 );
xor ( n15071 , n15070 , n13169 );
and ( n15072 , n15069 , n15071 );
xor ( n15073 , n13512 , n15072 );
xor ( n15074 , n15066 , n15073 );
xor ( n15075 , n9239 , n6947 );
xor ( n15076 , n15075 , n6963 );
not ( n15077 , n15076 );
xor ( n15078 , n12659 , n11739 );
xor ( n15079 , n15078 , n11761 );
and ( n15080 , n15077 , n15079 );
xor ( n15081 , n13562 , n15080 );
xor ( n15082 , n15074 , n15081 );
not ( n15083 , n15056 );
and ( n15084 , n15083 , n15058 );
xor ( n15085 , n13586 , n15084 );
xor ( n15086 , n15082 , n15085 );
xor ( n15087 , n7921 , n8908 );
xor ( n15088 , n15087 , n10642 );
not ( n15089 , n15088 );
xor ( n15090 , n6846 , n8807 );
xor ( n15091 , n15090 , n8822 );
and ( n15092 , n15089 , n15091 );
xor ( n15093 , n13596 , n15092 );
xor ( n15094 , n15086 , n15093 );
xor ( n15095 , n15061 , n15094 );
xor ( n15096 , n7028 , n14847 );
xor ( n15097 , n15096 , n11892 );
not ( n15098 , n15097 );
xor ( n15099 , n13524 , n7533 );
xor ( n15100 , n15099 , n7555 );
and ( n15101 , n15098 , n15100 );
xor ( n15102 , n13642 , n15101 );
xor ( n15103 , n12124 , n6819 );
xor ( n15104 , n15103 , n12347 );
not ( n15105 , n15104 );
xor ( n15106 , n8374 , n9384 );
xor ( n15107 , n15106 , n10530 );
and ( n15108 , n15105 , n15107 );
xor ( n15109 , n13658 , n15108 );
xor ( n15110 , n15102 , n15109 );
xor ( n15111 , n7515 , n9615 );
xor ( n15112 , n15111 , n8584 );
not ( n15113 , n15112 );
xor ( n15114 , n7541 , n8127 );
xor ( n15115 , n15114 , n8142 );
and ( n15116 , n15113 , n15115 );
xor ( n15117 , n13688 , n15116 );
xor ( n15118 , n15110 , n15117 );
xor ( n15119 , n9477 , n10034 );
xor ( n15120 , n15119 , n8505 );
not ( n15121 , n15120 );
xor ( n15122 , n14644 , n14444 );
xor ( n15123 , n15122 , n12393 );
and ( n15124 , n15121 , n15123 );
xor ( n15125 , n13740 , n15124 );
xor ( n15126 , n15118 , n15125 );
xor ( n15127 , n7124 , n10822 );
xor ( n15128 , n15127 , n10603 );
not ( n15129 , n15128 );
xor ( n15130 , n7081 , n13378 );
xor ( n15131 , n15130 , n13774 );
and ( n15132 , n15129 , n15131 );
xor ( n15133 , n13750 , n15132 );
xor ( n15134 , n15126 , n15133 );
xor ( n15135 , n15095 , n15134 );
not ( n15136 , n15135 );
xor ( n15137 , n7006 , n11866 );
xor ( n15138 , n15137 , n10845 );
xor ( n15139 , n13067 , n7579 );
xor ( n15140 , n15139 , n7600 );
not ( n15141 , n15140 );
and ( n15142 , n15141 , n14005 );
xor ( n15143 , n15138 , n15142 );
xor ( n15144 , n8971 , n12125 );
xor ( n15145 , n15144 , n8036 );
not ( n15146 , n15145 );
xor ( n15147 , n11512 , n10120 );
xor ( n15148 , n15147 , n10012 );
and ( n15149 , n15146 , n15148 );
xor ( n15150 , n13928 , n15149 );
xor ( n15151 , n9197 , n13652 );
xor ( n15152 , n15151 , n7677 );
not ( n15153 , n15152 );
xor ( n15154 , n12803 , n8886 );
xor ( n15155 , n15154 , n8908 );
and ( n15156 , n15153 , n15155 );
xor ( n15157 , n13937 , n15156 );
xor ( n15158 , n15150 , n15157 );
not ( n15159 , n13919 );
xor ( n15160 , n11804 , n9511 );
xor ( n15161 , n15160 , n9533 );
and ( n15162 , n15159 , n15161 );
xor ( n15163 , n13916 , n15162 );
xor ( n15164 , n15158 , n15163 );
xor ( n15165 , n13576 , n12696 );
xor ( n15166 , n15165 , n9478 );
not ( n15167 , n15166 );
xor ( n15168 , n9582 , n8552 );
xor ( n15169 , n15168 , n7737 );
and ( n15170 , n15167 , n15169 );
xor ( n15171 , n14000 , n15170 );
xor ( n15172 , n15164 , n15171 );
not ( n15173 , n15138 );
and ( n15174 , n15173 , n15140 );
xor ( n15175 , n14052 , n15174 );
xor ( n15176 , n15172 , n15175 );
xor ( n15177 , n15143 , n15176 );
xor ( n15178 , n7354 , n12160 );
xor ( n15179 , n15178 , n13068 );
not ( n15180 , n15179 );
xor ( n15181 , n9193 , n13652 );
xor ( n15182 , n15181 , n7677 );
and ( n15183 , n15180 , n15182 );
xor ( n15184 , n14083 , n15183 );
xor ( n15185 , n7696 , n11978 );
xor ( n15186 , n15185 , n11993 );
not ( n15187 , n15186 );
xor ( n15188 , n13352 , n8974 );
xor ( n15189 , n15188 , n7216 );
and ( n15190 , n15187 , n15189 );
xor ( n15191 , n14092 , n15190 );
xor ( n15192 , n15184 , n15191 );
xor ( n15193 , n13056 , n7579 );
xor ( n15194 , n15193 , n7600 );
not ( n15195 , n15194 );
xor ( n15196 , n8750 , n11710 );
xor ( n15197 , n15196 , n8460 );
and ( n15198 , n15195 , n15197 );
xor ( n15199 , n14102 , n15198 );
xor ( n15200 , n15192 , n15199 );
xor ( n15201 , n10611 , n7654 );
xor ( n15202 , n15201 , n12473 );
not ( n15203 , n15202 );
xor ( n15204 , n10692 , n7996 );
xor ( n15205 , n15204 , n10192 );
and ( n15206 , n15203 , n15205 );
xor ( n15207 , n14133 , n15206 );
xor ( n15208 , n15200 , n15207 );
xor ( n15209 , n9546 , n7948 );
xor ( n15210 , n15209 , n11650 );
not ( n15211 , n15210 );
xor ( n15212 , n9576 , n8552 );
xor ( n15213 , n15212 , n7737 );
and ( n15214 , n15211 , n15213 );
xor ( n15215 , n14144 , n15214 );
xor ( n15216 , n15208 , n15215 );
xor ( n15217 , n15177 , n15216 );
and ( n15218 , n15136 , n15217 );
xor ( n15219 , n15054 , n15218 );
and ( n15220 , n15219 , n6584 );
or ( n15221 , n14949 , n15220 );
and ( n15222 , n14947 , n15221 );
buf ( n15223 , n15222 );
buf ( n15224 , n15223 );
not ( n15225 , n6578 );
not ( n15226 , n6584 );
and ( n15227 , n15226 , n8165 );
xor ( n15228 , n10941 , n10797 );
xor ( n15229 , n15228 , n12804 );
xor ( n15230 , n7172 , n10388 );
xor ( n15231 , n15230 , n12015 );
not ( n15232 , n15231 );
xor ( n15233 , n10853 , n13104 );
xor ( n15234 , n15233 , n9178 );
and ( n15235 , n15232 , n15234 );
xor ( n15236 , n15229 , n15235 );
xor ( n15237 , n11431 , n7759 );
xor ( n15238 , n15237 , n10776 );
xor ( n15239 , n11471 , n7980 );
xor ( n15240 , n15239 , n7996 );
not ( n15241 , n15240 );
xor ( n15242 , n13822 , n7710 );
xor ( n15243 , n15242 , n6705 );
and ( n15244 , n15241 , n15243 );
xor ( n15245 , n15238 , n15244 );
xor ( n15246 , n11801 , n9511 );
xor ( n15247 , n15246 , n9533 );
not ( n15248 , n15229 );
and ( n15249 , n15248 , n15231 );
xor ( n15250 , n15247 , n15249 );
xor ( n15251 , n15245 , n15250 );
xor ( n15252 , n6982 , n11907 );
xor ( n15253 , n15252 , n11866 );
xor ( n15254 , n8989 , n13774 );
xor ( n15255 , n15254 , n13537 );
not ( n15256 , n15255 );
xor ( n15257 , n13686 , n9455 );
xor ( n15258 , n15257 , n11786 );
and ( n15259 , n15256 , n15258 );
xor ( n15260 , n15253 , n15259 );
xor ( n15261 , n15251 , n15260 );
xor ( n15262 , n7550 , n8127 );
xor ( n15263 , n15262 , n8142 );
xor ( n15264 , n12644 , n12954 );
xor ( n15265 , n15264 , n11739 );
not ( n15266 , n15265 );
xor ( n15267 , n12572 , n8757 );
xor ( n15268 , n15267 , n8766 );
and ( n15269 , n15266 , n15268 );
xor ( n15270 , n15263 , n15269 );
xor ( n15271 , n15261 , n15270 );
xor ( n15272 , n12995 , n8789 );
xor ( n15273 , n15272 , n8530 );
xor ( n15274 , n8838 , n6659 );
xor ( n15275 , n15274 , n6681 );
not ( n15276 , n15275 );
xor ( n15277 , n6895 , n9493 );
not ( n15278 , n6583 );
buf ( n15279 , n6575 );
and ( n15280 , n15278 , n15279 );
buf ( n15281 , n6576 );
xor ( n15282 , n15281 , n15279 );
and ( n15283 , n15282 , n6583 );
or ( n15284 , n15280 , n15283 );
xor ( n15285 , n7246 , n15284 );
xor ( n15286 , n15285 , n12043 );
xor ( n15287 , n15286 , n13386 );
xor ( n15288 , n15287 , n14598 );
xor ( n15289 , n15277 , n15288 );
and ( n15290 , n15276 , n15289 );
xor ( n15291 , n15273 , n15290 );
xor ( n15292 , n15271 , n15291 );
xor ( n15293 , n15236 , n15292 );
xor ( n15294 , n11992 , n11218 );
xor ( n15295 , n15294 , n7782 );
xor ( n15296 , n14069 , n12234 );
xor ( n15297 , n15296 , n6896 );
not ( n15298 , n15297 );
xor ( n15299 , n10937 , n10797 );
xor ( n15300 , n15299 , n12804 );
and ( n15301 , n15298 , n15300 );
xor ( n15302 , n15295 , n15301 );
xor ( n15303 , n11496 , n10098 );
xor ( n15304 , n15303 , n10120 );
xor ( n15305 , n8592 , n9761 );
xor ( n15306 , n15305 , n8083 );
not ( n15307 , n15306 );
xor ( n15308 , n13969 , n11474 );
xor ( n15309 , n15308 , n10698 );
and ( n15310 , n15307 , n15309 );
xor ( n15311 , n15304 , n15310 );
xor ( n15312 , n15302 , n15311 );
xor ( n15313 , n13713 , n12323 );
xor ( n15314 , n15313 , n11459 );
xor ( n15315 , n6882 , n9493 );
xor ( n15316 , n15315 , n15288 );
not ( n15317 , n15316 );
xor ( n15318 , n7088 , n13378 );
xor ( n15319 , n15318 , n13774 );
and ( n15320 , n15317 , n15319 );
xor ( n15321 , n15314 , n15320 );
xor ( n15322 , n15312 , n15321 );
xor ( n15323 , n8459 , n12978 );
xor ( n15324 , n15323 , n11325 );
xor ( n15325 , n7460 , n10867 );
xor ( n15326 , n15325 , n9920 );
not ( n15327 , n15326 );
xor ( n15328 , n12387 , n10260 );
xor ( n15329 , n15328 , n10282 );
and ( n15330 , n15327 , n15329 );
xor ( n15331 , n15324 , n15330 );
xor ( n15332 , n15322 , n15331 );
xor ( n15333 , n7266 , n11805 );
xor ( n15334 , n15333 , n11275 );
xor ( n15335 , n12833 , n9340 );
xor ( n15336 , n15335 , n12292 );
not ( n15337 , n15336 );
xor ( n15338 , n12567 , n8757 );
xor ( n15339 , n15338 , n8766 );
and ( n15340 , n15337 , n15339 );
xor ( n15341 , n15334 , n15340 );
xor ( n15342 , n15332 , n15341 );
xor ( n15343 , n15293 , n15342 );
xor ( n15344 , n9492 , n8505 );
xor ( n15345 , n15344 , n7267 );
xor ( n15346 , n7399 , n6849 );
xor ( n15347 , n15346 , n6871 );
not ( n15348 , n15347 );
xor ( n15349 , n13163 , n12433 );
xor ( n15350 , n15349 , n12447 );
and ( n15351 , n15348 , n15350 );
xor ( n15352 , n15345 , n15351 );
xor ( n15353 , n8015 , n12756 );
xor ( n15354 , n15353 , n13358 );
xor ( n15355 , n7188 , n12015 );
xor ( n15356 , n15355 , n12037 );
not ( n15357 , n15356 );
xor ( n15358 , n10628 , n9085 );
xor ( n15359 , n15358 , n7406 );
and ( n15360 , n15357 , n15359 );
xor ( n15361 , n15354 , n15360 );
xor ( n15362 , n11145 , n9920 );
xor ( n15363 , n15362 , n9942 );
xor ( n15364 , n12064 , n10944 );
xor ( n15365 , n15364 , n9140 );
not ( n15366 , n15365 );
xor ( n15367 , n7133 , n10603 );
xor ( n15368 , n15367 , n10619 );
and ( n15369 , n15366 , n15368 );
xor ( n15370 , n15363 , n15369 );
xor ( n15371 , n15361 , n15370 );
xor ( n15372 , n8425 , n12573 );
xor ( n15373 , n15372 , n14258 );
not ( n15374 , n15345 );
and ( n15375 , n15374 , n15347 );
xor ( n15376 , n15373 , n15375 );
xor ( n15377 , n15371 , n15376 );
xor ( n15378 , n12837 , n9340 );
xor ( n15379 , n15378 , n12292 );
xor ( n15380 , n9108 , n10142 );
xor ( n15381 , n15380 , n6659 );
not ( n15382 , n15381 );
xor ( n15383 , n12484 , n8635 );
xor ( n15384 , n15383 , n8705 );
and ( n15385 , n15382 , n15384 );
xor ( n15386 , n15379 , n15385 );
xor ( n15387 , n15377 , n15386 );
xor ( n15388 , n14048 , n14334 );
xor ( n15389 , n15388 , n10584 );
xor ( n15390 , n8821 , n7368 );
xor ( n15391 , n15390 , n7390 );
not ( n15392 , n15391 );
xor ( n15393 , n12798 , n8886 );
xor ( n15394 , n15393 , n8908 );
and ( n15395 , n15392 , n15394 );
xor ( n15396 , n15389 , n15395 );
xor ( n15397 , n15387 , n15396 );
xor ( n15398 , n15352 , n15397 );
xor ( n15399 , n15398 , n14055 );
not ( n15400 , n15399 );
not ( n15401 , n15205 );
and ( n15402 , n15401 , n14107 );
xor ( n15403 , n15202 , n15402 );
xor ( n15404 , n15403 , n15216 );
xor ( n15405 , n15404 , n13287 );
and ( n15406 , n15400 , n15405 );
xor ( n15407 , n15343 , n15406 );
and ( n15408 , n15407 , n6584 );
or ( n15409 , n15227 , n15408 );
and ( n15410 , n15225 , n15409 );
buf ( n15411 , n15410 );
buf ( n15412 , n15411 );
endmodule

