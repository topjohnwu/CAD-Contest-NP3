//
// Conformal-LEC Version 16.10-d005 ( 21-Apr-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 ;
output n2048 , n2049 ;

wire n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , 
     n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , 
     n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , 
     n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , 
     n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , 
     n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , 
     n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , 
     n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , 
     n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , 
     n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , 
     n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , 
     n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , 
     n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , 
     n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , 
     n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , 
     n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , 
     n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , 
     n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , 
     n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , 
     n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , 
     n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , 
     n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , 
     n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , 
     n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , 
     n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , 
     n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , 
     n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , 
     n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , 
     n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , 
     n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , 
     n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , 
     n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , 
     n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , 
     n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , 
     n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , 
     n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , 
     n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , 
     n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , 
     n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , 
     n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , 
     n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , 
     n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , 
     n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , 
     n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , 
     n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , 
     n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , 
     n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , 
     n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , 
     n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , 
     n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , 
     n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , 
     n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , 
     n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , 
     n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , 
     n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , 
     n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , 
     n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , 
     n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , 
     n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , 
     n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , 
     n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , 
     n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , 
     n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , 
     n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , 
     n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , 
     n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , 
     n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , 
     n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , 
     n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , 
     n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , 
     n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , 
     n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , 
     n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , 
     n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , 
     n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , 
     n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , 
     n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , 
     n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , 
     n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , 
     n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , 
     n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , 
     n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , 
     n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , 
     n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , 
     n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , 
     n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , 
     n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , 
     n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , 
     n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , 
     n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , 
     n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , 
     n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , 
     n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , 
     n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , 
     n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , 
     n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , 
     n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , 
     n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , 
     n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , 
     n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , 
     n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , 
     n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , 
     n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , 
     n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , 
     n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , 
     n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , 
     n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , 
     n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , 
     n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , 
     n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , 
     n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , 
     n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , 
     n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , 
     n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , 
     n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , 
     n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , 
     n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , 
     n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , 
     n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , 
     n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , 
     n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , 
     n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , 
     n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , 
     n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , 
     n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , 
     n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , 
     n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , 
     n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , 
     n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , 
     n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , 
     n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , 
     n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , 
     n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , 
     n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , 
     n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , 
     n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , 
     n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , 
     n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , 
     n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , 
     n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , 
     n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , 
     n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , 
     n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , 
     n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , 
     n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , 
     n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , 
     n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , 
     n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , 
     n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , 
     n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , 
     n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , 
     n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , 
     n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , 
     n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , 
     n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , 
     n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , 
     n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , 
     n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , 
     n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , 
     n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , 
     n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , 
     n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , 
     n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , 
     n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , 
     n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , 
     n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , 
     n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , 
     n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , 
     n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , 
     n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , 
     n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , 
     n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , 
     n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , 
     n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , 
     n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , 
     n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , 
     n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , 
     n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , 
     n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , 
     n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , 
     n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , 
     n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , 
     n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , 
     n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , 
     n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , 
     n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , 
     n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , 
     n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , 
     n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , 
     n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , 
     n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , 
     n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , 
     n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , 
     n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , 
     n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , 
     n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , 
     n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , 
     n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , 
     n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , 
     n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , 
     n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , 
     n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , 
     n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , 
     n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , 
     n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , 
     n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , 
     n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , 
     n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , 
     n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , 
     n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , 
     n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , 
     n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , 
     n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , 
     n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , 
     n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , 
     n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , 
     n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , 
     n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , 
     n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , 
     n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , 
     n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , 
     n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , 
     n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , 
     n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , 
     n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , 
     n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , 
     n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , 
     n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , 
     n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , 
     n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , 
     n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , 
     n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , 
     n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , 
     n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , 
     n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , 
     n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , 
     n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , 
     n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , 
     n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , 
     n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , 
     n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , 
     n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , 
     n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , 
     n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , 
     n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , 
     n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , 
     n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , 
     n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , 
     n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , 
     n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , 
     n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , 
     n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , 
     n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , 
     n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , 
     n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , 
     n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , 
     n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , 
     n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , 
     n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , 
     n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , 
     n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , 
     n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , 
     n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , 
     n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , 
     n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , 
     n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , 
     n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , 
     n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , 
     n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , 
     n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , 
     n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , 
     n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , 
     n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , 
     n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , 
     n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , 
     n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , 
     n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , 
     n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , 
     n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , 
     n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , 
     n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , 
     n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , 
     n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , 
     n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , 
     n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , 
     n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , 
     n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , 
     n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , 
     n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , 
     n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , 
     n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , 
     n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , 
     n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , 
     n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , 
     n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , 
     n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , 
     n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , 
     n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , 
     n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , 
     n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , 
     n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , 
     n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , 
     n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , 
     n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , 
     n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , 
     n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , 
     n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , 
     n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , 
     n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , 
     n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , 
     n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , 
     n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , 
     n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , 
     n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , 
     n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , 
     n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , 
     n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , 
     n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , 
     n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , 
     n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , 
     n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , 
     n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , 
     n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , 
     n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , 
     n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , 
     n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , 
     n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , 
     n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , 
     n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , 
     n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , 
     n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , 
     n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , 
     n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , 
     n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , 
     n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , 
     n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , 
     n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , 
     n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , 
     n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , 
     n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , 
     n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , 
     n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , 
     n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , 
     n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , 
     n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , 
     n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , 
     n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , 
     n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , 
     n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , 
     n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , 
     n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , 
     n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , 
     n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , 
     n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , 
     n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , 
     n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , 
     n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , 
     n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , 
     n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , 
     n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , 
     n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , 
     n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , 
     n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , 
     n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , 
     n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , 
     n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , 
     n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , 
     n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , 
     n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , 
     n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , 
     n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , 
     n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , 
     n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , 
     n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , 
     n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , 
     n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , 
     n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , 
     n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , 
     n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , 
     n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , 
     n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , 
     n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , 
     n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , 
     n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , 
     n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , 
     n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , 
     n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , 
     n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , 
     n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , 
     n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , 
     n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , 
     n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , 
     n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , 
     n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , 
     n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , 
     n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , 
     n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , 
     n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , 
     n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , 
     n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , 
     n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , 
     n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , 
     n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , 
     n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , 
     n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , 
     n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , 
     n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , 
     n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , 
     n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , 
     n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , 
     n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , 
     n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , 
     n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , 
     n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , 
     n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , 
     n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , 
     n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , 
     n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , 
     n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , 
     n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , 
     n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , 
     n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , 
     n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , 
     n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , 
     n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , 
     n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , 
     n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , 
     n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , 
     n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , 
     n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , 
     n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , 
     n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , 
     n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , 
     n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , 
     n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , 
     n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , 
     n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , 
     n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , 
     n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , 
     n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , 
     n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , 
     n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , 
     n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , 
     n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , 
     n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , 
     n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , 
     n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , 
     n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , 
     n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , 
     n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , 
     n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , 
     n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , 
     n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , 
     n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , 
     n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , 
     n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , 
     n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , 
     n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , 
     n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , 
     n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , 
     n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , 
     n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , 
     n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , 
     n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , 
     n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , 
     n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , 
     n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , 
     n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , 
     n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , 
     n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , 
     n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , 
     n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , 
     n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , 
     n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , 
     n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , 
     n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , 
     n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , 
     n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , 
     n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , 
     n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , 
     n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , 
     n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , 
     n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , 
     n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , 
     n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , 
     n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , 
     n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , 
     n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , 
     n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , 
     n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , 
     n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , 
     n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , 
     n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , 
     n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , 
     n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , 
     n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , 
     n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , 
     n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , 
     n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , 
     n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , 
     n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , 
     n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , 
     n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , 
     n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , 
     n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , 
     n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , 
     n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , 
     n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , 
     n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , 
     n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , 
     n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , 
     n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , 
     n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , 
     n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , 
     n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , 
     n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , 
     n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , 
     n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , 
     n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , 
     n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , 
     n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , 
     n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , 
     n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , 
     n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , 
     n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , 
     n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , 
     n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , 
     n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , 
     n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , 
     n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , 
     n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , 
     n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , 
     n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , 
     n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , 
     n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , 
     n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , 
     n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , 
     n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , 
     n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , 
     n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , 
     n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , 
     n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , 
     n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , 
     n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , 
     n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , 
     n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , 
     n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , 
     n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , 
     n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , 
     n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , 
     n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , 
     n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , 
     n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , 
     n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , 
     n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , 
     n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , 
     n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , 
     n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , 
     n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , 
     n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , 
     n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , 
     n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , 
     n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , 
     n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , 
     n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , 
     n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , 
     n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , 
     n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , 
     n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , 
     n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , 
     n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , 
     n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , 
     n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , 
     n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , 
     n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , 
     n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , 
     n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , 
     n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , 
     n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , 
     n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , 
     n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , 
     n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , 
     n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , 
     n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , 
     n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , 
     n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , 
     n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , 
     n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , 
     n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , 
     n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , 
     n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , 
     n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , 
     n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , 
     n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , 
     n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , 
     n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , 
     n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , 
     n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , 
     n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , 
     n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , 
     n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , 
     n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , 
     n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , 
     n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , 
     n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , 
     n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , 
     n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , 
     n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , 
     n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , 
     n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , 
     n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , 
     n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , 
     n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , 
     n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , 
     n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , 
     n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , 
     n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , 
     n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , 
     n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , 
     n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , 
     n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , 
     n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , 
     n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , 
     n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , 
     n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , 
     n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , 
     n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , 
     n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , 
     n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , 
     n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , 
     n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , 
     n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , 
     n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , 
     n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , 
     n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , 
     n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , 
     n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , 
     n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , 
     n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , 
     n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , 
     n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , 
     n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , 
     n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , 
     n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , 
     n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , 
     n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , 
     n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , 
     n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , 
     n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , 
     n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , 
     n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , 
     n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , 
     n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , 
     n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , 
     n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , 
     n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , 
     n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , 
     n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , 
     n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , 
     n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , 
     n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , 
     n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , 
     n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , 
     n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , 
     n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , 
     n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , 
     n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , 
     n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , 
     n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , 
     n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , 
     n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , 
     n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , 
     n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , 
     n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , 
     n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , 
     n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , 
     n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , 
     n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , 
     n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , 
     n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , 
     n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , 
     n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , 
     n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , 
     n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , 
     n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , 
     n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , 
     n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , 
     n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , 
     n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , 
     n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , 
     n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , 
     n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , 
     n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , 
     n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , 
     n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , 
     n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , 
     n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , 
     n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , 
     n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , 
     n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , 
     n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , 
     n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , 
     n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , 
     n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , 
     n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , 
     n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , 
     n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , 
     n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , 
     n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , 
     n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , 
     n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , 
     n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , 
     n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , 
     n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , 
     n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , 
     n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , 
     n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , 
     n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , 
     n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , 
     n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , 
     n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , 
     n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , 
     n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , 
     n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , 
     n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , 
     n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , 
     n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , 
     n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , 
     n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , 
     n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , 
     n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , 
     n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , 
     n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , 
     n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , 
     n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , 
     n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , 
     n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , 
     n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , 
     n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , 
     n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , 
     n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , 
     n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , 
     n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , 
     n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , 
     n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , 
     n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , 
     n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , 
     n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , 
     n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , 
     n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , 
     n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , 
     n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , 
     n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , 
     n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , 
     n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , 
     n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , 
     n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , 
     n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , 
     n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , 
     n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , 
     n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , 
     n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , 
     n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , 
     n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , 
     n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , 
     n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , 
     n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , 
     n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , 
     n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , 
     n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , 
     n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , 
     n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , 
     n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , 
     n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , 
     n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , 
     n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , 
     n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , 
     n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , 
     n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , 
     n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , 
     n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , 
     n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , 
     n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , 
     n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , 
     n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , 
     n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , 
     n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , 
     n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , 
     n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , 
     n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , 
     n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , 
     n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , 
     n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , 
     n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , 
     n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , 
     n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , 
     n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 ;
buf ( n2048 , n12065 );
buf ( n2049 , n12068 );
buf ( n4102 , n1087 );
buf ( n4103 , n1970 );
buf ( n4104 , n1014 );
buf ( n4105 , n484 );
buf ( n4106 , n1812 );
buf ( n4107 , n1992 );
buf ( n4108 , n764 );
buf ( n4109 , n1323 );
buf ( n4110 , n1191 );
buf ( n4111 , n2034 );
buf ( n4112 , n689 );
buf ( n4113 , n365 );
buf ( n4114 , n872 );
buf ( n4115 , n1178 );
buf ( n4116 , n1781 );
buf ( n4117 , n2014 );
buf ( n4118 , n843 );
buf ( n4119 , n1356 );
buf ( n4120 , n1196 );
buf ( n4121 , n339 );
buf ( n4122 , n699 );
buf ( n4123 , n54 );
buf ( n4124 , n958 );
buf ( n4125 , n1227 );
buf ( n4126 , n1525 );
buf ( n4127 , n1317 );
buf ( n4128 , n1389 );
buf ( n4129 , n1821 );
buf ( n4130 , n1845 );
buf ( n4131 , n684 );
buf ( n4132 , n902 );
buf ( n4133 , n975 );
buf ( n4134 , n41 );
buf ( n4135 , n1819 );
buf ( n4136 , n85 );
buf ( n4137 , n1456 );
buf ( n4138 , n768 );
buf ( n4139 , n1823 );
buf ( n4140 , n553 );
buf ( n4141 , n1335 );
buf ( n4142 , n1851 );
buf ( n4143 , n1099 );
buf ( n4144 , n159 );
buf ( n4145 , n1424 );
buf ( n4146 , n74 );
buf ( n4147 , n1991 );
buf ( n4148 , n910 );
buf ( n4149 , n636 );
buf ( n4150 , n720 );
buf ( n4151 , n1116 );
buf ( n4152 , n1990 );
buf ( n4153 , n1865 );
buf ( n4154 , n1403 );
buf ( n4155 , n1627 );
buf ( n4156 , n1901 );
buf ( n4157 , n1442 );
buf ( n4158 , n905 );
buf ( n4159 , n670 );
buf ( n4160 , n1844 );
buf ( n4161 , n1986 );
buf ( n4162 , n473 );
buf ( n4163 , n4 );
buf ( n4164 , n753 );
buf ( n4165 , n37 );
buf ( n4166 , n499 );
buf ( n4167 , n1390 );
buf ( n4168 , n154 );
buf ( n4169 , n774 );
buf ( n4170 , n144 );
buf ( n4171 , n751 );
buf ( n4172 , n1184 );
buf ( n4173 , n1300 );
buf ( n4174 , n348 );
buf ( n4175 , n375 );
buf ( n4176 , n1838 );
buf ( n4177 , n1194 );
buf ( n4178 , n687 );
buf ( n4179 , n743 );
buf ( n4180 , n2002 );
buf ( n4181 , n550 );
buf ( n4182 , n141 );
buf ( n4183 , n721 );
buf ( n4184 , n1949 );
buf ( n4185 , n271 );
buf ( n4186 , n291 );
buf ( n4187 , n58 );
buf ( n4188 , n1615 );
buf ( n4189 , n2019 );
buf ( n4190 , n1164 );
buf ( n4191 , n442 );
buf ( n4192 , n787 );
buf ( n4193 , n1120 );
buf ( n4194 , n1128 );
buf ( n4195 , n609 );
buf ( n4196 , n1364 );
buf ( n4197 , n856 );
buf ( n4198 , n1041 );
buf ( n4199 , n1719 );
buf ( n4200 , n681 );
buf ( n4201 , n1447 );
buf ( n4202 , n1349 );
buf ( n4203 , n1044 );
buf ( n4204 , n915 );
buf ( n4205 , n864 );
buf ( n4206 , n1514 );
buf ( n4207 , n28 );
buf ( n4208 , n1470 );
buf ( n4209 , n458 );
buf ( n4210 , n1828 );
buf ( n4211 , n505 );
buf ( n4212 , n493 );
buf ( n4213 , n1071 );
buf ( n4214 , n673 );
buf ( n4215 , n943 );
buf ( n4216 , n243 );
buf ( n4217 , n111 );
buf ( n4218 , n1051 );
buf ( n4219 , n657 );
buf ( n4220 , n1040 );
buf ( n4221 , n695 );
buf ( n4222 , n2013 );
buf ( n4223 , n371 );
buf ( n4224 , n1354 );
buf ( n4225 , n11 );
buf ( n4226 , n1493 );
buf ( n4227 , n240 );
buf ( n4228 , n1585 );
buf ( n4229 , n1136 );
buf ( n4230 , n302 );
buf ( n4231 , n1151 );
buf ( n4232 , n246 );
buf ( n4233 , n1211 );
buf ( n4234 , n1004 );
buf ( n4235 , n1291 );
buf ( n4236 , n1528 );
buf ( n4237 , n466 );
buf ( n4238 , n709 );
buf ( n4239 , n513 );
buf ( n4240 , n270 );
buf ( n4241 , n1353 );
buf ( n4242 , n1398 );
buf ( n4243 , n44 );
buf ( n4244 , n664 );
buf ( n4245 , n453 );
buf ( n4246 , n735 );
buf ( n4247 , n587 );
buf ( n4248 , n186 );
buf ( n4249 , n1135 );
buf ( n4250 , n1374 );
buf ( n4251 , n117 );
buf ( n4252 , n1422 );
buf ( n4253 , n1249 );
buf ( n4254 , n1799 );
buf ( n4255 , n1843 );
buf ( n4256 , n1898 );
buf ( n4257 , n671 );
buf ( n4258 , n969 );
buf ( n4259 , n1649 );
buf ( n4260 , n1558 );
buf ( n4261 , n1526 );
buf ( n4262 , n248 );
buf ( n4263 , n798 );
buf ( n4264 , n747 );
buf ( n4265 , n221 );
buf ( n4266 , n378 );
buf ( n4267 , n1182 );
buf ( n4268 , n1733 );
buf ( n4269 , n907 );
buf ( n4270 , n998 );
buf ( n4271 , n394 );
buf ( n4272 , n1973 );
buf ( n4273 , n462 );
buf ( n4274 , n1676 );
buf ( n4275 , n1878 );
buf ( n4276 , n794 );
buf ( n4277 , n912 );
buf ( n4278 , n1520 );
buf ( n4279 , n361 );
buf ( n4280 , n59 );
buf ( n4281 , n1953 );
buf ( n4282 , n1365 );
buf ( n4283 , n50 );
buf ( n4284 , n1460 );
buf ( n4285 , n1130 );
buf ( n4286 , n292 );
buf ( n4287 , n479 );
buf ( n4288 , n164 );
buf ( n4289 , n1825 );
buf ( n4290 , n250 );
buf ( n4291 , n767 );
buf ( n4292 , n1137 );
buf ( n4293 , n656 );
buf ( n4294 , n1325 );
buf ( n4295 , n539 );
buf ( n4296 , n1877 );
buf ( n4297 , n802 );
buf ( n4298 , n482 );
buf ( n4299 , n1327 );
buf ( n4300 , n96 );
buf ( n4301 , n771 );
buf ( n4302 , n807 );
buf ( n4303 , n153 );
buf ( n4304 , n1378 );
buf ( n4305 , n160 );
buf ( n4306 , n1033 );
buf ( n4307 , n1553 );
buf ( n4308 , n659 );
buf ( n4309 , n504 );
buf ( n4310 , n858 );
buf ( n4311 , n349 );
buf ( n4312 , n1414 );
buf ( n4313 , n901 );
buf ( n4314 , n1880 );
buf ( n4315 , n836 );
buf ( n4316 , n84 );
buf ( n4317 , n918 );
buf ( n4318 , n742 );
buf ( n4319 , n121 );
buf ( n4320 , n308 );
buf ( n4321 , n252 );
buf ( n4322 , n1421 );
buf ( n4323 , n1654 );
buf ( n4324 , n488 );
buf ( n4325 , n1542 );
buf ( n4326 , n495 );
buf ( n4327 , n1944 );
buf ( n4328 , n1757 );
buf ( n4329 , n238 );
buf ( n4330 , n384 );
buf ( n4331 , n541 );
buf ( n4332 , n210 );
buf ( n4333 , n33 );
buf ( n4334 , n306 );
buf ( n4335 , n459 );
buf ( n4336 , n1190 );
buf ( n4337 , n532 );
buf ( n4338 , n1797 );
buf ( n4339 , n408 );
buf ( n4340 , n1911 );
buf ( n4341 , n1018 );
buf ( n4342 , n108 );
buf ( n4343 , n486 );
buf ( n4344 , n1415 );
buf ( n4345 , n1074 );
buf ( n4346 , n1874 );
buf ( n4347 , n304 );
buf ( n4348 , n1482 );
buf ( n4349 , n318 );
buf ( n4350 , n886 );
buf ( n4351 , n1872 );
buf ( n4352 , n1305 );
buf ( n4353 , n2000 );
buf ( n4354 , n299 );
buf ( n4355 , n1740 );
buf ( n4356 , n307 );
buf ( n4357 , n1189 );
buf ( n4358 , n1622 );
buf ( n4359 , n274 );
buf ( n4360 , n1984 );
buf ( n4361 , n1771 );
buf ( n4362 , n1980 );
buf ( n4363 , n1269 );
buf ( n4364 , n1075 );
buf ( n4365 , n1634 );
buf ( n4366 , n512 );
buf ( n4367 , n1055 );
buf ( n4368 , n322 );
buf ( n4369 , n1009 );
buf ( n4370 , n407 );
buf ( n4371 , n1166 );
buf ( n4372 , n1332 );
buf ( n4373 , n2023 );
buf ( n4374 , n1203 );
buf ( n4375 , n1907 );
buf ( n4376 , n61 );
buf ( n4377 , n580 );
buf ( n4378 , n543 );
buf ( n4379 , n315 );
buf ( n4380 , n295 );
buf ( n4381 , n468 );
buf ( n4382 , n679 );
buf ( n4383 , n558 );
buf ( n4384 , n1271 );
buf ( n4385 , n1850 );
buf ( n4386 , n1406 );
buf ( n4387 , n529 );
buf ( n4388 , n264 );
buf ( n4389 , n545 );
buf ( n4390 , n1232 );
buf ( n4391 , n113 );
buf ( n4392 , n772 );
buf ( n4393 , n1265 );
buf ( n4394 , n518 );
buf ( n4395 , n1100 );
buf ( n4396 , n1814 );
buf ( n4397 , n874 );
buf ( n4398 , n919 );
buf ( n4399 , n1367 );
buf ( n4400 , n1253 );
buf ( n4401 , n1476 );
buf ( n4402 , n1707 );
buf ( n4403 , n913 );
buf ( n4404 , n1085 );
buf ( n4405 , n1724 );
buf ( n4406 , n341 );
buf ( n4407 , n489 );
buf ( n4408 , n1309 );
buf ( n4409 , n1494 );
buf ( n4410 , n1670 );
buf ( n4411 , n1708 );
buf ( n4412 , n1098 );
buf ( n4413 , n968 );
buf ( n4414 , n1048 );
buf ( n4415 , n98 );
buf ( n4416 , n1181 );
buf ( n4417 , n1604 );
buf ( n4418 , n773 );
buf ( n4419 , n1554 );
buf ( n4420 , n1505 );
buf ( n4421 , n1444 );
buf ( n4422 , n999 );
buf ( n4423 , n1225 );
buf ( n4424 , n1696 );
buf ( n4425 , n1152 );
buf ( n4426 , n1363 );
buf ( n4427 , n629 );
buf ( n4428 , n701 );
buf ( n4429 , n1220 );
buf ( n4430 , n1774 );
buf ( n4431 , n1250 );
buf ( n4432 , n10 );
buf ( n4433 , n1715 );
buf ( n4434 , n1320 );
buf ( n4435 , n1432 );
buf ( n4436 , n1139 );
buf ( n4437 , n953 );
buf ( n4438 , n601 );
buf ( n4439 , n200 );
buf ( n4440 , n498 );
buf ( n4441 , n1889 );
buf ( n4442 , n923 );
buf ( n4443 , n632 );
buf ( n4444 , n1789 );
buf ( n4445 , n754 );
buf ( n4446 , n1594 );
buf ( n4447 , n705 );
buf ( n4448 , n319 );
buf ( n4449 , n1875 );
buf ( n4450 , n1321 );
buf ( n4451 , n1223 );
buf ( n4452 , n2018 );
buf ( n4453 , n555 );
buf ( n4454 , n1836 );
buf ( n4455 , n1416 );
buf ( n4456 , n1782 );
buf ( n4457 , n675 );
buf ( n4458 , n961 );
buf ( n4459 , n390 );
buf ( n4460 , n178 );
buf ( n4461 , n1848 );
buf ( n4462 , n1729 );
buf ( n4463 , n211 );
buf ( n4464 , n1854 );
buf ( n4465 , n1668 );
buf ( n4466 , n1868 );
buf ( n4467 , n2 );
buf ( n4468 , n1837 );
buf ( n4469 , n1021 );
buf ( n4470 , n1258 );
buf ( n4471 , n599 );
buf ( n4472 , n1714 );
buf ( n4473 , n1652 );
buf ( n4474 , n1871 );
buf ( n4475 , n748 );
buf ( n4476 , n693 );
buf ( n4477 , n811 );
buf ( n4478 , n1971 );
buf ( n4479 , n1045 );
buf ( n4480 , n623 );
buf ( n4481 , n763 );
buf ( n4482 , n1695 );
buf ( n4483 , n1107 );
buf ( n4484 , n1070 );
buf ( n4485 , n1755 );
buf ( n4486 , n356 );
buf ( n4487 , n978 );
buf ( n4488 , n842 );
buf ( n4489 , n500 );
buf ( n4490 , n1589 );
buf ( n4491 , n133 );
buf ( n4492 , n575 );
buf ( n4493 , n382 );
buf ( n4494 , n337 );
buf ( n4495 , n522 );
buf ( n4496 , n2045 );
buf ( n4497 , n607 );
buf ( n4498 , n678 );
buf ( n4499 , n1308 );
buf ( n4500 , n2003 );
buf ( n4501 , n1013 );
buf ( n4502 , n717 );
buf ( n4503 , n2025 );
buf ( n4504 , n346 );
buf ( n4505 , n228 );
buf ( n4506 , n2030 );
buf ( n4507 , n921 );
buf ( n4508 , n487 );
buf ( n4509 , n651 );
buf ( n4510 , n665 );
buf ( n4511 , n860 );
buf ( n4512 , n1712 );
buf ( n4513 , n426 );
buf ( n4514 , n201 );
buf ( n4515 , n1985 );
buf ( n4516 , n1731 );
buf ( n4517 , n183 );
buf ( n4518 , n1028 );
buf ( n4519 , n866 );
buf ( n4520 , n233 );
buf ( n4521 , n301 );
buf ( n4522 , n281 );
buf ( n4523 , n272 );
buf ( n4524 , n951 );
buf ( n4525 , n142 );
buf ( n4526 , n1104 );
buf ( n4527 , n1728 );
buf ( n4528 , n1902 );
buf ( n4529 , n1785 );
buf ( n4530 , n23 );
buf ( n4531 , n317 );
buf ( n4532 , n1301 );
buf ( n4533 , n1656 );
buf ( n4534 , n1418 );
buf ( n4535 , n1884 );
buf ( n4536 , n1032 );
buf ( n4537 , n621 );
buf ( n4538 , n1611 );
buf ( n4539 , n520 );
buf ( n4540 , n1373 );
buf ( n4541 , n964 );
buf ( n4542 , n132 );
buf ( n4543 , n362 );
buf ( n4544 , n1472 );
buf ( n4545 , n1454 );
buf ( n4546 , n822 );
buf ( n4547 , n286 );
buf ( n4548 , n1133 );
buf ( n4549 , n20 );
buf ( n4550 , n166 );
buf ( n4551 , n1540 );
buf ( n4552 , n1326 );
buf ( n4553 , n654 );
buf ( n4554 , n963 );
buf ( n4555 , n715 );
buf ( n4556 , n1685 );
buf ( n4557 , n818 );
buf ( n4558 , n1701 );
buf ( n4559 , n577 );
buf ( n4560 , n1243 );
buf ( n4561 , n756 );
buf ( n4562 , n2005 );
buf ( n4563 , n437 );
buf ( n4564 , n1257 );
buf ( n4565 , n1951 );
buf ( n4566 , n1697 );
buf ( n4567 , n1228 );
buf ( n4568 , n199 );
buf ( n4569 , n1766 );
buf ( n4570 , n868 );
buf ( n4571 , n399 );
buf ( n4572 , n667 );
buf ( n4573 , n993 );
buf ( n4574 , n1034 );
buf ( n4575 , n120 );
buf ( n4576 , n1934 );
buf ( n4577 , n227 );
buf ( n4578 , n1 );
buf ( n4579 , n7 );
buf ( n4580 , n257 );
buf ( n4581 , n1538 );
buf ( n4582 , n282 );
buf ( n4583 , n1739 );
buf ( n4584 , n1645 );
buf ( n4585 , n1966 );
buf ( n4586 , n853 );
buf ( n4587 , n206 );
buf ( n4588 , n1276 );
buf ( n4589 , n728 );
buf ( n4590 , n1709 );
buf ( n4591 , n691 );
buf ( n4592 , n2033 );
buf ( n4593 , n224 );
buf ( n4594 , n1340 );
buf ( n4595 , n1144 );
buf ( n4596 , n1175 );
buf ( n4597 , n1050 );
buf ( n4598 , n175 );
buf ( n4599 , n1508 );
buf ( n4600 , n1273 );
buf ( n4601 , n704 );
buf ( n4602 , n436 );
buf ( n4603 , n1012 );
buf ( n4604 , n1433 );
buf ( n4605 , n1337 );
buf ( n4606 , n1815 );
buf ( n4607 , n1052 );
buf ( n4608 , n1420 );
buf ( n4609 , n63 );
buf ( n4610 , n1929 );
buf ( n4611 , n2011 );
buf ( n4612 , n1109 );
buf ( n4613 , n109 );
buf ( n4614 , n1921 );
buf ( n4615 , n1895 );
buf ( n4616 , n1219 );
buf ( n4617 , n1576 );
buf ( n4618 , n1173 );
buf ( n4619 , n1684 );
buf ( n4620 , n696 );
buf ( n4621 , n1142 );
buf ( n4622 , n401 );
buf ( n4623 , n994 );
buf ( n4624 , n491 );
buf ( n4625 , n503 );
buf ( n4626 , n1794 );
buf ( n4627 , n1671 );
buf ( n4628 , n589 );
buf ( n4629 , n283 );
buf ( n4630 , n411 );
buf ( n4631 , n597 );
buf ( n4632 , n107 );
buf ( n4633 , n1464 );
buf ( n4634 , n1648 );
buf ( n4635 , n335 );
buf ( n4636 , n1234 );
buf ( n4637 , n841 );
buf ( n4638 , n1593 );
buf ( n4639 , n1503 );
buf ( n4640 , n955 );
buf ( n4641 , n1483 );
buf ( n4642 , n1629 );
buf ( n4643 , n1762 );
buf ( n4644 , n1283 );
buf ( n4645 , n752 );
buf ( n4646 , n1148 );
buf ( n4647 , n494 );
buf ( n4648 , n628 );
buf ( n4649 , n1093 );
buf ( n4650 , n99 );
buf ( n4651 , n1820 );
buf ( n4652 , n1431 );
buf ( n4653 , n455 );
buf ( n4654 , n1333 );
buf ( n4655 , n1847 );
buf ( n4656 , n276 );
buf ( n4657 , n25 );
buf ( n4658 , n1726 );
buf ( n4659 , n27 );
buf ( n4660 , n95 );
buf ( n4661 , n176 );
buf ( n4662 , n1858 );
buf ( n4663 , n602 );
buf ( n4664 , n1002 );
buf ( n4665 , n1926 );
buf ( n4666 , n1060 );
buf ( n4667 , n1817 );
buf ( n4668 , n1519 );
buf ( n4669 , n548 );
buf ( n4670 , n987 );
buf ( n4671 , n1072 );
buf ( n4672 , n2028 );
buf ( n4673 , n406 );
buf ( n4674 , n93 );
buf ( n4675 , n846 );
buf ( n4676 , n852 );
buf ( n4677 , n1555 );
buf ( n4678 , n1818 );
buf ( n4679 , n1600 );
buf ( n4680 , n1123 );
buf ( n4681 , n1610 );
buf ( n4682 , n899 );
buf ( n4683 , n538 );
buf ( n4684 , n829 );
buf ( n4685 , n1924 );
buf ( n4686 , n1653 );
buf ( n4687 , n372 );
buf ( n4688 , n1206 );
buf ( n4689 , n1029 );
buf ( n4690 , n1678 );
buf ( n4691 , n959 );
buf ( n4692 , n1094 );
buf ( n4693 , n834 );
buf ( n4694 , n260 );
buf ( n4695 , n1480 );
buf ( n4696 , n104 );
buf ( n4697 , n820 );
buf ( n4698 , n576 );
buf ( n4699 , n592 );
buf ( n4700 , n103 );
buf ( n4701 , n396 );
buf ( n4702 , n388 );
buf ( n4703 , n1246 );
buf ( n4704 , n2029 );
buf ( n4705 , n582 );
buf ( n4706 , n1037 );
buf ( n4707 , n509 );
buf ( n4708 , n13 );
buf ( n4709 , n168 );
buf ( n4710 , n1428 );
buf ( n4711 , n22 );
buf ( n4712 , n1570 );
buf ( n4713 , n1743 );
buf ( n4714 , n1643 );
buf ( n4715 , n1853 );
buf ( n4716 , n757 );
buf ( n4717 , n1955 );
buf ( n4718 , n981 );
buf ( n4719 , n941 );
buf ( n4720 , n561 );
buf ( n4721 , n1964 );
buf ( n4722 , n564 );
buf ( n4723 , n979 );
buf ( n4724 , n563 );
buf ( n4725 , n719 );
buf ( n4726 , n1609 );
buf ( n4727 , n106 );
buf ( n4728 , n32 );
buf ( n4729 , n62 );
buf ( n4730 , n1746 );
buf ( n4731 , n42 );
buf ( n4732 , n514 );
buf ( n4733 , n21 );
buf ( n4734 , n583 );
buf ( n4735 , n1459 );
buf ( n4736 , n1376 );
buf ( n4737 , n1703 );
buf ( n4738 , n929 );
buf ( n4739 , n631 );
buf ( n4740 , n1019 );
buf ( n4741 , n1391 );
buf ( n4742 , n793 );
buf ( n4743 , n1958 );
buf ( n4744 , n151 );
buf ( n4745 , n1198 );
buf ( n4746 , n1150 );
buf ( n4747 , n380 );
buf ( n4748 , n497 );
buf ( n4749 , n1122 );
buf ( n4750 , n1727 );
buf ( n4751 , n634 );
buf ( n4752 , n660 );
buf ( n4753 , n88 );
buf ( n4754 , n1068 );
buf ( n4755 , n507 );
buf ( n4756 , n983 );
buf ( n4757 , n1942 );
buf ( n4758 , n1550 );
buf ( n4759 , n1575 );
buf ( n4760 , n1950 );
buf ( n4761 , n926 );
buf ( n4762 , n700 );
buf ( n4763 , n415 );
buf ( n4764 , n1097 );
buf ( n4765 , n851 );
buf ( n4766 , n2040 );
buf ( n4767 , n418 );
buf ( n4768 , n1690 );
buf ( n4769 , n930 );
buf ( n4770 , n305 );
buf ( n4771 , n1336 );
buf ( n4772 , n616 );
buf ( n4773 , n1434 );
buf ( n4774 , n31 );
buf ( n4775 , n460 );
buf ( n4776 , n1530 );
buf ( n4777 , n796 );
buf ( n4778 , n197 );
buf ( n4779 , n1382 );
buf ( n4780 , n1084 );
buf ( n4781 , n1761 );
buf ( n4782 , n803 );
buf ( n4783 , n1972 );
buf ( n4784 , n17 );
buf ( n4785 , n765 );
buf ( n4786 , n136 );
buf ( n4787 , n1487 );
buf ( n4788 , n26 );
buf ( n4789 , n1026 );
buf ( n4790 , n1461 );
buf ( n4791 , n1229 );
buf ( n4792 , n1736 );
buf ( n4793 , n683 );
buf ( n4794 , n540 );
buf ( n4795 , n1486 );
buf ( n4796 , n862 );
buf ( n4797 , n1778 );
buf ( n4798 , n1607 );
buf ( n4799 , n703 );
buf ( n4800 , n888 );
buf ( n4801 , n1800 );
buf ( n4802 , n1010 );
buf ( n4803 , n966 );
buf ( n4804 , n1210 );
buf ( n4805 , n1711 );
buf ( n4806 , n729 );
buf ( n4807 , n674 );
buf ( n4808 , n69 );
buf ( n4809 , n1891 );
buf ( n4810 , n76 );
buf ( n4811 , n658 );
buf ( n4812 , n1568 );
buf ( n4813 , n1202 );
buf ( n4814 , n1205 );
buf ( n4815 , n311 );
buf ( n4816 , n284 );
buf ( n4817 , n896 );
buf ( n4818 , n448 );
buf ( n4819 , n1822 );
buf ( n4820 , n1215 );
buf ( n4821 , n82 );
buf ( n4822 , n1038 );
buf ( n4823 , n1282 );
buf ( n4824 , n1485 );
buf ( n4825 , n1020 );
buf ( n4826 , n1466 );
buf ( n4827 , n1260 );
buf ( n4828 , n770 );
buf ( n4829 , n105 );
buf ( n4830 , n1939 );
buf ( n4831 , n1601 );
buf ( n4832 , n710 );
buf ( n4833 , n1764 );
buf ( n4834 , n1932 );
buf ( n4835 , n1125 );
buf ( n4836 , n472 );
buf ( n4837 , n52 );
buf ( n4838 , n112 );
buf ( n4839 , n179 );
buf ( n4840 , n1439 );
buf ( n4841 , n1295 );
buf ( n4842 , n43 );
buf ( n4843 , n1718 );
buf ( n4844 , n1298 );
buf ( n4845 , n973 );
buf ( n4846 , n156 );
buf ( n4847 , n65 );
buf ( n4848 , n739 );
buf ( n4849 , n1890 );
buf ( n4850 , n413 );
buf ( n4851 , n1752 );
buf ( n4852 , n551 );
buf ( n4853 , n1941 );
buf ( n4854 , n1830 );
buf ( n4855 , n1056 );
buf ( n4856 , n1169 );
buf ( n4857 , n1413 );
buf ( n4858 , n1968 );
buf ( n4859 , n417 );
buf ( n4860 , n452 );
buf ( n4861 , n680 );
buf ( n4862 , n934 );
buf ( n4863 , n219 );
buf ( n4864 , n2016 );
buf ( n4865 , n1446 );
buf ( n4866 , n6 );
buf ( n4867 , n1174 );
buf ( n4868 , n931 );
buf ( n4869 , n1999 );
buf ( n4870 , n731 );
buf ( n4871 , n556 );
buf ( n4872 , n1905 );
buf ( n4873 , n1769 );
buf ( n4874 , n1277 );
buf ( n4875 , n1088 );
buf ( n4876 , n1448 );
buf ( n4877 , n1974 );
buf ( n4878 , n414 );
buf ( n4879 , n1281 );
buf ( n4880 , n1165 );
buf ( n4881 , n158 );
buf ( n4882 , n1686 );
buf ( n4883 , n1650 );
buf ( n4884 , n204 );
buf ( n4885 , n1552 );
buf ( n4886 , n1887 );
buf ( n4887 , n1304 );
buf ( n4888 , n1209 );
buf ( n4889 , n1348 );
buf ( n4890 , n1946 );
buf ( n4891 , n554 );
buf ( n4892 , n944 );
buf ( n4893 , n1183 );
buf ( n4894 , n1179 );
buf ( n4895 , n278 );
buf ( n4896 , n789 );
buf ( n4897 , n1744 );
buf ( n4898 , n1914 );
buf ( n4899 , n936 );
buf ( n4900 , n1680 );
buf ( n4901 , n932 );
buf ( n4902 , n761 );
buf ( n4903 , n1319 );
buf ( n4904 , n230 );
buf ( n4905 , n892 );
buf ( n4906 , n620 );
buf ( n4907 , n245 );
buf ( n4908 , n110 );
buf ( n4909 , n783 );
buf ( n4910 , n1831 );
buf ( n4911 , n1560 );
buf ( n4912 , n702 );
buf ( n4913 , n135 );
buf ( n4914 , n269 );
buf ( n4915 , n323 );
buf ( n4916 , n1780 );
buf ( n4917 , n805 );
buf ( n4918 , n711 );
buf ( n4919 , n1866 );
buf ( n4920 , n1532 );
buf ( n4921 , n1621 );
buf ( n4922 , n1000 );
buf ( n4923 , n1252 );
buf ( n4924 , n644 );
buf ( n4925 , n1141 );
buf ( n4926 , n835 );
buf ( n4927 , n1919 );
buf ( n4928 , n212 );
buf ( n4929 , n1734 );
buf ( n4930 , n769 );
buf ( n4931 , n1763 );
buf ( n4932 , n123 );
buf ( n4933 , n444 );
buf ( n4934 , n78 );
buf ( n4935 , n287 );
buf ( n4936 , n430 );
buf ( n4937 , n2032 );
buf ( n4938 , n454 );
buf ( n4939 , n1917 );
buf ( n4940 , n440 );
buf ( n4941 , n358 );
buf ( n4942 , n1379 );
buf ( n4943 , n1278 );
buf ( n4944 , n1313 );
buf ( n4945 , n714 );
buf ( n4946 , n828 );
buf ( n4947 , n277 );
buf ( n4948 , n1126 );
buf ( n4949 , n690 );
buf ( n4950 , n546 );
buf ( n4951 , n1140 );
buf ( n4952 , n392 );
buf ( n4953 , n855 );
buf ( n4954 , n1846 );
buf ( n4955 , n1943 );
buf ( n4956 , n1360 );
buf ( n4957 , n155 );
buf ( n4958 , n359 );
buf ( n4959 , n1691 );
buf ( n4960 , n1092 );
buf ( n4961 , n226 );
buf ( n4962 , n2001 );
buf ( n4963 , n445 );
buf ( n4964 , n1386 );
buf ( n4965 , n1938 );
buf ( n4966 , n1900 );
buf ( n4967 , n1147 );
buf ( n4968 , n1279 );
buf ( n4969 , n1543 );
buf ( n4970 , n647 );
buf ( n4971 , n1153 );
buf ( n4972 , n333 );
buf ( n4973 , n310 );
buf ( n4974 , n639 );
buf ( n4975 , n971 );
buf ( n4976 , n1510 );
buf ( n4977 , n1748 );
buf ( n4978 , n1419 );
buf ( n4979 , n937 );
buf ( n4980 , n1081 );
buf ( n4981 , n1810 );
buf ( n4982 , n1637 );
buf ( n4983 , n935 );
buf ( n4984 , n1860 );
buf ( n4985 , n662 );
buf ( n4986 , n900 );
buf ( n4987 , n1384 );
buf ( n4988 , n126 );
buf ( n4989 , n235 );
buf ( n4990 , n1145 );
buf ( n4991 , n573 );
buf ( n4992 , n1162 );
buf ( n4993 , n724 );
buf ( n4994 , n1867 );
buf ( n4995 , n1082 );
buf ( n4996 , n697 );
buf ( n4997 , n1963 );
buf ( n4998 , n191 );
buf ( n4999 , n1438 );
buf ( n5000 , n1358 );
buf ( n5001 , n1467 );
buf ( n5002 , n1784 );
buf ( n5003 , n496 );
buf ( n5004 , n2027 );
buf ( n5005 , n140 );
buf ( n5006 , n1638 );
buf ( n5007 , n861 );
buf ( n5008 , n942 );
buf ( n5009 , n1534 );
buf ( n5010 , n649 );
buf ( n5011 , n1710 );
buf ( n5012 , n1616 );
buf ( n5013 , n766 );
buf ( n5014 , n909 );
buf ( n5015 , n1046 );
buf ( n5016 , n363 );
buf ( n5017 , n619 );
buf ( n5018 , n1591 );
buf ( n5019 , n1411 );
buf ( n5020 , n1569 );
buf ( n5021 , n1338 );
buf ( n5022 , n925 );
buf ( n5023 , n1108 );
buf ( n5024 , n1161 );
buf ( n5025 , n1387 );
buf ( n5026 , n1381 );
buf ( n5027 , n637 );
buf ( n5028 , n1346 );
buf ( n5029 , n429 );
buf ( n5030 , n605 );
buf ( n5031 , n1222 );
buf ( n5032 , n1952 );
buf ( n5033 , n1073 );
buf ( n5034 , n741 );
buf ( n5035 , n736 );
buf ( n5036 , n184 );
buf ( n5037 , n830 );
buf ( n5038 , n1400 );
buf ( n5039 , n1635 );
buf ( n5040 , n1978 );
buf ( n5041 , n73 );
buf ( n5042 , n1549 );
buf ( n5043 , n1588 );
buf ( n5044 , n379 );
buf ( n5045 , n1006 );
buf ( n5046 , n1647 );
buf ( n5047 , n410 );
buf ( n5048 , n476 );
buf ( n5049 , n1172 );
buf ( n5050 , n1993 );
buf ( n5051 , n222 );
buf ( n5052 , n606 );
buf ( n5053 , n1256 );
buf ( n5054 , n1267 );
buf ( n5055 , n579 );
buf ( n5056 , n531 );
buf ( n5057 , n1347 );
buf ( n5058 , n878 );
buf ( n5059 , n1054 );
buf ( n5060 , n1912 );
buf ( n5061 , n1016 );
buf ( n5062 , n14 );
buf ( n5063 , n1582 );
buf ( n5064 , n1156 );
buf ( n5065 , n1674 );
buf ( n5066 , n457 );
buf ( n5067 , n526 );
buf ( n5068 , n775 );
buf ( n5069 , n1523 );
buf ( n5070 , n2037 );
buf ( n5071 , n517 );
buf ( n5072 , n1790 );
buf ( n5073 , n1357 );
buf ( n5074 , n1931 );
buf ( n5075 , n880 );
buf ( n5076 , n972 );
buf ( n5077 , n1535 );
buf ( n5078 , n35 );
buf ( n5079 , n97 );
buf ( n5080 , n1940 );
buf ( n5081 , n837 );
buf ( n5082 , n485 );
buf ( n5083 , n321 );
buf ( n5084 , n1630 );
buf ( n5085 , n799 );
buf ( n5086 , n1813 );
buf ( n5087 , n1001 );
buf ( n5088 , n1079 );
buf ( n5089 , n813 );
buf ( n5090 , n1673 );
buf ( n5091 , n648 );
buf ( n5092 , n122 );
buf ( n5093 , n1773 );
buf ( n5094 , n279 );
buf ( n5095 , n1160 );
buf ( n5096 , n1641 );
buf ( n5097 , n642 );
buf ( n5098 , n2004 );
buf ( n5099 , n334 );
buf ( n5100 , n1511 );
buf ( n5101 , n1385 );
buf ( n5102 , n1965 );
buf ( n5103 , n231 );
buf ( n5104 , n446 );
buf ( n5105 , n1592 );
buf ( n5106 , n1956 );
buf ( n5107 , n949 );
buf ( n5108 , n947 );
buf ( n5109 , n330 );
buf ( n5110 , n139 );
buf ( n5111 , n119 );
buf ( n5112 , n60 );
buf ( n5113 , n1443 );
buf ( n5114 , n1584 );
buf ( n5115 , n351 );
buf ( n5116 , n1863 );
buf ( n5117 , n1248 );
buf ( n5118 , n984 );
buf ( n5119 , n1612 );
buf ( n5120 , n225 );
buf ( n5121 , n1617 );
buf ( n5122 , n370 );
buf ( n5123 , n463 );
buf ( n5124 , n147 );
buf ( n5125 , n604 );
buf ( n5126 , n1529 );
buf ( n5127 , n1826 );
buf ( n5128 , n1613 );
buf ( n5129 , n1185 );
buf ( n5130 , n1791 );
buf ( n5131 , n624 );
buf ( n5132 , n977 );
buf ( n5133 , n1168 );
buf ( n5134 , n524 );
buf ( n5135 , n1987 );
buf ( n5136 , n1188 );
buf ( n5137 , n1566 );
buf ( n5138 , n1722 );
buf ( n5139 , n24 );
buf ( n5140 , n521 );
buf ( n5141 , n1015 );
buf ( n5142 , n706 );
buf ( n5143 , n1027 );
buf ( n5144 , n885 );
buf ( n5145 , n1977 );
buf ( n5146 , n1361 );
buf ( n5147 , n1275 );
buf ( n5148 , n733 );
buf ( n5149 , n970 );
buf ( n5150 , n530 );
buf ( n5151 , n962 );
buf ( n5152 , n633 );
buf ( n5153 , n1264 );
buf ( n5154 , n409 );
buf ( n5155 , n1435 );
buf ( n5156 , n1565 );
buf ( n5157 , n1005 );
buf ( n5158 , n1064 );
buf ( n5159 , n1672 );
buf ( n5160 , n297 );
buf ( n5161 , n1692 );
buf ( n5162 , n433 );
buf ( n5163 , n46 );
buf ( n5164 , n461 );
buf ( n5165 , n613 );
buf ( n5166 , n884 );
buf ( n5167 , n911 );
buf ( n5168 , n3 );
buf ( n5169 , n1240 );
buf ( n5170 , n1192 );
buf ( n5171 , n1661 );
buf ( n5172 , n1475 );
buf ( n5173 , n786 );
buf ( n5174 , n572 );
buf ( n5175 , n1341 );
buf ( n5176 , n181 );
buf ( n5177 , n1134 );
buf ( n5178 , n1628 );
buf ( n5179 , n1839 );
buf ( n5180 , n650 );
buf ( n5181 , n873 );
buf ( n5182 , n1788 );
buf ( n5183 , n1735 );
buf ( n5184 , n1557 );
buf ( n5185 , n173 );
buf ( n5186 , n991 );
buf ( n5187 , n1217 );
buf ( n5188 , n332 );
buf ( n5189 , n328 );
buf ( n5190 , n1401 );
buf ( n5191 , n1423 );
buf ( n5192 , n1124 );
buf ( n5193 , n1700 );
buf ( n5194 , n614 );
buf ( n5195 , n760 );
buf ( n5196 , n1042 );
buf ( n5197 , n383 );
buf ( n5198 , n1266 );
buf ( n5199 , n920 );
buf ( n5200 , n825 );
buf ( n5201 , n1103 );
buf ( n5202 , n265 );
buf ( n5203 , n1372 );
buf ( n5204 , n938 );
buf ( n5205 , n234 );
buf ( n5206 , n1577 );
buf ( n5207 , n1078 );
buf ( n5208 , n169 );
buf ( n5209 , n474 );
buf ( n5210 , n1329 );
buf ( n5211 , n266 );
buf ( n5212 , n557 );
buf ( n5213 , n1767 );
buf ( n5214 , n1669 );
buf ( n5215 , n1177 );
buf ( n5216 , n1368 );
buf ( n5217 , n1515 );
buf ( n5218 , n343 );
buf ( n5219 , n1207 );
buf ( n5220 , n1808 );
buf ( n5221 , n1783 );
buf ( n5222 , n134 );
buf ( n5223 , n814 );
buf ( n5224 , n5 );
buf ( n5225 , n627 );
buf ( n5226 , n1948 );
buf ( n5227 , n1869 );
buf ( n5228 , n1720 );
buf ( n5229 , n145 );
buf ( n5230 , n1352 );
buf ( n5231 , n738 );
buf ( n5232 , n1286 );
buf ( n5233 , n172 );
buf ( n5234 , n1396 );
buf ( n5235 , n867 );
buf ( n5236 , n995 );
buf ( n5237 , n1402 );
buf ( n5238 , n1682 );
buf ( n5239 , n996 );
buf ( n5240 , n125 );
buf ( n5241 , n38 );
buf ( n5242 , n432 );
buf ( n5243 , n570 );
buf ( n5244 , n598 );
buf ( n5245 , n1187 );
buf ( n5246 , n1312 );
buf ( n5247 , n584 );
buf ( n5248 , n40 );
buf ( n5249 , n585 );
buf ( n5250 , n1539 );
buf ( n5251 , n256 );
buf ( n5252 , n922 );
buf ( n5253 , n102 );
buf ( n5254 , n847 );
buf ( n5255 , n1732 );
buf ( n5256 , n75 );
buf ( n5257 , n2010 );
buf ( n5258 , n324 );
buf ( n5259 , n779 );
buf ( n5260 , n1294 );
buf ( n5261 , n1614 );
buf ( n5262 , n1377 );
buf ( n5263 , n1201 );
buf ( n5264 , n1631 );
buf ( n5265 , n694 );
buf ( n5266 , n1412 );
buf ( n5267 , n1573 );
buf ( n5268 , n100 );
buf ( n5269 , n1025 );
buf ( n5270 , n1285 );
buf ( n5271 , n1981 );
buf ( n5272 , n1105 );
buf ( n5273 , n1500 );
buf ( n5274 , n1681 );
buf ( n5275 , n2036 );
buf ( n5276 , n1798 );
buf ( n5277 , n1666 );
buf ( n5278 , n1910 );
buf ( n5279 , n2041 );
buf ( n5280 , n1859 );
buf ( n5281 , n713 );
buf ( n5282 , n1303 );
buf ( n5283 , n1501 );
buf ( n5284 , n1302 );
buf ( n5285 , n1399 );
buf ( n5286 , n1053 );
buf ( n5287 , n745 );
buf ( n5288 , n1504 );
buf ( n5289 , n171 );
buf ( n5290 , n622 );
buf ( n5291 , n894 );
buf ( n5292 , n47 );
buf ( n5293 , n1531 );
buf ( n5294 , n1114 );
buf ( n5295 , n115 );
buf ( n5296 , n1102 );
buf ( n5297 , n933 );
buf ( n5298 , n1989 );
buf ( n5299 , n387 );
buf ( n5300 , n832 );
buf ( n5301 , n268 );
buf ( n5302 , n1765 );
buf ( n5303 , n1003 );
buf ( n5304 , n1598 );
buf ( n5305 , n954 );
buf ( n5306 , n1959 );
buf ( n5307 , n1675 );
buf ( n5308 , n508 );
buf ( n5309 , n1430 );
buf ( n5310 , n67 );
buf ( n5311 , n1429 );
buf ( n5312 , n131 );
buf ( n5313 , n56 );
buf ( n5314 , n612 );
buf ( n5315 , n247 );
buf ( n5316 , n1835 );
buf ( n5317 , n1067 );
buf ( n5318 , n1129 );
buf ( n5319 , n1270 );
buf ( n5320 , n1693 );
buf ( n5321 , n354 );
buf ( n5322 , n1506 );
buf ( n5323 , n1199 );
buf ( n5324 , n1197 );
buf ( n5325 , n190 );
buf ( n5326 , n1745 );
buf ( n5327 , n1587 );
buf ( n5328 , n1827 );
buf ( n5329 , n782 );
buf ( n5330 , n1477 );
buf ( n5331 , n138 );
buf ( n5332 , n1235 );
buf ( n5333 , n1545 );
buf ( n5334 , n1662 );
buf ( n5335 , n1975 );
buf ( n5336 , n1138 );
buf ( n5337 , n331 );
buf ( n5338 , n810 );
buf ( n5339 , n844 );
buf ( n5340 , n209 );
buf ( n5341 , n55 );
buf ( n5342 , n1117 );
buf ( n5343 , n1288 );
buf ( n5344 , n1086 );
buf ( n5345 , n965 );
buf ( n5346 , n916 );
buf ( n5347 , n220 );
buf ( n5348 , n86 );
buf ( n5349 , n1426 );
buf ( n5350 , n288 );
buf ( n5351 , n1284 );
buf ( n5352 , n727 );
buf ( n5353 , n2020 );
buf ( n5354 , n1925 );
buf ( n5355 , n1478 );
buf ( n5356 , n1876 );
buf ( n5357 , n1463 );
buf ( n5358 , n1742 );
buf ( n5359 , n870 );
buf ( n5360 , n165 );
buf ( n5361 , n788 );
buf ( n5362 , n1343 );
buf ( n5363 , n1954 );
buf ( n5364 , n1920 );
buf ( n5365 , n1238 );
buf ( n5366 , n16 );
buf ( n5367 , n549 );
buf ( n5368 , n1772 );
buf ( n5369 , n1706 );
buf ( n5370 , n1121 );
buf ( n5371 , n471 );
buf ( n5372 , n2044 );
buf ( n5373 , n1608 );
buf ( n5374 , n1721 );
buf ( n5375 , n750 );
buf ( n5376 , n1289 );
buf ( n5377 , n1299 );
buf ( n5378 , n1596 );
buf ( n5379 , n1119 );
buf ( n5380 , n483 );
buf ( n5381 , n1111 );
buf ( n5382 , n1747 );
buf ( n5383 , n2047 );
buf ( n5384 , n1410 );
buf ( n5385 , n1417 );
buf ( n5386 , n1131 );
buf ( n5387 , n1328 );
buf ( n5388 , n1473 );
buf ( n5389 , n781 );
buf ( n5390 , n1049 );
buf ( n5391 , n824 );
buf ( n5392 , n403 );
buf ( n5393 , n2022 );
buf ( n5394 , n646 );
buf ( n5395 , n1908 );
buf ( n5396 , n603 );
buf ( n5397 , n68 );
buf ( n5398 , n1787 );
buf ( n5399 , n215 );
buf ( n5400 , n1663 );
buf ( n5401 , n980 );
buf ( n5402 , n1713 );
buf ( n5403 , n523 );
buf ( n5404 , n1095 );
buf ( n5405 , n800 );
buf ( n5406 , n1563 );
buf ( n5407 , n1106 );
buf ( n5408 , n708 );
buf ( n5409 , n875 );
buf ( n5410 , n12 );
buf ( n5411 , n39 );
buf ( n5412 , n707 );
buf ( n5413 , n1268 );
buf ( n5414 , n1345 );
buf ( n5415 , n1832 );
buf ( n5416 , n641 );
buf ( n5417 , n1306 );
buf ( n5418 , n1311 );
buf ( n5419 , n369 );
buf ( n5420 , n778 );
buf ( n5421 , n982 );
buf ( n5422 , n1171 );
buf ( n5423 , n1779 );
buf ( n5424 , n1751 );
buf ( n5425 , n1132 );
buf ( n5426 , n595 );
buf ( n5427 , n1375 );
buf ( n5428 , n1567 );
buf ( n5429 , n1509 );
buf ( n5430 , n1659 );
buf ( n5431 , n1262 );
buf ( n5432 , n298 );
buf ( n5433 , n1492 );
buf ( n5434 , n192 );
buf ( n5435 , n1259 );
buf ( n5436 , n1170 );
buf ( n5437 , n188 );
buf ( n5438 , n1502 );
buf ( n5439 , n730 );
buf ( n5440 , n1982 );
buf ( n5441 , n1768 );
buf ( n5442 , n1888 );
buf ( n5443 , n986 );
buf ( n5444 , n127 );
buf ( n5445 , n1922 );
buf ( n5446 , n590 );
buf ( n5447 , n515 );
buf ( n5448 , n1517 );
buf ( n5449 , n1469 );
buf ( n5450 , n313 );
buf ( n5451 , n116 );
buf ( n5452 , n1918 );
buf ( n5453 , n150 );
buf ( n5454 , n1792 );
buf ( n5455 , n1091 );
buf ( n5456 , n1307 );
buf ( n5457 , n869 );
buf ( n5458 , n535 );
buf ( n5459 , n1829 );
buf ( n5460 , n280 );
buf ( n5461 , n422 );
buf ( n5462 , n490 );
buf ( n5463 , n777 );
buf ( n5464 , n1069 );
buf ( n5465 , n1886 );
buf ( n5466 , n216 );
buf ( n5467 , n2043 );
buf ( n5468 , n1436 );
buf ( n5469 , n967 );
buf ( n5470 , n808 );
buf ( n5471 , n990 );
buf ( n5472 , n1449 );
buf ( n5473 , n904 );
buf ( n5474 , n1405 );
buf ( n5475 , n391 );
buf ( n5476 , n434 );
buf ( n5477 , n1625 );
buf ( n5478 , n1497 );
buf ( n5479 , n574 );
buf ( n5480 , n1870 );
buf ( n5481 , n865 );
buf ( n5482 , n381 );
buf ( n5483 , n876 );
buf ( n5484 , n685 );
buf ( n5485 , n565 );
buf ( n5486 , n467 );
buf ( n5487 , n1897 );
buf ( n5488 , n101 );
buf ( n5489 , n1058 );
buf ( n5490 , n625 );
buf ( n5491 , n36 );
buf ( n5492 , n49 );
buf ( n5493 , n1857 );
buf ( n5494 , n945 );
buf ( n5495 , n1274 );
buf ( n5496 , n882 );
buf ( n5497 , n229 );
buf ( n5498 , n1683 );
buf ( n5499 , n533 );
buf ( n5500 , n1513 );
buf ( n5501 , n327 );
buf ( n5502 , n1660 );
buf ( n5503 , n237 );
buf ( n5504 , n1705 );
buf ( n5505 , n478 );
buf ( n5506 , n1796 );
buf ( n5507 , n780 );
buf ( n5508 , n129 );
buf ( n5509 , n1688 );
buf ( n5510 , n1590 );
buf ( n5511 , n1244 );
buf ( n5512 , n626 );
buf ( n5513 , n1620 );
buf ( n5514 , n423 );
buf ( n5515 , n1842 );
buf ( n5516 , n661 );
buf ( n5517 , n797 );
buf ( n5518 , n1110 );
buf ( n5519 , n249 );
buf ( n5520 , n94 );
buf ( n5521 , n755 );
buf ( n5522 , n1885 );
buf ( n5523 , n1224 );
buf ( n5524 , n501 );
buf ( n5525 , n666 );
buf ( n5526 , n1490 );
buf ( n5527 , n91 );
buf ( n5528 , n898 );
buf ( n5529 , n903 );
buf ( n5530 , n336 );
buf ( n5531 , n946 );
buf ( n5532 , n326 );
buf ( n5533 , n817 );
buf ( n5534 , n2024 );
buf ( n5535 , n823 );
buf ( n5536 , n1516 );
buf ( n5537 , n1961 );
buf ( n5538 , n1579 );
buf ( n5539 , n1527 );
buf ( n5540 , n924 );
buf ( n5541 , n87 );
buf ( n5542 , n889 );
buf ( n5543 , n242 );
buf ( n5544 , n1619 );
buf ( n5545 , n1581 );
buf ( n5546 , n863 );
buf ( n5547 , n1393 );
buf ( n5548 , n1218 );
buf ( n5549 , n1664 );
buf ( n5550 , n393 );
buf ( n5551 , n263 );
buf ( n5552 , n1759 );
buf ( n5553 , n143 );
buf ( n5554 , n1899 );
buf ( n5555 , n1957 );
buf ( n5556 , n1180 );
buf ( n5557 , n1380 );
buf ( n5558 , n450 );
buf ( n5559 , n1394 );
buf ( n5560 , n443 );
buf ( n5561 , n1541 );
buf ( n5562 , n1292 );
buf ( n5563 , n163 );
buf ( n5564 , n189 );
buf ( n5565 , n1988 );
buf ( n5566 , n424 );
buf ( n5567 , n1024 );
buf ( n5568 , n350 );
buf ( n5569 , n1626 );
buf ( n5570 , n1061 );
buf ( n5571 , n402 );
buf ( n5572 , n239 );
buf ( n5573 , n80 );
buf ( n5574 , n1564 );
buf ( n5575 , n1521 );
buf ( n5576 , n2007 );
buf ( n5577 , n1795 );
buf ( n5578 , n352 );
buf ( n5579 , n149 );
buf ( n5580 , n806 );
buf ( n5581 , n130 );
buf ( n5582 , n1802 );
buf ( n5583 , n1484 );
buf ( n5584 , n1314 );
buf ( n5585 , n71 );
buf ( n5586 , n477 );
buf ( n5587 , n1090 );
buf ( n5588 , n1066 );
buf ( n5589 , n289 );
buf ( n5590 , n718 );
buf ( n5591 , n1369 );
buf ( n5592 , n1556 );
buf ( n5593 , n1602 );
buf ( n5594 , n1080 );
buf ( n5595 , n1351 );
buf ( n5596 , n871 );
buf ( n5597 , n1651 );
buf ( n5598 , n516 );
buf ( n5599 , n1548 );
buf ( n5600 , n833 );
buf ( n5601 , n676 );
buf ( n5602 , n464 );
buf ( n5603 , n1427 );
buf ( n5604 , n1639 );
buf ( n5605 , n1409 );
buf ( n5606 , n569 );
buf ( n5607 , n725 );
buf ( n5608 , n425 );
buf ( n5609 , n1896 );
buf ( n5610 , n1221 );
buf ( n5611 , n1008 );
buf ( n5612 , n1623 );
buf ( n5613 , n859 );
buf ( n5614 , n376 );
buf ( n5615 , n722 );
buf ( n5616 , n2039 );
buf ( n5617 , n534 );
buf ( n5618 , n1297 );
buf ( n5619 , n421 );
buf ( n5620 , n428 );
buf ( n5621 , n427 );
buf ( n5622 , n527 );
buf ( n5623 , n1247 );
buf ( n5624 , n939 );
buf ( n5625 , n79 );
buf ( n5626 , n682 );
buf ( n5627 , n66 );
buf ( n5628 , n740 );
buf ( n5629 , n2006 );
buf ( n5630 , n267 );
buf ( n5631 , n1272 );
buf ( n5632 , n1873 );
buf ( n5633 , n1770 );
buf ( n5634 , n758 );
buf ( n5635 , n1879 );
buf ( n5636 , n956 );
buf ( n5637 , n1362 );
buf ( n5638 , n1065 );
buf ( n5639 , n525 );
buf ( n5640 , n1583 );
buf ( n5641 , n1862 );
buf ( n5642 , n1642 );
buf ( n5643 , n1906 );
buf ( n5644 , n456 );
buf ( n5645 , n398 );
buf ( n5646 , n81 );
buf ( n5647 , n668 );
buf ( n5648 , n831 );
buf ( n5649 , n72 );
buf ( n5650 , n1524 );
buf ( n5651 , n839 );
buf ( n5652 , n511 );
buf ( n5653 , n838 );
buf ( n5654 , n1574 );
buf ( n5655 , n92 );
buf ( n5656 , n1355 );
buf ( n5657 , n217 );
buf ( n5658 , n1687 );
buf ( n5659 , n784 );
buf ( n5660 , n1840 );
buf ( n5661 , n1457 );
buf ( n5662 , n906 );
buf ( n5663 , n1913 );
buf ( n5664 , n1230 );
buf ( n5665 , n1881 );
buf ( n5666 , n566 );
buf ( n5667 , n1499 );
buf ( n5668 , n451 );
buf ( n5669 , n1462 );
buf ( n5670 , n536 );
buf ( n5671 , n1915 );
buf ( n5672 , n1893 );
buf ( n5673 , n157 );
buf ( n5674 , n1293 );
buf ( n5675 , n357 );
buf ( n5676 , n1440 );
buf ( n5677 , n1233 );
buf ( n5678 , n812 );
buf ( n5679 , n615 );
buf ( n5680 , n438 );
buf ( n5681 , n364 );
buf ( n5682 , n1537 );
buf ( n5683 , n1488 );
buf ( n5684 , n571 );
buf ( n5685 , n950 );
buf ( n5686 , n1489 );
buf ( n5687 , n213 );
buf ( n5688 , n849 );
buf ( n5689 , n70 );
buf ( n5690 , n989 );
buf ( n5691 , n397 );
buf ( n5692 , n1039 );
buf ( n5693 , n1344 );
buf ( n5694 , n653 );
buf ( n5695 , n1115 );
buf ( n5696 , n492 );
buf ( n5697 , n1599 );
buf ( n5698 , n1894 );
buf ( n5699 , n312 );
buf ( n5700 , n1603 );
buf ( n5701 , n908 );
buf ( n5702 , n325 );
buf ( n5703 , n146 );
buf ( n5704 , n506 );
buf ( n5705 , n1498 );
buf ( n5706 , n89 );
buf ( n5707 , n1741 );
buf ( n5708 , n617 );
buf ( n5709 , n293 );
buf ( n5710 , n465 );
buf ( n5711 , n1976 );
buf ( n5712 , n1969 );
buf ( n5713 , n57 );
buf ( n5714 , n259 );
buf ( n5715 , n1236 );
buf ( n5716 , n635 );
buf ( n5717 , n1231 );
buf ( n5718 , n167 );
buf ( n5719 , n1699 );
buf ( n5720 , n948 );
buf ( n5721 , n1495 );
buf ( n5722 , n1035 );
buf ( n5723 , n1479 );
buf ( n5724 , n1994 );
buf ( n5725 , n342 );
buf ( n5726 , n182 );
buf ( n5727 , n610 );
buf ( n5728 , n1754 );
buf ( n5729 , n2015 );
buf ( n5730 , n320 );
buf ( n5731 , n1546 );
buf ( n5732 , n340 );
buf ( n5733 , n202 );
buf ( n5734 , n1453 );
buf ( n5735 , n643 );
buf ( n5736 , n1923 );
buf ( n5737 , n1962 );
buf ( n5738 , n1458 );
buf ( n5739 , n895 );
buf ( n5740 , n1947 );
buf ( n5741 , n1062 );
buf ( n5742 , n1655 );
buf ( n5743 , n385 );
buf ( n5744 , n1186 );
buf ( n5745 , n790 );
buf ( n5746 , n275 );
buf ( n5747 , n1451 );
buf ( n5748 , n652 );
buf ( n5749 , n1679 );
buf ( n5750 , n1334 );
buf ( n5751 , n404 );
buf ( n5752 , n1158 );
buf ( n5753 , n881 );
buf ( n5754 , n809 );
buf ( n5755 , n746 );
buf ( n5756 , n255 );
buf ( n5757 , n552 );
buf ( n5758 , n1011 );
buf ( n5759 , n1445 );
buf ( n5760 , n1737 );
buf ( n5761 , n1892 );
buf ( n5762 , n195 );
buf ( n5763 , n90 );
buf ( n5764 , n1595 );
buf ( n5765 , n2009 );
buf ( n5766 , n716 );
buf ( n5767 , n997 );
buf ( n5768 , n431 );
buf ( n5769 , n759 );
buf ( n5770 , n373 );
buf ( n5771 , n1471 );
buf ( n5772 , n1155 );
buf ( n5773 , n377 );
buf ( n5774 , n439 );
buf ( n5775 , n1786 );
buf ( n5776 , n669 );
buf ( n5777 , n30 );
buf ( n5778 , n355 );
buf ( n5779 , n258 );
buf ( n5780 , n1330 );
buf ( n5781 , n568 );
buf ( n5782 , n1809 );
buf ( n5783 , n559 );
buf ( n5784 , n1359 );
buf ( n5785 , n845 );
buf ( n5786 , n591 );
buf ( n5787 , n1036 );
buf ( n5788 , n1849 );
buf ( n5789 , n1468 );
buf ( n5790 , n1927 );
buf ( n5791 , n1315 );
buf ( n5792 , n640 );
buf ( n5793 , n416 );
buf ( n5794 , n1388 );
buf ( n5795 , n2012 );
buf ( n5796 , n1723 );
buf ( n5797 , n137 );
buf ( n5798 , n475 );
buf ( n5799 , n1775 );
buf ( n5800 , n205 );
buf ( n5801 , n1758 );
buf ( n5802 , n1760 );
buf ( n5803 , n8 );
buf ( n5804 , n1118 );
buf ( n5805 , n593 );
buf ( n5806 , n161 );
buf ( n5807 , n368 );
buf ( n5808 , n2026 );
buf ( n5809 , n1030 );
buf ( n5810 , n917 );
buf ( n5811 , n1756 );
buf ( n5812 , n618 );
buf ( n5813 , n1632 );
buf ( n5814 , n850 );
buf ( n5815 , n441 );
buf ( n5816 , n594 );
buf ( n5817 , n77 );
buf ( n5818 , n1753 );
buf ( n5819 , n2042 );
buf ( n5820 , n608 );
buf ( n5821 , n180 );
buf ( n5822 , n1193 );
buf ( n5823 , n395 );
buf ( n5824 , n1263 );
buf ( n5825 , n1254 );
buf ( n5826 , n1544 );
buf ( n5827 , n1805 );
buf ( n5828 , n1371 );
buf ( n5829 , n1318 );
buf ( n5830 , n1395 );
buf ( n5831 , n329 );
buf ( n5832 , n241 );
buf ( n5833 , n698 );
buf ( n5834 , n64 );
buf ( n5835 , n1059 );
buf ( n5836 , n1216 );
buf ( n5837 , n801 );
buf ( n5838 , n596 );
buf ( n5839 , n128 );
buf ( n5840 , n214 );
buf ( n5841 , n1983 );
buf ( n5842 , n1450 );
buf ( n5843 , n1665 );
buf ( n5844 , n196 );
buf ( n5845 , n1667 );
buf ( n5846 , n1618 );
buf ( n5847 , n1167 );
buf ( n5848 , n1370 );
buf ( n5849 , n510 );
buf ( n5850 , n1163 );
buf ( n5851 , n1043 );
buf ( n5852 , n1730 );
buf ( n5853 , n1089 );
buf ( n5854 , n29 );
buf ( n5855 , n1928 );
buf ( n5856 , n251 );
buf ( n5857 , n1571 );
buf ( n5858 , n2017 );
buf ( n5859 , n481 );
buf ( n5860 , n854 );
buf ( n5861 , n1324 );
buf ( n5862 , n1455 );
buf ( n5863 , n400 );
buf ( n5864 , n1143 );
buf ( n5865 , n1606 );
buf ( n5866 , n1127 );
buf ( n5867 , n1261 );
buf ( n5868 , n1624 );
buf ( n5869 , n1204 );
buf ( n5870 , n1200 );
buf ( n5871 , n1640 );
buf ( n5872 , n1176 );
buf ( n5873 , n992 );
buf ( n5874 , n560 );
buf ( n5875 , n762 );
buf ( n5876 , n1750 );
buf ( n5877 , n480 );
buf ( n5878 , n542 );
buf ( n5879 , n1749 );
buf ( n5880 , n1704 );
buf ( n5881 , n1597 );
buf ( n5882 , n1437 );
buf ( n5883 , n848 );
buf ( n5884 , n734 );
buf ( n5885 , n1967 );
buf ( n5886 , n1644 );
buf ( n5887 , n1559 );
buf ( n5888 , n1580 );
buf ( n5889 , n218 );
buf ( n5890 , n435 );
buf ( n5891 , n83 );
buf ( n5892 , n821 );
buf ( n5893 , n567 );
buf ( n5894 , n586 );
buf ( n5895 , n236 );
buf ( n5896 , n1997 );
buf ( n5897 , n1425 );
buf ( n5898 , n1979 );
buf ( n5899 , n890 );
buf ( n5900 , n1512 );
buf ( n5901 , n891 );
buf ( n5902 , n1154 );
buf ( n5903 , n1226 );
buf ( n5904 , n1861 );
buf ( n5905 , n1316 );
buf ( n5906 , n877 );
buf ( n5907 , n985 );
buf ( n5908 , n1366 );
buf ( n5909 , n749 );
buf ( n5910 , n309 );
buf ( n5911 , n1776 );
buf ( n5912 , n914 );
buf ( n5913 , n1507 );
buf ( n5914 , n1241 );
buf ( n5915 , n988 );
buf ( n5916 , n48 );
buf ( n5917 , n502 );
buf ( n5918 , n887 );
buf ( n5919 , n1383 );
buf ( n5920 , n0 );
buf ( n5921 , n1255 );
buf ( n5922 , n208 );
buf ( n5923 , n386 );
buf ( n5924 , n261 );
buf ( n5925 , n1022 );
buf ( n5926 , n360 );
buf ( n5927 , n1657 );
buf ( n5928 , n1157 );
buf ( n5929 , n1698 );
buf ( n5930 , n1533 );
buf ( n5931 , n207 );
buf ( n5932 , n232 );
buf ( n5933 , n185 );
buf ( n5934 , n883 );
buf ( n5935 , n124 );
buf ( n5936 , n1824 );
buf ( n5937 , n1474 );
buf ( n5938 , n148 );
buf ( n5939 , n578 );
buf ( n5940 , n1547 );
buf ( n5941 , n960 );
buf ( n5942 , n1960 );
buf ( n5943 , n1945 );
buf ( n5944 , n547 );
buf ( n5945 , n1658 );
buf ( n5946 , n2035 );
buf ( n5947 , n51 );
buf ( n5948 , n857 );
buf ( n5949 , n303 );
buf ( n5950 , n1816 );
buf ( n5951 , n1930 );
buf ( n5952 , n296 );
buf ( n5953 , n1057 );
buf ( n5954 , n1242 );
buf ( n5955 , n45 );
buf ( n5956 , n940 );
buf ( n5957 , n420 );
buf ( n5958 , n1578 );
buf ( n5959 , n2021 );
buf ( n5960 , n655 );
buf ( n5961 , n1407 );
buf ( n5962 , n1725 );
buf ( n5963 , n389 );
buf ( n5964 , n957 );
buf ( n5965 , n1811 );
buf ( n5966 , n1077 );
buf ( n5967 , n1392 );
buf ( n5968 , n1452 );
buf ( n5969 , n34 );
buf ( n5970 , n1536 );
buf ( n5971 , n815 );
buf ( n5972 , n170 );
buf ( n5973 , n203 );
buf ( n5974 , n1804 );
buf ( n5975 , n1239 );
buf ( n5976 , n1083 );
buf ( n5977 , n1777 );
buf ( n5978 , n688 );
buf ( n5979 , n1331 );
buf ( n5980 , n1245 );
buf ( n5981 , n737 );
buf ( n5982 , n1689 );
buf ( n5983 , n785 );
buf ( n5984 , n1694 );
buf ( n5985 , n1101 );
buf ( n5986 , n1996 );
buf ( n5987 , n1646 );
buf ( n5988 , n374 );
buf ( n5989 , n405 );
buf ( n5990 , n1562 );
buf ( n5991 , n1465 );
buf ( n5992 , n1518 );
buf ( n5993 , n519 );
buf ( n5994 , n816 );
buf ( n5995 , n1936 );
buf ( n5996 , n1856 );
buf ( n5997 , n447 );
buf ( n5998 , n1717 );
buf ( n5999 , n686 );
buf ( n6000 , n927 );
buf ( n6001 , n1159 );
buf ( n6002 , n177 );
buf ( n6003 , n1935 );
buf ( n6004 , n1007 );
buf ( n6005 , n1909 );
buf ( n6006 , n692 );
buf ( n6007 , n2008 );
buf ( n6008 , n2031 );
buf ( n6009 , n827 );
buf ( n6010 , n1882 );
buf ( n6011 , n1793 );
buf ( n6012 , n879 );
buf ( n6013 , n253 );
buf ( n6014 , n630 );
buf ( n6015 , n1883 );
buf ( n6016 , n1852 );
buf ( n6017 , n1841 );
buf ( n6018 , n712 );
buf ( n6019 , n366 );
buf ( n6020 , n1290 );
buf ( n6021 , n1807 );
buf ( n6022 , n1113 );
buf ( n6023 , n1017 );
buf ( n6024 , n974 );
buf ( n6025 , n1481 );
buf ( n6026 , n562 );
buf ( n6027 , n1237 );
buf ( n6028 , n928 );
buf ( n6029 , n194 );
buf ( n6030 , n588 );
buf ( n6031 , n174 );
buf ( n6032 , n1636 );
buf ( n6033 , n254 );
buf ( n6034 , n795 );
buf ( n6035 , n353 );
buf ( n6036 , n976 );
buf ( n6037 , n1339 );
buf ( n6038 , n449 );
buf ( n6039 , n663 );
buf ( n6040 , n198 );
buf ( n6041 , n223 );
buf ( n6042 , n152 );
buf ( n6043 , n1322 );
buf ( n6044 , n367 );
buf ( n6045 , n1296 );
buf ( n6046 , n1031 );
buf ( n6047 , n1208 );
buf ( n6048 , n344 );
buf ( n6049 , n581 );
buf ( n6050 , n819 );
buf ( n6051 , n118 );
buf ( n6052 , n1496 );
buf ( n6053 , n1047 );
buf ( n6054 , n1491 );
buf ( n6055 , n187 );
buf ( n6056 , n1633 );
buf ( n6057 , n1096 );
buf ( n6058 , n1063 );
buf ( n6059 , n1522 );
buf ( n6060 , n53 );
buf ( n6061 , n1350 );
buf ( n6062 , n1213 );
buf ( n6063 , n316 );
buf ( n6064 , n1995 );
buf ( n6065 , n1677 );
buf ( n6066 , n1280 );
buf ( n6067 , n1404 );
buf ( n6068 , n1251 );
buf ( n6069 , n1904 );
buf ( n6070 , n273 );
buf ( n6071 , n792 );
buf ( n6072 , n15 );
buf ( n6073 , n1149 );
buf ( n6074 , n294 );
buf ( n6075 , n338 );
buf ( n6076 , n544 );
buf ( n6077 , n1702 );
buf ( n6078 , n893 );
buf ( n6079 , n1076 );
buf ( n6080 , n1310 );
buf ( n6081 , n193 );
buf ( n6082 , n1855 );
buf ( n6083 , n412 );
buf ( n6084 , n1803 );
buf ( n6085 , n1833 );
buf ( n6086 , n469 );
buf ( n6087 , n1214 );
buf ( n6088 , n804 );
buf ( n6089 , n1864 );
buf ( n6090 , n1586 );
buf ( n6091 , n672 );
buf ( n6092 , n776 );
buf ( n6093 , n162 );
buf ( n6094 , n826 );
buf ( n6095 , n470 );
buf ( n6096 , n1605 );
buf ( n6097 , n347 );
buf ( n6098 , n732 );
buf ( n6099 , n1937 );
buf ( n6100 , n114 );
buf ( n6101 , n528 );
buf ( n6102 , n262 );
buf ( n6103 , n897 );
buf ( n6104 , n791 );
buf ( n6105 , n840 );
buf ( n6106 , n1834 );
buf ( n6107 , n1287 );
buf ( n6108 , n2038 );
buf ( n6109 , n1572 );
buf ( n6110 , n244 );
buf ( n6111 , n345 );
buf ( n6112 , n1023 );
buf ( n6113 , n1195 );
buf ( n6114 , n1397 );
buf ( n6115 , n1738 );
buf ( n6116 , n1408 );
buf ( n6117 , n1801 );
buf ( n6118 , n1933 );
buf ( n6119 , n1903 );
buf ( n6120 , n537 );
buf ( n6121 , n726 );
buf ( n6122 , n638 );
buf ( n6123 , n419 );
buf ( n6124 , n611 );
buf ( n6125 , n744 );
buf ( n6126 , n723 );
buf ( n6127 , n1916 );
buf ( n6128 , n600 );
buf ( n6129 , n1212 );
buf ( n6130 , n1146 );
buf ( n6131 , n9 );
buf ( n6132 , n314 );
buf ( n6133 , n290 );
buf ( n6134 , n677 );
buf ( n6135 , n300 );
buf ( n6136 , n952 );
buf ( n6137 , n1806 );
buf ( n6138 , n1342 );
buf ( n6139 , n1998 );
buf ( n6140 , n285 );
buf ( n6141 , n1716 );
buf ( n6142 , n2046 );
buf ( n6143 , n1112 );
buf ( n6144 , n645 );
buf ( n6145 , n1441 );
buf ( n6146 , n18 );
buf ( n6147 , n1561 );
buf ( n6148 , n19 );
buf ( n6149 , n1551 );
not ( n6150 , n5155 );
not ( n6151 , n4131 );
or ( n6152 , n6150 , n6151 );
or ( n6153 , n4131 , n5155 );
nand ( n6154 , n6152 , n6153 );
not ( n6155 , n5154 );
not ( n6156 , n4130 );
or ( n6157 , n6155 , n6156 );
or ( n6158 , n4130 , n5154 );
nand ( n6159 , n6157 , n6158 );
nand ( n6160 , n6154 , n6159 );
not ( n6161 , n5157 );
not ( n6162 , n4133 );
or ( n6163 , n6161 , n6162 );
or ( n6164 , n4133 , n5157 );
nand ( n6165 , n6163 , n6164 );
not ( n6166 , n5156 );
not ( n6167 , n4132 );
or ( n6168 , n6166 , n6167 );
or ( n6169 , n4132 , n5156 );
nand ( n6170 , n6168 , n6169 );
nand ( n6171 , n6165 , n6170 );
nor ( n6172 , n6160 , n6171 );
not ( n6173 , n5151 );
not ( n6174 , n4127 );
or ( n6175 , n6173 , n6174 );
or ( n6176 , n4127 , n5151 );
nand ( n6177 , n6175 , n6176 );
not ( n6178 , n5150 );
not ( n6179 , n4126 );
or ( n6180 , n6178 , n6179 );
or ( n6181 , n4126 , n5150 );
nand ( n6182 , n6180 , n6181 );
nand ( n6183 , n6177 , n6182 );
not ( n6184 , n5153 );
not ( n6185 , n4129 );
or ( n6186 , n6184 , n6185 );
or ( n6187 , n4129 , n5153 );
nand ( n6188 , n6186 , n6187 );
not ( n6189 , n5152 );
not ( n6190 , n4128 );
or ( n6191 , n6189 , n6190 );
or ( n6192 , n4128 , n5152 );
nand ( n6193 , n6191 , n6192 );
nand ( n6194 , n6188 , n6193 );
nor ( n6195 , n6183 , n6194 );
not ( n6196 , n5147 );
not ( n6197 , n4123 );
or ( n6198 , n6196 , n6197 );
or ( n6199 , n4123 , n5147 );
nand ( n6200 , n6198 , n6199 );
not ( n6201 , n5146 );
not ( n6202 , n4122 );
or ( n6203 , n6201 , n6202 );
or ( n6204 , n4122 , n5146 );
nand ( n6205 , n6203 , n6204 );
nand ( n6206 , n6200 , n6205 );
not ( n6207 , n5149 );
not ( n6208 , n4125 );
or ( n6209 , n6207 , n6208 );
or ( n6210 , n4125 , n5149 );
nand ( n6211 , n6209 , n6210 );
not ( n6212 , n5148 );
not ( n6213 , n4124 );
or ( n6214 , n6212 , n6213 );
or ( n6215 , n4124 , n5148 );
nand ( n6216 , n6214 , n6215 );
nand ( n6217 , n6211 , n6216 );
nor ( n6218 , n6206 , n6217 );
not ( n6219 , n5143 );
not ( n6220 , n4119 );
or ( n6221 , n6219 , n6220 );
or ( n6222 , n4119 , n5143 );
nand ( n6223 , n6221 , n6222 );
not ( n6224 , n5142 );
not ( n6225 , n4118 );
or ( n6226 , n6224 , n6225 );
or ( n6227 , n4118 , n5142 );
nand ( n6228 , n6226 , n6227 );
nand ( n6229 , n6223 , n6228 );
not ( n6230 , n5145 );
not ( n6231 , n4121 );
or ( n6232 , n6230 , n6231 );
or ( n6233 , n4121 , n5145 );
nand ( n6234 , n6232 , n6233 );
not ( n6235 , n5144 );
not ( n6236 , n4120 );
or ( n6237 , n6235 , n6236 );
or ( n6238 , n4120 , n5144 );
nand ( n6239 , n6237 , n6238 );
nand ( n6240 , n6234 , n6239 );
nor ( n6241 , n6229 , n6240 );
nand ( n6242 , n6172 , n6195 , n6218 , n6241 );
not ( n6243 , n5139 );
not ( n6244 , n4115 );
or ( n6245 , n6243 , n6244 );
or ( n6246 , n4115 , n5139 );
nand ( n6247 , n6245 , n6246 );
not ( n6248 , n5138 );
not ( n6249 , n4114 );
or ( n6250 , n6248 , n6249 );
or ( n6251 , n4114 , n5138 );
nand ( n6252 , n6250 , n6251 );
nand ( n6253 , n6247 , n6252 );
not ( n6254 , n5141 );
not ( n6255 , n4117 );
or ( n6256 , n6254 , n6255 );
or ( n6257 , n4117 , n5141 );
nand ( n6258 , n6256 , n6257 );
not ( n6259 , n5140 );
not ( n6260 , n4116 );
or ( n6261 , n6259 , n6260 );
or ( n6262 , n4116 , n5140 );
nand ( n6263 , n6261 , n6262 );
nand ( n6264 , n6258 , n6263 );
nor ( n6265 , n6253 , n6264 );
not ( n6266 , n5135 );
not ( n6267 , n4111 );
or ( n6268 , n6266 , n6267 );
or ( n6269 , n4111 , n5135 );
nand ( n6270 , n6268 , n6269 );
not ( n6271 , n5134 );
not ( n6272 , n4110 );
or ( n6273 , n6271 , n6272 );
or ( n6274 , n4110 , n5134 );
nand ( n6275 , n6273 , n6274 );
nand ( n6276 , n6270 , n6275 );
not ( n6277 , n5137 );
not ( n6278 , n4113 );
or ( n6279 , n6277 , n6278 );
or ( n6280 , n4113 , n5137 );
nand ( n6281 , n6279 , n6280 );
not ( n6282 , n5136 );
not ( n6283 , n4112 );
or ( n6284 , n6282 , n6283 );
or ( n6285 , n4112 , n5136 );
nand ( n6286 , n6284 , n6285 );
nand ( n6287 , n6281 , n6286 );
nor ( n6288 , n6276 , n6287 );
not ( n6289 , n5131 );
not ( n6290 , n4107 );
or ( n6291 , n6289 , n6290 );
or ( n6292 , n4107 , n5131 );
nand ( n6293 , n6291 , n6292 );
not ( n6294 , n5130 );
not ( n6295 , n4106 );
or ( n6296 , n6294 , n6295 );
or ( n6297 , n4106 , n5130 );
nand ( n6298 , n6296 , n6297 );
nand ( n6299 , n6293 , n6298 );
not ( n6300 , n5133 );
not ( n6301 , n4109 );
or ( n6302 , n6300 , n6301 );
or ( n6303 , n4109 , n5133 );
nand ( n6304 , n6302 , n6303 );
not ( n6305 , n5132 );
not ( n6306 , n4108 );
or ( n6307 , n6305 , n6306 );
or ( n6308 , n4108 , n5132 );
nand ( n6309 , n6307 , n6308 );
nand ( n6310 , n6304 , n6309 );
nor ( n6311 , n6299 , n6310 );
not ( n6312 , n5127 );
not ( n6313 , n4103 );
or ( n6314 , n6312 , n6313 );
or ( n6315 , n4103 , n5127 );
nand ( n6316 , n6314 , n6315 );
not ( n6317 , n5126 );
not ( n6318 , n4102 );
or ( n6319 , n6317 , n6318 );
or ( n6320 , n4102 , n5126 );
nand ( n6321 , n6319 , n6320 );
nand ( n6322 , n6316 , n6321 );
not ( n6323 , n5129 );
not ( n6324 , n4105 );
or ( n6325 , n6323 , n6324 );
or ( n6326 , n4105 , n5129 );
nand ( n6327 , n6325 , n6326 );
not ( n6328 , n5128 );
not ( n6329 , n4104 );
or ( n6330 , n6328 , n6329 );
or ( n6331 , n4104 , n5128 );
nand ( n6332 , n6330 , n6331 );
nand ( n6333 , n6327 , n6332 );
nor ( n6334 , n6322 , n6333 );
nand ( n6335 , n6265 , n6288 , n6311 , n6334 );
nor ( n6336 , n6242 , n6335 );
not ( n6337 , n5171 );
not ( n6338 , n4147 );
or ( n6339 , n6337 , n6338 );
or ( n6340 , n4147 , n5171 );
nand ( n6341 , n6339 , n6340 );
not ( n6342 , n5172 );
not ( n6343 , n4148 );
or ( n6344 , n6342 , n6343 );
or ( n6345 , n4148 , n5172 );
nand ( n6346 , n6344 , n6345 );
not ( n6347 , n5173 );
not ( n6348 , n4149 );
or ( n6349 , n6347 , n6348 );
or ( n6350 , n4149 , n5173 );
nand ( n6351 , n6349 , n6350 );
not ( n6352 , n5170 );
not ( n6353 , n4146 );
or ( n6354 , n6352 , n6353 );
or ( n6355 , n4146 , n5170 );
nand ( n6356 , n6354 , n6355 );
and ( n6357 , n6341 , n6346 , n6351 , n6356 );
not ( n6358 , n5167 );
not ( n6359 , n4143 );
or ( n6360 , n6358 , n6359 );
or ( n6361 , n4143 , n5167 );
nand ( n6362 , n6360 , n6361 );
not ( n6363 , n5166 );
not ( n6364 , n4142 );
or ( n6365 , n6363 , n6364 );
or ( n6366 , n4142 , n5166 );
nand ( n6367 , n6365 , n6366 );
nand ( n6368 , n6362 , n6367 );
not ( n6369 , n5169 );
not ( n6370 , n4145 );
or ( n6371 , n6369 , n6370 );
or ( n6372 , n4145 , n5169 );
nand ( n6373 , n6371 , n6372 );
not ( n6374 , n5168 );
not ( n6375 , n4144 );
or ( n6376 , n6374 , n6375 );
or ( n6377 , n4144 , n5168 );
nand ( n6378 , n6376 , n6377 );
nand ( n6379 , n6373 , n6378 );
nor ( n6380 , n6368 , n6379 );
not ( n6381 , n5159 );
not ( n6382 , n4135 );
or ( n6383 , n6381 , n6382 );
or ( n6384 , n4135 , n5159 );
nand ( n6385 , n6383 , n6384 );
not ( n6386 , n5158 );
not ( n6387 , n4134 );
or ( n6388 , n6386 , n6387 );
or ( n6389 , n4134 , n5158 );
nand ( n6390 , n6388 , n6389 );
nand ( n6391 , n6385 , n6390 );
not ( n6392 , n5161 );
not ( n6393 , n4137 );
or ( n6394 , n6392 , n6393 );
or ( n6395 , n4137 , n5161 );
nand ( n6396 , n6394 , n6395 );
not ( n6397 , n5160 );
not ( n6398 , n4136 );
or ( n6399 , n6397 , n6398 );
or ( n6400 , n4136 , n5160 );
nand ( n6401 , n6399 , n6400 );
nand ( n6402 , n6396 , n6401 );
nor ( n6403 , n6391 , n6402 );
not ( n6404 , n5165 );
not ( n6405 , n4141 );
or ( n6406 , n6404 , n6405 );
or ( n6407 , n4141 , n5165 );
nand ( n6408 , n6406 , n6407 );
not ( n6409 , n5164 );
not ( n6410 , n4140 );
or ( n6411 , n6409 , n6410 );
or ( n6412 , n4140 , n5164 );
nand ( n6413 , n6411 , n6412 );
nand ( n6414 , n6408 , n6413 );
not ( n6415 , n5163 );
not ( n6416 , n4139 );
or ( n6417 , n6415 , n6416 );
or ( n6418 , n4139 , n5163 );
nand ( n6419 , n6417 , n6418 );
not ( n6420 , n5162 );
not ( n6421 , n4138 );
or ( n6422 , n6420 , n6421 );
or ( n6423 , n4138 , n5162 );
nand ( n6424 , n6422 , n6423 );
nand ( n6425 , n6419 , n6424 );
nor ( n6426 , n6414 , n6425 );
nand ( n6427 , n6357 , n6380 , n6403 , n6426 );
not ( n6428 , n5187 );
not ( n6429 , n4163 );
or ( n6430 , n6428 , n6429 );
or ( n6431 , n4163 , n5187 );
nand ( n6432 , n6430 , n6431 );
not ( n6433 , n5186 );
not ( n6434 , n4162 );
or ( n6435 , n6433 , n6434 );
or ( n6436 , n4162 , n5186 );
nand ( n6437 , n6435 , n6436 );
nand ( n6438 , n6432 , n6437 );
not ( n6439 , n5189 );
not ( n6440 , n4165 );
or ( n6441 , n6439 , n6440 );
or ( n6442 , n4165 , n5189 );
nand ( n6443 , n6441 , n6442 );
not ( n6444 , n5188 );
not ( n6445 , n4164 );
or ( n6446 , n6444 , n6445 );
or ( n6447 , n4164 , n5188 );
nand ( n6448 , n6446 , n6447 );
nand ( n6449 , n6443 , n6448 );
nor ( n6450 , n6438 , n6449 );
not ( n6451 , n5183 );
not ( n6452 , n4159 );
or ( n6453 , n6451 , n6452 );
or ( n6454 , n4159 , n5183 );
nand ( n6455 , n6453 , n6454 );
not ( n6456 , n5182 );
not ( n6457 , n4158 );
or ( n6458 , n6456 , n6457 );
or ( n6459 , n4158 , n5182 );
nand ( n6460 , n6458 , n6459 );
nand ( n6461 , n6455 , n6460 );
not ( n6462 , n5185 );
not ( n6463 , n4161 );
or ( n6464 , n6462 , n6463 );
or ( n6465 , n4161 , n5185 );
nand ( n6466 , n6464 , n6465 );
not ( n6467 , n5184 );
not ( n6468 , n4160 );
or ( n6469 , n6467 , n6468 );
or ( n6470 , n4160 , n5184 );
nand ( n6471 , n6469 , n6470 );
nand ( n6472 , n6466 , n6471 );
nor ( n6473 , n6461 , n6472 );
not ( n6474 , n5179 );
not ( n6475 , n4155 );
or ( n6476 , n6474 , n6475 );
or ( n6477 , n4155 , n5179 );
nand ( n6478 , n6476 , n6477 );
not ( n6479 , n5178 );
not ( n6480 , n4154 );
or ( n6481 , n6479 , n6480 );
or ( n6482 , n4154 , n5178 );
nand ( n6483 , n6481 , n6482 );
nand ( n6484 , n6478 , n6483 );
not ( n6485 , n5181 );
not ( n6486 , n4157 );
or ( n6487 , n6485 , n6486 );
or ( n6488 , n4157 , n5181 );
nand ( n6489 , n6487 , n6488 );
not ( n6490 , n5180 );
not ( n6491 , n4156 );
or ( n6492 , n6490 , n6491 );
or ( n6493 , n4156 , n5180 );
nand ( n6494 , n6492 , n6493 );
nand ( n6495 , n6489 , n6494 );
nor ( n6496 , n6484 , n6495 );
not ( n6497 , n5175 );
not ( n6498 , n4151 );
or ( n6499 , n6497 , n6498 );
or ( n6500 , n4151 , n5175 );
nand ( n6501 , n6499 , n6500 );
not ( n6502 , n5174 );
not ( n6503 , n4150 );
or ( n6504 , n6502 , n6503 );
or ( n6505 , n4150 , n5174 );
nand ( n6506 , n6504 , n6505 );
nand ( n6507 , n6501 , n6506 );
not ( n6508 , n5177 );
not ( n6509 , n4153 );
or ( n6510 , n6508 , n6509 );
or ( n6511 , n4153 , n5177 );
nand ( n6512 , n6510 , n6511 );
not ( n6513 , n5176 );
not ( n6514 , n4152 );
or ( n6515 , n6513 , n6514 );
or ( n6516 , n4152 , n5176 );
nand ( n6517 , n6515 , n6516 );
nand ( n6518 , n6512 , n6517 );
nor ( n6519 , n6507 , n6518 );
nand ( n6520 , n6450 , n6473 , n6496 , n6519 );
nor ( n6521 , n6427 , n6520 );
not ( n6522 , n5192 );
not ( n6523 , n4168 );
or ( n6524 , n6522 , n6523 );
or ( n6525 , n4168 , n5192 );
nand ( n6526 , n6524 , n6525 );
not ( n6527 , n5193 );
not ( n6528 , n4169 );
or ( n6529 , n6527 , n6528 );
or ( n6530 , n4169 , n5193 );
nand ( n6531 , n6529 , n6530 );
not ( n6532 , n5190 );
not ( n6533 , n4166 );
or ( n6534 , n6532 , n6533 );
or ( n6535 , n4166 , n5190 );
nand ( n6536 , n6534 , n6535 );
not ( n6537 , n5191 );
not ( n6538 , n4167 );
or ( n6539 , n6537 , n6538 );
or ( n6540 , n4167 , n5191 );
nand ( n6541 , n6539 , n6540 );
nand ( n6542 , n6526 , n6531 , n6536 , n6541 );
not ( n6543 , n5203 );
not ( n6544 , n4179 );
or ( n6545 , n6543 , n6544 );
or ( n6546 , n4179 , n5203 );
nand ( n6547 , n6545 , n6546 );
not ( n6548 , n5205 );
not ( n6549 , n4181 );
or ( n6550 , n6548 , n6549 );
or ( n6551 , n4181 , n5205 );
nand ( n6552 , n6550 , n6551 );
not ( n6553 , n5202 );
not ( n6554 , n4178 );
or ( n6555 , n6553 , n6554 );
or ( n6556 , n4178 , n5202 );
nand ( n6557 , n6555 , n6556 );
not ( n6558 , n5204 );
not ( n6559 , n4180 );
or ( n6560 , n6558 , n6559 );
or ( n6561 , n4180 , n5204 );
nand ( n6562 , n6560 , n6561 );
nand ( n6563 , n6547 , n6552 , n6557 , n6562 );
nor ( n6564 , n6542 , n6563 );
not ( n6565 , n5200 );
not ( n6566 , n4176 );
or ( n6567 , n6565 , n6566 );
or ( n6568 , n4176 , n5200 );
nand ( n6569 , n6567 , n6568 );
not ( n6570 , n5201 );
not ( n6571 , n4177 );
or ( n6572 , n6570 , n6571 );
or ( n6573 , n4177 , n5201 );
nand ( n6574 , n6572 , n6573 );
not ( n6575 , n5198 );
not ( n6576 , n4174 );
or ( n6577 , n6575 , n6576 );
or ( n6578 , n4174 , n5198 );
nand ( n6579 , n6577 , n6578 );
not ( n6580 , n5199 );
not ( n6581 , n4175 );
or ( n6582 , n6580 , n6581 );
or ( n6583 , n4175 , n5199 );
nand ( n6584 , n6582 , n6583 );
nand ( n6585 , n6569 , n6574 , n6579 , n6584 );
not ( n6586 , n4172 );
not ( n6587 , n5196 );
or ( n6588 , n6586 , n6587 );
or ( n6589 , n5196 , n4172 );
nand ( n6590 , n6588 , n6589 );
not ( n6591 , n4173 );
not ( n6592 , n5197 );
or ( n6593 , n6591 , n6592 );
or ( n6594 , n5197 , n4173 );
nand ( n6595 , n6593 , n6594 );
not ( n6596 , n4170 );
not ( n6597 , n5194 );
or ( n6598 , n6596 , n6597 );
or ( n6599 , n5194 , n4170 );
nand ( n6600 , n6598 , n6599 );
not ( n6601 , n4171 );
not ( n6602 , n5195 );
or ( n6603 , n6601 , n6602 );
or ( n6604 , n5195 , n4171 );
nand ( n6605 , n6603 , n6604 );
nand ( n6606 , n6590 , n6595 , n6600 , n6605 );
nor ( n6607 , n6585 , n6606 );
nand ( n6608 , n6564 , n6607 );
not ( n6609 , n5215 );
not ( n6610 , n4191 );
or ( n6611 , n6609 , n6610 );
or ( n6612 , n4191 , n5215 );
nand ( n6613 , n6611 , n6612 );
not ( n6614 , n5214 );
not ( n6615 , n4190 );
or ( n6616 , n6614 , n6615 );
or ( n6617 , n4190 , n5214 );
nand ( n6618 , n6616 , n6617 );
nand ( n6619 , n6613 , n6618 );
not ( n6620 , n5217 );
not ( n6621 , n4193 );
or ( n6622 , n6620 , n6621 );
or ( n6623 , n4193 , n5217 );
nand ( n6624 , n6622 , n6623 );
not ( n6625 , n5216 );
not ( n6626 , n4192 );
or ( n6627 , n6625 , n6626 );
or ( n6628 , n4192 , n5216 );
nand ( n6629 , n6627 , n6628 );
nand ( n6630 , n6624 , n6629 );
nor ( n6631 , n6619 , n6630 );
not ( n6632 , n5211 );
not ( n6633 , n4187 );
or ( n6634 , n6632 , n6633 );
or ( n6635 , n4187 , n5211 );
nand ( n6636 , n6634 , n6635 );
not ( n6637 , n5210 );
not ( n6638 , n4186 );
or ( n6639 , n6637 , n6638 );
or ( n6640 , n4186 , n5210 );
nand ( n6641 , n6639 , n6640 );
nand ( n6642 , n6636 , n6641 );
not ( n6643 , n5213 );
not ( n6644 , n4189 );
or ( n6645 , n6643 , n6644 );
or ( n6646 , n4189 , n5213 );
nand ( n6647 , n6645 , n6646 );
not ( n6648 , n5212 );
not ( n6649 , n4188 );
or ( n6650 , n6648 , n6649 );
or ( n6651 , n4188 , n5212 );
nand ( n6652 , n6650 , n6651 );
nand ( n6653 , n6647 , n6652 );
nor ( n6654 , n6642 , n6653 );
not ( n6655 , n5220 );
not ( n6656 , n4196 );
or ( n6657 , n6655 , n6656 );
or ( n6658 , n4196 , n5220 );
nand ( n6659 , n6657 , n6658 );
not ( n6660 , n5221 );
not ( n6661 , n4197 );
or ( n6662 , n6660 , n6661 );
or ( n6663 , n4197 , n5221 );
nand ( n6664 , n6662 , n6663 );
not ( n6665 , n5218 );
not ( n6666 , n4194 );
or ( n6667 , n6665 , n6666 );
or ( n6668 , n4194 , n5218 );
nand ( n6669 , n6667 , n6668 );
not ( n6670 , n5219 );
not ( n6671 , n4195 );
or ( n6672 , n6670 , n6671 );
or ( n6673 , n4195 , n5219 );
nand ( n6674 , n6672 , n6673 );
nand ( n6675 , n6659 , n6664 , n6669 , n6674 );
not ( n6676 , n6675 );
not ( n6677 , n5207 );
not ( n6678 , n4183 );
or ( n6679 , n6677 , n6678 );
or ( n6680 , n4183 , n5207 );
nand ( n6681 , n6679 , n6680 );
not ( n6682 , n5206 );
not ( n6683 , n4182 );
or ( n6684 , n6682 , n6683 );
or ( n6685 , n4182 , n5206 );
nand ( n6686 , n6684 , n6685 );
nand ( n6687 , n6681 , n6686 );
not ( n6688 , n5209 );
not ( n6689 , n4185 );
or ( n6690 , n6688 , n6689 );
or ( n6691 , n4185 , n5209 );
nand ( n6692 , n6690 , n6691 );
not ( n6693 , n5208 );
not ( n6694 , n4184 );
or ( n6695 , n6693 , n6694 );
or ( n6696 , n4184 , n5208 );
nand ( n6697 , n6695 , n6696 );
nand ( n6698 , n6692 , n6697 );
nor ( n6699 , n6687 , n6698 );
nand ( n6700 , n6631 , n6654 , n6676 , n6699 );
nor ( n6701 , n6608 , n6700 );
not ( n6702 , n5235 );
not ( n6703 , n4211 );
or ( n6704 , n6702 , n6703 );
or ( n6705 , n4211 , n5235 );
nand ( n6706 , n6704 , n6705 );
not ( n6707 , n5234 );
not ( n6708 , n4210 );
or ( n6709 , n6707 , n6708 );
or ( n6710 , n4210 , n5234 );
nand ( n6711 , n6709 , n6710 );
nand ( n6712 , n6706 , n6711 );
not ( n6713 , n5237 );
not ( n6714 , n4213 );
or ( n6715 , n6713 , n6714 );
or ( n6716 , n4213 , n5237 );
nand ( n6717 , n6715 , n6716 );
not ( n6718 , n5236 );
not ( n6719 , n4212 );
or ( n6720 , n6718 , n6719 );
or ( n6721 , n4212 , n5236 );
nand ( n6722 , n6720 , n6721 );
nand ( n6723 , n6717 , n6722 );
nor ( n6724 , n6712 , n6723 );
not ( n6725 , n5231 );
not ( n6726 , n4207 );
or ( n6727 , n6725 , n6726 );
or ( n6728 , n4207 , n5231 );
nand ( n6729 , n6727 , n6728 );
not ( n6730 , n5230 );
not ( n6731 , n4206 );
or ( n6732 , n6730 , n6731 );
or ( n6733 , n4206 , n5230 );
nand ( n6734 , n6732 , n6733 );
nand ( n6735 , n6729 , n6734 );
not ( n6736 , n5233 );
not ( n6737 , n4209 );
or ( n6738 , n6736 , n6737 );
or ( n6739 , n4209 , n5233 );
nand ( n6740 , n6738 , n6739 );
not ( n6741 , n5232 );
not ( n6742 , n4208 );
or ( n6743 , n6741 , n6742 );
or ( n6744 , n4208 , n5232 );
nand ( n6745 , n6743 , n6744 );
nand ( n6746 , n6740 , n6745 );
nor ( n6747 , n6735 , n6746 );
not ( n6748 , n5227 );
not ( n6749 , n4203 );
or ( n6750 , n6748 , n6749 );
or ( n6751 , n4203 , n5227 );
nand ( n6752 , n6750 , n6751 );
not ( n6753 , n5226 );
not ( n6754 , n4202 );
or ( n6755 , n6753 , n6754 );
or ( n6756 , n4202 , n5226 );
nand ( n6757 , n6755 , n6756 );
nand ( n6758 , n6752 , n6757 );
not ( n6759 , n5229 );
not ( n6760 , n4205 );
or ( n6761 , n6759 , n6760 );
or ( n6762 , n4205 , n5229 );
nand ( n6763 , n6761 , n6762 );
not ( n6764 , n5228 );
not ( n6765 , n4204 );
or ( n6766 , n6764 , n6765 );
or ( n6767 , n4204 , n5228 );
nand ( n6768 , n6766 , n6767 );
nand ( n6769 , n6763 , n6768 );
nor ( n6770 , n6758 , n6769 );
not ( n6771 , n5223 );
not ( n6772 , n4199 );
or ( n6773 , n6771 , n6772 );
or ( n6774 , n4199 , n5223 );
nand ( n6775 , n6773 , n6774 );
not ( n6776 , n5222 );
not ( n6777 , n4198 );
or ( n6778 , n6776 , n6777 );
or ( n6779 , n4198 , n5222 );
nand ( n6780 , n6778 , n6779 );
nand ( n6781 , n6775 , n6780 );
not ( n6782 , n5225 );
not ( n6783 , n4201 );
or ( n6784 , n6782 , n6783 );
or ( n6785 , n4201 , n5225 );
nand ( n6786 , n6784 , n6785 );
not ( n6787 , n5224 );
not ( n6788 , n4200 );
or ( n6789 , n6787 , n6788 );
or ( n6790 , n4200 , n5224 );
nand ( n6791 , n6789 , n6790 );
nand ( n6792 , n6786 , n6791 );
nor ( n6793 , n6781 , n6792 );
nand ( n6794 , n6724 , n6747 , n6770 , n6793 );
not ( n6795 , n5251 );
not ( n6796 , n4227 );
or ( n6797 , n6795 , n6796 );
or ( n6798 , n4227 , n5251 );
nand ( n6799 , n6797 , n6798 );
not ( n6800 , n5250 );
not ( n6801 , n4226 );
or ( n6802 , n6800 , n6801 );
or ( n6803 , n4226 , n5250 );
nand ( n6804 , n6802 , n6803 );
nand ( n6805 , n6799 , n6804 );
not ( n6806 , n5253 );
not ( n6807 , n4229 );
or ( n6808 , n6806 , n6807 );
or ( n6809 , n4229 , n5253 );
nand ( n6810 , n6808 , n6809 );
not ( n6811 , n5252 );
not ( n6812 , n4228 );
or ( n6813 , n6811 , n6812 );
or ( n6814 , n4228 , n5252 );
nand ( n6815 , n6813 , n6814 );
nand ( n6816 , n6810 , n6815 );
nor ( n6817 , n6805 , n6816 );
not ( n6818 , n5247 );
not ( n6819 , n4223 );
or ( n6820 , n6818 , n6819 );
or ( n6821 , n4223 , n5247 );
nand ( n6822 , n6820 , n6821 );
not ( n6823 , n5246 );
not ( n6824 , n4222 );
or ( n6825 , n6823 , n6824 );
or ( n6826 , n4222 , n5246 );
nand ( n6827 , n6825 , n6826 );
nand ( n6828 , n6822 , n6827 );
not ( n6829 , n5249 );
not ( n6830 , n4225 );
or ( n6831 , n6829 , n6830 );
or ( n6832 , n4225 , n5249 );
nand ( n6833 , n6831 , n6832 );
not ( n6834 , n5248 );
not ( n6835 , n4224 );
or ( n6836 , n6834 , n6835 );
or ( n6837 , n4224 , n5248 );
nand ( n6838 , n6836 , n6837 );
nand ( n6839 , n6833 , n6838 );
nor ( n6840 , n6828 , n6839 );
not ( n6841 , n5243 );
not ( n6842 , n4219 );
or ( n6843 , n6841 , n6842 );
or ( n6844 , n4219 , n5243 );
nand ( n6845 , n6843 , n6844 );
not ( n6846 , n5242 );
not ( n6847 , n4218 );
or ( n6848 , n6846 , n6847 );
or ( n6849 , n4218 , n5242 );
nand ( n6850 , n6848 , n6849 );
nand ( n6851 , n6845 , n6850 );
not ( n6852 , n5245 );
not ( n6853 , n4221 );
or ( n6854 , n6852 , n6853 );
or ( n6855 , n4221 , n5245 );
nand ( n6856 , n6854 , n6855 );
not ( n6857 , n5244 );
not ( n6858 , n4220 );
or ( n6859 , n6857 , n6858 );
or ( n6860 , n4220 , n5244 );
nand ( n6861 , n6859 , n6860 );
nand ( n6862 , n6856 , n6861 );
nor ( n6863 , n6851 , n6862 );
not ( n6864 , n5239 );
not ( n6865 , n4215 );
or ( n6866 , n6864 , n6865 );
or ( n6867 , n4215 , n5239 );
nand ( n6868 , n6866 , n6867 );
not ( n6869 , n5238 );
not ( n6870 , n4214 );
or ( n6871 , n6869 , n6870 );
or ( n6872 , n4214 , n5238 );
nand ( n6873 , n6871 , n6872 );
nand ( n6874 , n6868 , n6873 );
not ( n6875 , n5241 );
not ( n6876 , n4217 );
or ( n6877 , n6875 , n6876 );
or ( n6878 , n4217 , n5241 );
nand ( n6879 , n6877 , n6878 );
not ( n6880 , n5240 );
not ( n6881 , n4216 );
or ( n6882 , n6880 , n6881 );
or ( n6883 , n4216 , n5240 );
nand ( n6884 , n6882 , n6883 );
nand ( n6885 , n6879 , n6884 );
nor ( n6886 , n6874 , n6885 );
nand ( n6887 , n6817 , n6840 , n6863 , n6886 );
nor ( n6888 , n6794 , n6887 );
nand ( n6889 , n6336 , n6521 , n6701 , n6888 );
not ( n6890 , n5263 );
not ( n6891 , n4239 );
or ( n6892 , n6890 , n6891 );
or ( n6893 , n4239 , n5263 );
nand ( n6894 , n6892 , n6893 );
not ( n6895 , n5262 );
not ( n6896 , n4238 );
or ( n6897 , n6895 , n6896 );
or ( n6898 , n4238 , n5262 );
nand ( n6899 , n6897 , n6898 );
nand ( n6900 , n6894 , n6899 );
not ( n6901 , n5265 );
not ( n6902 , n4241 );
or ( n6903 , n6901 , n6902 );
or ( n6904 , n4241 , n5265 );
nand ( n6905 , n6903 , n6904 );
not ( n6906 , n5264 );
not ( n6907 , n4240 );
or ( n6908 , n6906 , n6907 );
or ( n6909 , n4240 , n5264 );
nand ( n6910 , n6908 , n6909 );
nand ( n6911 , n6905 , n6910 );
nor ( n6912 , n6900 , n6911 );
not ( n6913 , n5267 );
not ( n6914 , n4243 );
or ( n6915 , n6913 , n6914 );
or ( n6916 , n4243 , n5267 );
nand ( n6917 , n6915 , n6916 );
not ( n6918 , n5266 );
not ( n6919 , n4242 );
or ( n6920 , n6918 , n6919 );
or ( n6921 , n4242 , n5266 );
nand ( n6922 , n6920 , n6921 );
nand ( n6923 , n6917 , n6922 );
not ( n6924 , n5269 );
not ( n6925 , n4245 );
or ( n6926 , n6924 , n6925 );
or ( n6927 , n4245 , n5269 );
nand ( n6928 , n6926 , n6927 );
not ( n6929 , n5268 );
not ( n6930 , n4244 );
or ( n6931 , n6929 , n6930 );
or ( n6932 , n4244 , n5268 );
nand ( n6933 , n6931 , n6932 );
nand ( n6934 , n6928 , n6933 );
nor ( n6935 , n6923 , n6934 );
not ( n6936 , n5259 );
not ( n6937 , n4235 );
or ( n6938 , n6936 , n6937 );
or ( n6939 , n4235 , n5259 );
nand ( n6940 , n6938 , n6939 );
not ( n6941 , n5258 );
not ( n6942 , n4234 );
or ( n6943 , n6941 , n6942 );
or ( n6944 , n4234 , n5258 );
nand ( n6945 , n6943 , n6944 );
nand ( n6946 , n6940 , n6945 );
not ( n6947 , n5261 );
not ( n6948 , n4237 );
or ( n6949 , n6947 , n6948 );
or ( n6950 , n4237 , n5261 );
nand ( n6951 , n6949 , n6950 );
not ( n6952 , n5260 );
not ( n6953 , n4236 );
or ( n6954 , n6952 , n6953 );
or ( n6955 , n4236 , n5260 );
nand ( n6956 , n6954 , n6955 );
nand ( n6957 , n6951 , n6956 );
nor ( n6958 , n6946 , n6957 );
not ( n6959 , n5257 );
not ( n6960 , n4233 );
or ( n6961 , n6959 , n6960 );
or ( n6962 , n4233 , n5257 );
nand ( n6963 , n6961 , n6962 );
not ( n6964 , n5256 );
not ( n6965 , n4232 );
or ( n6966 , n6964 , n6965 );
or ( n6967 , n4232 , n5256 );
nand ( n6968 , n6966 , n6967 );
nand ( n6969 , n6963 , n6968 );
not ( n6970 , n5255 );
not ( n6971 , n4231 );
or ( n6972 , n6970 , n6971 );
or ( n6973 , n4231 , n5255 );
nand ( n6974 , n6972 , n6973 );
not ( n6975 , n5254 );
not ( n6976 , n4230 );
or ( n6977 , n6975 , n6976 );
or ( n6978 , n4230 , n5254 );
nand ( n6979 , n6977 , n6978 );
nand ( n6980 , n6974 , n6979 );
nor ( n6981 , n6969 , n6980 );
nand ( n6982 , n6912 , n6935 , n6958 , n6981 );
not ( n6983 , n5279 );
not ( n6984 , n4255 );
or ( n6985 , n6983 , n6984 );
or ( n6986 , n4255 , n5279 );
nand ( n6987 , n6985 , n6986 );
not ( n6988 , n5278 );
not ( n6989 , n4254 );
or ( n6990 , n6988 , n6989 );
or ( n6991 , n4254 , n5278 );
nand ( n6992 , n6990 , n6991 );
nand ( n6993 , n6987 , n6992 );
not ( n6994 , n5281 );
not ( n6995 , n4257 );
or ( n6996 , n6994 , n6995 );
or ( n6997 , n4257 , n5281 );
nand ( n6998 , n6996 , n6997 );
not ( n6999 , n5280 );
not ( n7000 , n4256 );
or ( n7001 , n6999 , n7000 );
or ( n7002 , n4256 , n5280 );
nand ( n7003 , n7001 , n7002 );
nand ( n7004 , n6998 , n7003 );
nor ( n7005 , n6993 , n7004 );
not ( n7006 , n5283 );
not ( n7007 , n4259 );
or ( n7008 , n7006 , n7007 );
or ( n7009 , n4259 , n5283 );
nand ( n7010 , n7008 , n7009 );
not ( n7011 , n5282 );
not ( n7012 , n4258 );
or ( n7013 , n7011 , n7012 );
or ( n7014 , n4258 , n5282 );
nand ( n7015 , n7013 , n7014 );
nand ( n7016 , n7010 , n7015 );
not ( n7017 , n5285 );
not ( n7018 , n4261 );
or ( n7019 , n7017 , n7018 );
or ( n7020 , n4261 , n5285 );
nand ( n7021 , n7019 , n7020 );
not ( n7022 , n5284 );
not ( n7023 , n4260 );
or ( n7024 , n7022 , n7023 );
or ( n7025 , n4260 , n5284 );
nand ( n7026 , n7024 , n7025 );
nand ( n7027 , n7021 , n7026 );
nor ( n7028 , n7016 , n7027 );
not ( n7029 , n5275 );
not ( n7030 , n4251 );
or ( n7031 , n7029 , n7030 );
or ( n7032 , n4251 , n5275 );
nand ( n7033 , n7031 , n7032 );
not ( n7034 , n5274 );
not ( n7035 , n4250 );
or ( n7036 , n7034 , n7035 );
or ( n7037 , n4250 , n5274 );
nand ( n7038 , n7036 , n7037 );
nand ( n7039 , n7033 , n7038 );
not ( n7040 , n5277 );
not ( n7041 , n4253 );
or ( n7042 , n7040 , n7041 );
or ( n7043 , n4253 , n5277 );
nand ( n7044 , n7042 , n7043 );
not ( n7045 , n5276 );
not ( n7046 , n4252 );
or ( n7047 , n7045 , n7046 );
or ( n7048 , n4252 , n5276 );
nand ( n7049 , n7047 , n7048 );
nand ( n7050 , n7044 , n7049 );
nor ( n7051 , n7039 , n7050 );
not ( n7052 , n5271 );
not ( n7053 , n4247 );
or ( n7054 , n7052 , n7053 );
or ( n7055 , n4247 , n5271 );
nand ( n7056 , n7054 , n7055 );
not ( n7057 , n5270 );
not ( n7058 , n4246 );
or ( n7059 , n7057 , n7058 );
or ( n7060 , n4246 , n5270 );
nand ( n7061 , n7059 , n7060 );
nand ( n7062 , n7056 , n7061 );
not ( n7063 , n5273 );
not ( n7064 , n4249 );
or ( n7065 , n7063 , n7064 );
or ( n7066 , n4249 , n5273 );
nand ( n7067 , n7065 , n7066 );
not ( n7068 , n5272 );
not ( n7069 , n4248 );
or ( n7070 , n7068 , n7069 );
or ( n7071 , n4248 , n5272 );
nand ( n7072 , n7070 , n7071 );
nand ( n7073 , n7067 , n7072 );
nor ( n7074 , n7062 , n7073 );
nand ( n7075 , n7005 , n7028 , n7051 , n7074 );
nor ( n7076 , n6982 , n7075 );
not ( n7077 , n5299 );
not ( n7078 , n4275 );
or ( n7079 , n7077 , n7078 );
or ( n7080 , n4275 , n5299 );
nand ( n7081 , n7079 , n7080 );
not ( n7082 , n5298 );
not ( n7083 , n4274 );
or ( n7084 , n7082 , n7083 );
or ( n7085 , n4274 , n5298 );
nand ( n7086 , n7084 , n7085 );
nand ( n7087 , n7081 , n7086 );
not ( n7088 , n5301 );
not ( n7089 , n4277 );
or ( n7090 , n7088 , n7089 );
or ( n7091 , n4277 , n5301 );
nand ( n7092 , n7090 , n7091 );
not ( n7093 , n5300 );
not ( n7094 , n4276 );
or ( n7095 , n7093 , n7094 );
or ( n7096 , n4276 , n5300 );
nand ( n7097 , n7095 , n7096 );
nand ( n7098 , n7092 , n7097 );
nor ( n7099 , n7087 , n7098 );
not ( n7100 , n5295 );
not ( n7101 , n4271 );
or ( n7102 , n7100 , n7101 );
or ( n7103 , n4271 , n5295 );
nand ( n7104 , n7102 , n7103 );
not ( n7105 , n5294 );
not ( n7106 , n4270 );
or ( n7107 , n7105 , n7106 );
or ( n7108 , n4270 , n5294 );
nand ( n7109 , n7107 , n7108 );
nand ( n7110 , n7104 , n7109 );
not ( n7111 , n5297 );
not ( n7112 , n4273 );
or ( n7113 , n7111 , n7112 );
or ( n7114 , n4273 , n5297 );
nand ( n7115 , n7113 , n7114 );
not ( n7116 , n5296 );
not ( n7117 , n4272 );
or ( n7118 , n7116 , n7117 );
or ( n7119 , n4272 , n5296 );
nand ( n7120 , n7118 , n7119 );
nand ( n7121 , n7115 , n7120 );
nor ( n7122 , n7110 , n7121 );
not ( n7123 , n5291 );
not ( n7124 , n4267 );
or ( n7125 , n7123 , n7124 );
or ( n7126 , n4267 , n5291 );
nand ( n7127 , n7125 , n7126 );
not ( n7128 , n5290 );
not ( n7129 , n4266 );
or ( n7130 , n7128 , n7129 );
or ( n7131 , n4266 , n5290 );
nand ( n7132 , n7130 , n7131 );
nand ( n7133 , n7127 , n7132 );
not ( n7134 , n5293 );
not ( n7135 , n4269 );
or ( n7136 , n7134 , n7135 );
or ( n7137 , n4269 , n5293 );
nand ( n7138 , n7136 , n7137 );
not ( n7139 , n5292 );
not ( n7140 , n4268 );
or ( n7141 , n7139 , n7140 );
or ( n7142 , n4268 , n5292 );
nand ( n7143 , n7141 , n7142 );
nand ( n7144 , n7138 , n7143 );
nor ( n7145 , n7133 , n7144 );
not ( n7146 , n5287 );
not ( n7147 , n4263 );
or ( n7148 , n7146 , n7147 );
or ( n7149 , n4263 , n5287 );
nand ( n7150 , n7148 , n7149 );
not ( n7151 , n5286 );
not ( n7152 , n4262 );
or ( n7153 , n7151 , n7152 );
or ( n7154 , n4262 , n5286 );
nand ( n7155 , n7153 , n7154 );
nand ( n7156 , n7150 , n7155 );
not ( n7157 , n5289 );
not ( n7158 , n4265 );
or ( n7159 , n7157 , n7158 );
or ( n7160 , n4265 , n5289 );
nand ( n7161 , n7159 , n7160 );
not ( n7162 , n5288 );
not ( n7163 , n4264 );
or ( n7164 , n7162 , n7163 );
or ( n7165 , n4264 , n5288 );
nand ( n7166 , n7164 , n7165 );
nand ( n7167 , n7161 , n7166 );
nor ( n7168 , n7156 , n7167 );
nand ( n7169 , n7099 , n7122 , n7145 , n7168 );
not ( n7170 , n5316 );
not ( n7171 , n4292 );
or ( n7172 , n7170 , n7171 );
or ( n7173 , n4292 , n5316 );
nand ( n7174 , n7172 , n7173 );
not ( n7175 , n5317 );
not ( n7176 , n4293 );
or ( n7177 , n7175 , n7176 );
or ( n7178 , n4293 , n5317 );
nand ( n7179 , n7177 , n7178 );
not ( n7180 , n5314 );
not ( n7181 , n4290 );
or ( n7182 , n7180 , n7181 );
or ( n7183 , n4290 , n5314 );
nand ( n7184 , n7182 , n7183 );
not ( n7185 , n5315 );
not ( n7186 , n4291 );
or ( n7187 , n7185 , n7186 );
or ( n7188 , n4291 , n5315 );
nand ( n7189 , n7187 , n7188 );
and ( n7190 , n7174 , n7179 , n7184 , n7189 );
not ( n7191 , n5308 );
not ( n7192 , n4284 );
or ( n7193 , n7191 , n7192 );
or ( n7194 , n4284 , n5308 );
nand ( n7195 , n7193 , n7194 );
not ( n7196 , n5309 );
not ( n7197 , n4285 );
or ( n7198 , n7196 , n7197 );
or ( n7199 , n4285 , n5309 );
nand ( n7200 , n7198 , n7199 );
not ( n7201 , n5306 );
not ( n7202 , n4282 );
or ( n7203 , n7201 , n7202 );
or ( n7204 , n4282 , n5306 );
nand ( n7205 , n7203 , n7204 );
not ( n7206 , n5307 );
not ( n7207 , n4283 );
or ( n7208 , n7206 , n7207 );
or ( n7209 , n4283 , n5307 );
nand ( n7210 , n7208 , n7209 );
and ( n7211 , n7195 , n7200 , n7205 , n7210 );
not ( n7212 , n5312 );
not ( n7213 , n4288 );
or ( n7214 , n7212 , n7213 );
or ( n7215 , n4288 , n5312 );
nand ( n7216 , n7214 , n7215 );
not ( n7217 , n5313 );
not ( n7218 , n4289 );
or ( n7219 , n7217 , n7218 );
or ( n7220 , n4289 , n5313 );
nand ( n7221 , n7219 , n7220 );
not ( n7222 , n5310 );
not ( n7223 , n4286 );
or ( n7224 , n7222 , n7223 );
or ( n7225 , n4286 , n5310 );
nand ( n7226 , n7224 , n7225 );
not ( n7227 , n5311 );
not ( n7228 , n4287 );
or ( n7229 , n7227 , n7228 );
or ( n7230 , n4287 , n5311 );
nand ( n7231 , n7229 , n7230 );
and ( n7232 , n7216 , n7221 , n7226 , n7231 );
not ( n7233 , n4278 );
not ( n7234 , n5302 );
or ( n7235 , n7233 , n7234 );
or ( n7236 , n5302 , n4278 );
nand ( n7237 , n7235 , n7236 );
not ( n7238 , n4279 );
not ( n7239 , n5303 );
or ( n7240 , n7238 , n7239 );
or ( n7241 , n5303 , n4279 );
nand ( n7242 , n7240 , n7241 );
nand ( n7243 , n7237 , n7242 );
not ( n7244 , n4280 );
not ( n7245 , n5304 );
or ( n7246 , n7244 , n7245 );
or ( n7247 , n5304 , n4280 );
nand ( n7248 , n7246 , n7247 );
not ( n7249 , n4281 );
not ( n7250 , n5305 );
or ( n7251 , n7249 , n7250 );
or ( n7252 , n5305 , n4281 );
nand ( n7253 , n7251 , n7252 );
nand ( n7254 , n7248 , n7253 );
nor ( n7255 , n7243 , n7254 );
nand ( n7256 , n7190 , n7211 , n7232 , n7255 );
nor ( n7257 , n7169 , n7256 );
not ( n7258 , n5324 );
not ( n7259 , n4300 );
or ( n7260 , n7258 , n7259 );
or ( n7261 , n4300 , n5324 );
nand ( n7262 , n7260 , n7261 );
not ( n7263 , n5325 );
not ( n7264 , n4301 );
or ( n7265 , n7263 , n7264 );
or ( n7266 , n4301 , n5325 );
nand ( n7267 , n7265 , n7266 );
not ( n7268 , n5322 );
not ( n7269 , n4298 );
or ( n7270 , n7268 , n7269 );
or ( n7271 , n4298 , n5322 );
nand ( n7272 , n7270 , n7271 );
not ( n7273 , n5323 );
not ( n7274 , n4299 );
or ( n7275 , n7273 , n7274 );
or ( n7276 , n4299 , n5323 );
nand ( n7277 , n7275 , n7276 );
nand ( n7278 , n7262 , n7267 , n7272 , n7277 );
not ( n7279 , n5327 );
not ( n7280 , n4303 );
or ( n7281 , n7279 , n7280 );
or ( n7282 , n4303 , n5327 );
nand ( n7283 , n7281 , n7282 );
not ( n7284 , n5329 );
not ( n7285 , n4305 );
or ( n7286 , n7284 , n7285 );
or ( n7287 , n4305 , n5329 );
nand ( n7288 , n7286 , n7287 );
not ( n7289 , n5326 );
not ( n7290 , n4302 );
or ( n7291 , n7289 , n7290 );
or ( n7292 , n4302 , n5326 );
nand ( n7293 , n7291 , n7292 );
not ( n7294 , n5328 );
not ( n7295 , n4304 );
or ( n7296 , n7294 , n7295 );
or ( n7297 , n4304 , n5328 );
nand ( n7298 , n7296 , n7297 );
nand ( n7299 , n7283 , n7288 , n7293 , n7298 );
nor ( n7300 , n7278 , n7299 );
not ( n7301 , n5332 );
not ( n7302 , n4308 );
or ( n7303 , n7301 , n7302 );
or ( n7304 , n4308 , n5332 );
nand ( n7305 , n7303 , n7304 );
not ( n7306 , n5333 );
not ( n7307 , n4309 );
or ( n7308 , n7306 , n7307 );
or ( n7309 , n4309 , n5333 );
nand ( n7310 , n7308 , n7309 );
not ( n7311 , n5330 );
not ( n7312 , n4306 );
or ( n7313 , n7311 , n7312 );
or ( n7314 , n4306 , n5330 );
nand ( n7315 , n7313 , n7314 );
not ( n7316 , n5331 );
not ( n7317 , n4307 );
or ( n7318 , n7316 , n7317 );
or ( n7319 , n4307 , n5331 );
nand ( n7320 , n7318 , n7319 );
nand ( n7321 , n7305 , n7310 , n7315 , n7320 );
not ( n7322 , n4296 );
not ( n7323 , n5320 );
or ( n7324 , n7322 , n7323 );
or ( n7325 , n5320 , n4296 );
nand ( n7326 , n7324 , n7325 );
not ( n7327 , n4297 );
not ( n7328 , n5321 );
or ( n7329 , n7327 , n7328 );
or ( n7330 , n5321 , n4297 );
nand ( n7331 , n7329 , n7330 );
not ( n7332 , n4294 );
not ( n7333 , n5318 );
or ( n7334 , n7332 , n7333 );
or ( n7335 , n5318 , n4294 );
nand ( n7336 , n7334 , n7335 );
not ( n7337 , n4295 );
not ( n7338 , n5319 );
or ( n7339 , n7337 , n7338 );
or ( n7340 , n5319 , n4295 );
nand ( n7341 , n7339 , n7340 );
nand ( n7342 , n7326 , n7331 , n7336 , n7341 );
nor ( n7343 , n7321 , n7342 );
nand ( n7344 , n7300 , n7343 );
not ( n7345 , n5347 );
not ( n7346 , n4323 );
or ( n7347 , n7345 , n7346 );
or ( n7348 , n4323 , n5347 );
nand ( n7349 , n7347 , n7348 );
not ( n7350 , n5346 );
not ( n7351 , n4322 );
or ( n7352 , n7350 , n7351 );
or ( n7353 , n4322 , n5346 );
nand ( n7354 , n7352 , n7353 );
nand ( n7355 , n7349 , n7354 );
not ( n7356 , n5349 );
not ( n7357 , n4325 );
or ( n7358 , n7356 , n7357 );
or ( n7359 , n4325 , n5349 );
nand ( n7360 , n7358 , n7359 );
not ( n7361 , n5348 );
not ( n7362 , n4324 );
or ( n7363 , n7361 , n7362 );
or ( n7364 , n4324 , n5348 );
nand ( n7365 , n7363 , n7364 );
nand ( n7366 , n7360 , n7365 );
nor ( n7367 , n7355 , n7366 );
not ( n7368 , n5343 );
not ( n7369 , n4319 );
or ( n7370 , n7368 , n7369 );
or ( n7371 , n4319 , n5343 );
nand ( n7372 , n7370 , n7371 );
not ( n7373 , n5342 );
not ( n7374 , n4318 );
or ( n7375 , n7373 , n7374 );
or ( n7376 , n4318 , n5342 );
nand ( n7377 , n7375 , n7376 );
nand ( n7378 , n7372 , n7377 );
not ( n7379 , n5345 );
not ( n7380 , n4321 );
or ( n7381 , n7379 , n7380 );
or ( n7382 , n4321 , n5345 );
nand ( n7383 , n7381 , n7382 );
not ( n7384 , n5344 );
not ( n7385 , n4320 );
or ( n7386 , n7384 , n7385 );
or ( n7387 , n4320 , n5344 );
nand ( n7388 , n7386 , n7387 );
nand ( n7389 , n7383 , n7388 );
nor ( n7390 , n7378 , n7389 );
not ( n7391 , n5339 );
not ( n7392 , n4315 );
or ( n7393 , n7391 , n7392 );
or ( n7394 , n4315 , n5339 );
nand ( n7395 , n7393 , n7394 );
not ( n7396 , n5338 );
not ( n7397 , n4314 );
or ( n7398 , n7396 , n7397 );
or ( n7399 , n4314 , n5338 );
nand ( n7400 , n7398 , n7399 );
nand ( n7401 , n7395 , n7400 );
not ( n7402 , n5341 );
not ( n7403 , n4317 );
or ( n7404 , n7402 , n7403 );
or ( n7405 , n4317 , n5341 );
nand ( n7406 , n7404 , n7405 );
not ( n7407 , n5340 );
not ( n7408 , n4316 );
or ( n7409 , n7407 , n7408 );
or ( n7410 , n4316 , n5340 );
nand ( n7411 , n7409 , n7410 );
nand ( n7412 , n7406 , n7411 );
nor ( n7413 , n7401 , n7412 );
not ( n7414 , n5335 );
not ( n7415 , n4311 );
or ( n7416 , n7414 , n7415 );
or ( n7417 , n4311 , n5335 );
nand ( n7418 , n7416 , n7417 );
not ( n7419 , n5334 );
not ( n7420 , n4310 );
or ( n7421 , n7419 , n7420 );
or ( n7422 , n4310 , n5334 );
nand ( n7423 , n7421 , n7422 );
nand ( n7424 , n7418 , n7423 );
not ( n7425 , n5337 );
not ( n7426 , n4313 );
or ( n7427 , n7425 , n7426 );
or ( n7428 , n4313 , n5337 );
nand ( n7429 , n7427 , n7428 );
not ( n7430 , n5336 );
not ( n7431 , n4312 );
or ( n7432 , n7430 , n7431 );
or ( n7433 , n4312 , n5336 );
nand ( n7434 , n7432 , n7433 );
nand ( n7435 , n7429 , n7434 );
nor ( n7436 , n7424 , n7435 );
nand ( n7437 , n7367 , n7390 , n7413 , n7436 );
nor ( n7438 , n7344 , n7437 );
not ( n7439 , n5358 );
not ( n7440 , n4334 );
or ( n7441 , n7439 , n7440 );
or ( n7442 , n4334 , n5358 );
nand ( n7443 , n7441 , n7442 );
not ( n7444 , n5359 );
not ( n7445 , n4335 );
or ( n7446 , n7444 , n7445 );
or ( n7447 , n4335 , n5359 );
nand ( n7448 , n7446 , n7447 );
not ( n7449 , n5360 );
not ( n7450 , n4336 );
or ( n7451 , n7449 , n7450 );
or ( n7452 , n4336 , n5360 );
nand ( n7453 , n7451 , n7452 );
not ( n7454 , n5361 );
not ( n7455 , n4337 );
or ( n7456 , n7454 , n7455 );
or ( n7457 , n4337 , n5361 );
nand ( n7458 , n7456 , n7457 );
nand ( n7459 , n7443 , n7448 , n7453 , n7458 );
not ( n7460 , n5364 );
not ( n7461 , n4340 );
or ( n7462 , n7460 , n7461 );
or ( n7463 , n4340 , n5364 );
nand ( n7464 , n7462 , n7463 );
not ( n7465 , n5365 );
not ( n7466 , n4341 );
or ( n7467 , n7465 , n7466 );
or ( n7468 , n4341 , n5365 );
nand ( n7469 , n7467 , n7468 );
not ( n7470 , n5362 );
not ( n7471 , n4338 );
or ( n7472 , n7470 , n7471 );
or ( n7473 , n4338 , n5362 );
nand ( n7474 , n7472 , n7473 );
not ( n7475 , n5363 );
not ( n7476 , n4339 );
or ( n7477 , n7475 , n7476 );
or ( n7478 , n4339 , n5363 );
nand ( n7479 , n7477 , n7478 );
nand ( n7480 , n7464 , n7469 , n7474 , n7479 );
nor ( n7481 , n7459 , n7480 );
not ( n7482 , n5356 );
not ( n7483 , n4332 );
or ( n7484 , n7482 , n7483 );
or ( n7485 , n4332 , n5356 );
nand ( n7486 , n7484 , n7485 );
not ( n7487 , n5357 );
not ( n7488 , n4333 );
or ( n7489 , n7487 , n7488 );
or ( n7490 , n4333 , n5357 );
nand ( n7491 , n7489 , n7490 );
not ( n7492 , n5354 );
not ( n7493 , n4330 );
or ( n7494 , n7492 , n7493 );
or ( n7495 , n4330 , n5354 );
nand ( n7496 , n7494 , n7495 );
not ( n7497 , n5355 );
not ( n7498 , n4331 );
or ( n7499 , n7497 , n7498 );
or ( n7500 , n4331 , n5355 );
nand ( n7501 , n7499 , n7500 );
nand ( n7502 , n7486 , n7491 , n7496 , n7501 );
not ( n7503 , n5352 );
not ( n7504 , n4328 );
or ( n7505 , n7503 , n7504 );
or ( n7506 , n4328 , n5352 );
nand ( n7507 , n7505 , n7506 );
not ( n7508 , n5353 );
not ( n7509 , n4329 );
or ( n7510 , n7508 , n7509 );
or ( n7511 , n4329 , n5353 );
nand ( n7512 , n7510 , n7511 );
not ( n7513 , n5350 );
not ( n7514 , n4326 );
or ( n7515 , n7513 , n7514 );
or ( n7516 , n4326 , n5350 );
nand ( n7517 , n7515 , n7516 );
not ( n7518 , n5351 );
not ( n7519 , n4327 );
or ( n7520 , n7518 , n7519 );
or ( n7521 , n4327 , n5351 );
nand ( n7522 , n7520 , n7521 );
nand ( n7523 , n7507 , n7512 , n7517 , n7522 );
nor ( n7524 , n7502 , n7523 );
nand ( n7525 , n7481 , n7524 );
not ( n7526 , n5379 );
not ( n7527 , n4355 );
or ( n7528 , n7526 , n7527 );
or ( n7529 , n4355 , n5379 );
nand ( n7530 , n7528 , n7529 );
not ( n7531 , n5378 );
not ( n7532 , n4354 );
or ( n7533 , n7531 , n7532 );
or ( n7534 , n4354 , n5378 );
nand ( n7535 , n7533 , n7534 );
nand ( n7536 , n7530 , n7535 );
not ( n7537 , n5381 );
not ( n7538 , n4357 );
or ( n7539 , n7537 , n7538 );
or ( n7540 , n4357 , n5381 );
nand ( n7541 , n7539 , n7540 );
not ( n7542 , n5380 );
not ( n7543 , n4356 );
or ( n7544 , n7542 , n7543 );
or ( n7545 , n4356 , n5380 );
nand ( n7546 , n7544 , n7545 );
nand ( n7547 , n7541 , n7546 );
nor ( n7548 , n7536 , n7547 );
not ( n7549 , n5375 );
not ( n7550 , n4351 );
or ( n7551 , n7549 , n7550 );
or ( n7552 , n4351 , n5375 );
nand ( n7553 , n7551 , n7552 );
not ( n7554 , n5374 );
not ( n7555 , n4350 );
or ( n7556 , n7554 , n7555 );
or ( n7557 , n4350 , n5374 );
nand ( n7558 , n7556 , n7557 );
nand ( n7559 , n7553 , n7558 );
not ( n7560 , n5377 );
not ( n7561 , n4353 );
or ( n7562 , n7560 , n7561 );
or ( n7563 , n4353 , n5377 );
nand ( n7564 , n7562 , n7563 );
not ( n7565 , n5376 );
not ( n7566 , n4352 );
or ( n7567 , n7565 , n7566 );
or ( n7568 , n4352 , n5376 );
nand ( n7569 , n7567 , n7568 );
nand ( n7570 , n7564 , n7569 );
nor ( n7571 , n7559 , n7570 );
not ( n7572 , n5367 );
not ( n7573 , n4343 );
or ( n7574 , n7572 , n7573 );
or ( n7575 , n4343 , n5367 );
nand ( n7576 , n7574 , n7575 );
not ( n7577 , n5366 );
not ( n7578 , n4342 );
or ( n7579 , n7577 , n7578 );
or ( n7580 , n4342 , n5366 );
nand ( n7581 , n7579 , n7580 );
nand ( n7582 , n7576 , n7581 );
not ( n7583 , n5369 );
not ( n7584 , n4345 );
or ( n7585 , n7583 , n7584 );
or ( n7586 , n4345 , n5369 );
nand ( n7587 , n7585 , n7586 );
not ( n7588 , n5368 );
not ( n7589 , n4344 );
or ( n7590 , n7588 , n7589 );
or ( n7591 , n4344 , n5368 );
nand ( n7592 , n7590 , n7591 );
nand ( n7593 , n7587 , n7592 );
nor ( n7594 , n7582 , n7593 );
not ( n7595 , n5373 );
not ( n7596 , n4349 );
or ( n7597 , n7595 , n7596 );
or ( n7598 , n4349 , n5373 );
nand ( n7599 , n7597 , n7598 );
not ( n7600 , n5372 );
not ( n7601 , n4348 );
or ( n7602 , n7600 , n7601 );
or ( n7603 , n4348 , n5372 );
nand ( n7604 , n7602 , n7603 );
nand ( n7605 , n7599 , n7604 );
not ( n7606 , n5371 );
not ( n7607 , n4347 );
or ( n7608 , n7606 , n7607 );
or ( n7609 , n4347 , n5371 );
nand ( n7610 , n7608 , n7609 );
not ( n7611 , n5370 );
not ( n7612 , n4346 );
or ( n7613 , n7611 , n7612 );
or ( n7614 , n4346 , n5370 );
nand ( n7615 , n7613 , n7614 );
nand ( n7616 , n7610 , n7615 );
nor ( n7617 , n7605 , n7616 );
nand ( n7618 , n7548 , n7571 , n7594 , n7617 );
nor ( n7619 , n7525 , n7618 );
nand ( n7620 , n7076 , n7257 , n7438 , n7619 );
nor ( n7621 , n6889 , n7620 );
not ( n7622 , n5391 );
not ( n7623 , n4367 );
or ( n7624 , n7622 , n7623 );
or ( n7625 , n4367 , n5391 );
nand ( n7626 , n7624 , n7625 );
not ( n7627 , n5390 );
not ( n7628 , n4366 );
or ( n7629 , n7627 , n7628 );
or ( n7630 , n4366 , n5390 );
nand ( n7631 , n7629 , n7630 );
nand ( n7632 , n7626 , n7631 );
not ( n7633 , n5393 );
not ( n7634 , n4369 );
or ( n7635 , n7633 , n7634 );
or ( n7636 , n4369 , n5393 );
nand ( n7637 , n7635 , n7636 );
not ( n7638 , n5392 );
not ( n7639 , n4368 );
or ( n7640 , n7638 , n7639 );
or ( n7641 , n4368 , n5392 );
nand ( n7642 , n7640 , n7641 );
nand ( n7643 , n7637 , n7642 );
nor ( n7644 , n7632 , n7643 );
not ( n7645 , n5387 );
not ( n7646 , n4363 );
or ( n7647 , n7645 , n7646 );
or ( n7648 , n4363 , n5387 );
nand ( n7649 , n7647 , n7648 );
not ( n7650 , n5386 );
not ( n7651 , n4362 );
or ( n7652 , n7650 , n7651 );
or ( n7653 , n4362 , n5386 );
nand ( n7654 , n7652 , n7653 );
nand ( n7655 , n7649 , n7654 );
not ( n7656 , n5389 );
not ( n7657 , n4365 );
or ( n7658 , n7656 , n7657 );
or ( n7659 , n4365 , n5389 );
nand ( n7660 , n7658 , n7659 );
not ( n7661 , n5388 );
not ( n7662 , n4364 );
or ( n7663 , n7661 , n7662 );
or ( n7664 , n4364 , n5388 );
nand ( n7665 , n7663 , n7664 );
nand ( n7666 , n7660 , n7665 );
nor ( n7667 , n7655 , n7666 );
not ( n7668 , n5385 );
not ( n7669 , n4361 );
or ( n7670 , n7668 , n7669 );
or ( n7671 , n4361 , n5385 );
nand ( n7672 , n7670 , n7671 );
not ( n7673 , n5384 );
not ( n7674 , n4360 );
or ( n7675 , n7673 , n7674 );
or ( n7676 , n4360 , n5384 );
nand ( n7677 , n7675 , n7676 );
nand ( n7678 , n7672 , n7677 );
not ( n7679 , n5383 );
not ( n7680 , n4359 );
or ( n7681 , n7679 , n7680 );
or ( n7682 , n4359 , n5383 );
nand ( n7683 , n7681 , n7682 );
not ( n7684 , n5382 );
not ( n7685 , n4358 );
or ( n7686 , n7684 , n7685 );
or ( n7687 , n4358 , n5382 );
nand ( n7688 , n7686 , n7687 );
nand ( n7689 , n7683 , n7688 );
nor ( n7690 , n7678 , n7689 );
not ( n7691 , n5396 );
not ( n7692 , n4372 );
or ( n7693 , n7691 , n7692 );
or ( n7694 , n4372 , n5396 );
nand ( n7695 , n7693 , n7694 );
not ( n7696 , n5397 );
not ( n7697 , n4373 );
or ( n7698 , n7696 , n7697 );
or ( n7699 , n4373 , n5397 );
nand ( n7700 , n7698 , n7699 );
not ( n7701 , n5394 );
not ( n7702 , n4370 );
or ( n7703 , n7701 , n7702 );
or ( n7704 , n4370 , n5394 );
nand ( n7705 , n7703 , n7704 );
not ( n7706 , n5395 );
not ( n7707 , n4371 );
or ( n7708 , n7706 , n7707 );
or ( n7709 , n4371 , n5395 );
nand ( n7710 , n7708 , n7709 );
and ( n7711 , n7695 , n7700 , n7705 , n7710 );
nand ( n7712 , n7644 , n7667 , n7690 , n7711 );
not ( n7713 , n5411 );
not ( n7714 , n4387 );
or ( n7715 , n7713 , n7714 );
or ( n7716 , n4387 , n5411 );
nand ( n7717 , n7715 , n7716 );
not ( n7718 , n5410 );
not ( n7719 , n4386 );
or ( n7720 , n7718 , n7719 );
or ( n7721 , n4386 , n5410 );
nand ( n7722 , n7720 , n7721 );
nand ( n7723 , n7717 , n7722 );
not ( n7724 , n5413 );
not ( n7725 , n4389 );
or ( n7726 , n7724 , n7725 );
or ( n7727 , n4389 , n5413 );
nand ( n7728 , n7726 , n7727 );
not ( n7729 , n5412 );
not ( n7730 , n4388 );
or ( n7731 , n7729 , n7730 );
or ( n7732 , n4388 , n5412 );
nand ( n7733 , n7731 , n7732 );
nand ( n7734 , n7728 , n7733 );
nor ( n7735 , n7723 , n7734 );
not ( n7736 , n5407 );
not ( n7737 , n4383 );
or ( n7738 , n7736 , n7737 );
or ( n7739 , n4383 , n5407 );
nand ( n7740 , n7738 , n7739 );
not ( n7741 , n5406 );
not ( n7742 , n4382 );
or ( n7743 , n7741 , n7742 );
or ( n7744 , n4382 , n5406 );
nand ( n7745 , n7743 , n7744 );
nand ( n7746 , n7740 , n7745 );
not ( n7747 , n5409 );
not ( n7748 , n4385 );
or ( n7749 , n7747 , n7748 );
or ( n7750 , n4385 , n5409 );
nand ( n7751 , n7749 , n7750 );
not ( n7752 , n5408 );
not ( n7753 , n4384 );
or ( n7754 , n7752 , n7753 );
or ( n7755 , n4384 , n5408 );
nand ( n7756 , n7754 , n7755 );
nand ( n7757 , n7751 , n7756 );
nor ( n7758 , n7746 , n7757 );
not ( n7759 , n5403 );
not ( n7760 , n4379 );
or ( n7761 , n7759 , n7760 );
or ( n7762 , n4379 , n5403 );
nand ( n7763 , n7761 , n7762 );
not ( n7764 , n5402 );
not ( n7765 , n4378 );
or ( n7766 , n7764 , n7765 );
or ( n7767 , n4378 , n5402 );
nand ( n7768 , n7766 , n7767 );
nand ( n7769 , n7763 , n7768 );
not ( n7770 , n5405 );
not ( n7771 , n4381 );
or ( n7772 , n7770 , n7771 );
or ( n7773 , n4381 , n5405 );
nand ( n7774 , n7772 , n7773 );
not ( n7775 , n5404 );
not ( n7776 , n4380 );
or ( n7777 , n7775 , n7776 );
or ( n7778 , n4380 , n5404 );
nand ( n7779 , n7777 , n7778 );
nand ( n7780 , n7774 , n7779 );
nor ( n7781 , n7769 , n7780 );
not ( n7782 , n5399 );
not ( n7783 , n4375 );
or ( n7784 , n7782 , n7783 );
or ( n7785 , n4375 , n5399 );
nand ( n7786 , n7784 , n7785 );
not ( n7787 , n5398 );
not ( n7788 , n4374 );
or ( n7789 , n7787 , n7788 );
or ( n7790 , n4374 , n5398 );
nand ( n7791 , n7789 , n7790 );
nand ( n7792 , n7786 , n7791 );
not ( n7793 , n5401 );
not ( n7794 , n4377 );
or ( n7795 , n7793 , n7794 );
or ( n7796 , n4377 , n5401 );
nand ( n7797 , n7795 , n7796 );
not ( n7798 , n5400 );
not ( n7799 , n4376 );
or ( n7800 , n7798 , n7799 );
or ( n7801 , n4376 , n5400 );
nand ( n7802 , n7800 , n7801 );
nand ( n7803 , n7797 , n7802 );
nor ( n7804 , n7792 , n7803 );
nand ( n7805 , n7735 , n7758 , n7781 , n7804 );
nor ( n7806 , n7712 , n7805 );
not ( n7807 , n5419 );
not ( n7808 , n4395 );
or ( n7809 , n7807 , n7808 );
or ( n7810 , n4395 , n5419 );
nand ( n7811 , n7809 , n7810 );
not ( n7812 , n5418 );
not ( n7813 , n4394 );
or ( n7814 , n7812 , n7813 );
or ( n7815 , n4394 , n5418 );
nand ( n7816 , n7814 , n7815 );
nand ( n7817 , n7811 , n7816 );
not ( n7818 , n5421 );
not ( n7819 , n4397 );
or ( n7820 , n7818 , n7819 );
or ( n7821 , n4397 , n5421 );
nand ( n7822 , n7820 , n7821 );
not ( n7823 , n5420 );
not ( n7824 , n4396 );
or ( n7825 , n7823 , n7824 );
or ( n7826 , n4396 , n5420 );
nand ( n7827 , n7825 , n7826 );
nand ( n7828 , n7822 , n7827 );
nor ( n7829 , n7817 , n7828 );
not ( n7830 , n5427 );
not ( n7831 , n4403 );
or ( n7832 , n7830 , n7831 );
or ( n7833 , n4403 , n5427 );
nand ( n7834 , n7832 , n7833 );
not ( n7835 , n5426 );
not ( n7836 , n4402 );
or ( n7837 , n7835 , n7836 );
or ( n7838 , n4402 , n5426 );
nand ( n7839 , n7837 , n7838 );
nand ( n7840 , n7834 , n7839 );
not ( n7841 , n5429 );
not ( n7842 , n4405 );
or ( n7843 , n7841 , n7842 );
or ( n7844 , n4405 , n5429 );
nand ( n7845 , n7843 , n7844 );
not ( n7846 , n5428 );
not ( n7847 , n4404 );
or ( n7848 , n7846 , n7847 );
or ( n7849 , n4404 , n5428 );
nand ( n7850 , n7848 , n7849 );
nand ( n7851 , n7845 , n7850 );
nor ( n7852 , n7840 , n7851 );
not ( n7853 , n5415 );
not ( n7854 , n4391 );
or ( n7855 , n7853 , n7854 );
or ( n7856 , n4391 , n5415 );
nand ( n7857 , n7855 , n7856 );
not ( n7858 , n5414 );
not ( n7859 , n4390 );
or ( n7860 , n7858 , n7859 );
or ( n7861 , n4390 , n5414 );
nand ( n7862 , n7860 , n7861 );
nand ( n7863 , n7857 , n7862 );
not ( n7864 , n5417 );
not ( n7865 , n4393 );
or ( n7866 , n7864 , n7865 );
or ( n7867 , n4393 , n5417 );
nand ( n7868 , n7866 , n7867 );
not ( n7869 , n5416 );
not ( n7870 , n4392 );
or ( n7871 , n7869 , n7870 );
or ( n7872 , n4392 , n5416 );
nand ( n7873 , n7871 , n7872 );
nand ( n7874 , n7868 , n7873 );
nor ( n7875 , n7863 , n7874 );
not ( n7876 , n5423 );
not ( n7877 , n4399 );
or ( n7878 , n7876 , n7877 );
or ( n7879 , n4399 , n5423 );
nand ( n7880 , n7878 , n7879 );
not ( n7881 , n5425 );
not ( n7882 , n4401 );
or ( n7883 , n7881 , n7882 );
or ( n7884 , n4401 , n5425 );
nand ( n7885 , n7883 , n7884 );
not ( n7886 , n5422 );
not ( n7887 , n4398 );
or ( n7888 , n7886 , n7887 );
or ( n7889 , n4398 , n5422 );
nand ( n7890 , n7888 , n7889 );
not ( n7891 , n5424 );
not ( n7892 , n4400 );
or ( n7893 , n7891 , n7892 );
or ( n7894 , n4400 , n5424 );
nand ( n7895 , n7893 , n7894 );
and ( n7896 , n7880 , n7885 , n7890 , n7895 );
nand ( n7897 , n7829 , n7852 , n7875 , n7896 );
not ( n7898 , n5443 );
not ( n7899 , n4419 );
or ( n7900 , n7898 , n7899 );
or ( n7901 , n4419 , n5443 );
nand ( n7902 , n7900 , n7901 );
not ( n7903 , n5442 );
not ( n7904 , n4418 );
or ( n7905 , n7903 , n7904 );
or ( n7906 , n4418 , n5442 );
nand ( n7907 , n7905 , n7906 );
nand ( n7908 , n7902 , n7907 );
not ( n7909 , n5445 );
not ( n7910 , n4421 );
or ( n7911 , n7909 , n7910 );
or ( n7912 , n4421 , n5445 );
nand ( n7913 , n7911 , n7912 );
not ( n7914 , n5444 );
not ( n7915 , n4420 );
or ( n7916 , n7914 , n7915 );
or ( n7917 , n4420 , n5444 );
nand ( n7918 , n7916 , n7917 );
nand ( n7919 , n7913 , n7918 );
nor ( n7920 , n7908 , n7919 );
not ( n7921 , n5439 );
not ( n7922 , n4415 );
or ( n7923 , n7921 , n7922 );
or ( n7924 , n4415 , n5439 );
nand ( n7925 , n7923 , n7924 );
not ( n7926 , n5438 );
not ( n7927 , n4414 );
or ( n7928 , n7926 , n7927 );
or ( n7929 , n4414 , n5438 );
nand ( n7930 , n7928 , n7929 );
nand ( n7931 , n7925 , n7930 );
not ( n7932 , n5441 );
not ( n7933 , n4417 );
or ( n7934 , n7932 , n7933 );
or ( n7935 , n4417 , n5441 );
nand ( n7936 , n7934 , n7935 );
not ( n7937 , n5440 );
not ( n7938 , n4416 );
or ( n7939 , n7937 , n7938 );
or ( n7940 , n4416 , n5440 );
nand ( n7941 , n7939 , n7940 );
nand ( n7942 , n7936 , n7941 );
nor ( n7943 , n7931 , n7942 );
not ( n7944 , n5435 );
not ( n7945 , n4411 );
or ( n7946 , n7944 , n7945 );
or ( n7947 , n4411 , n5435 );
nand ( n7948 , n7946 , n7947 );
not ( n7949 , n5434 );
not ( n7950 , n4410 );
or ( n7951 , n7949 , n7950 );
or ( n7952 , n4410 , n5434 );
nand ( n7953 , n7951 , n7952 );
nand ( n7954 , n7948 , n7953 );
not ( n7955 , n5437 );
not ( n7956 , n4413 );
or ( n7957 , n7955 , n7956 );
or ( n7958 , n4413 , n5437 );
nand ( n7959 , n7957 , n7958 );
not ( n7960 , n5436 );
not ( n7961 , n4412 );
or ( n7962 , n7960 , n7961 );
or ( n7963 , n4412 , n5436 );
nand ( n7964 , n7962 , n7963 );
nand ( n7965 , n7959 , n7964 );
nor ( n7966 , n7954 , n7965 );
not ( n7967 , n5431 );
not ( n7968 , n4407 );
or ( n7969 , n7967 , n7968 );
or ( n7970 , n4407 , n5431 );
nand ( n7971 , n7969 , n7970 );
not ( n7972 , n5430 );
not ( n7973 , n4406 );
or ( n7974 , n7972 , n7973 );
or ( n7975 , n4406 , n5430 );
nand ( n7976 , n7974 , n7975 );
nand ( n7977 , n7971 , n7976 );
not ( n7978 , n5433 );
not ( n7979 , n4409 );
or ( n7980 , n7978 , n7979 );
or ( n7981 , n4409 , n5433 );
nand ( n7982 , n7980 , n7981 );
not ( n7983 , n5432 );
not ( n7984 , n4408 );
or ( n7985 , n7983 , n7984 );
or ( n7986 , n4408 , n5432 );
nand ( n7987 , n7985 , n7986 );
nand ( n7988 , n7982 , n7987 );
nor ( n7989 , n7977 , n7988 );
nand ( n7990 , n7920 , n7943 , n7966 , n7989 );
nor ( n7991 , n7897 , n7990 );
not ( n7992 , n5507 );
not ( n7993 , n4483 );
or ( n7994 , n7992 , n7993 );
or ( n7995 , n4483 , n5507 );
nand ( n7996 , n7994 , n7995 );
not ( n7997 , n5506 );
not ( n7998 , n4482 );
or ( n7999 , n7997 , n7998 );
or ( n8000 , n4482 , n5506 );
nand ( n8001 , n7999 , n8000 );
nand ( n8002 , n7996 , n8001 );
not ( n8003 , n5509 );
not ( n8004 , n4485 );
or ( n8005 , n8003 , n8004 );
or ( n8006 , n4485 , n5509 );
nand ( n8007 , n8005 , n8006 );
not ( n8008 , n5508 );
not ( n8009 , n4484 );
or ( n8010 , n8008 , n8009 );
or ( n8011 , n4484 , n5508 );
nand ( n8012 , n8010 , n8011 );
nand ( n8013 , n8007 , n8012 );
nor ( n8014 , n8002 , n8013 );
not ( n8015 , n5503 );
not ( n8016 , n4479 );
or ( n8017 , n8015 , n8016 );
or ( n8018 , n4479 , n5503 );
nand ( n8019 , n8017 , n8018 );
not ( n8020 , n5502 );
not ( n8021 , n4478 );
or ( n8022 , n8020 , n8021 );
or ( n8023 , n4478 , n5502 );
nand ( n8024 , n8022 , n8023 );
nand ( n8025 , n8019 , n8024 );
not ( n8026 , n5505 );
not ( n8027 , n4481 );
or ( n8028 , n8026 , n8027 );
or ( n8029 , n4481 , n5505 );
nand ( n8030 , n8028 , n8029 );
not ( n8031 , n5504 );
not ( n8032 , n4480 );
or ( n8033 , n8031 , n8032 );
or ( n8034 , n4480 , n5504 );
nand ( n8035 , n8033 , n8034 );
nand ( n8036 , n8030 , n8035 );
nor ( n8037 , n8025 , n8036 );
not ( n8038 , n5499 );
not ( n8039 , n4475 );
or ( n8040 , n8038 , n8039 );
or ( n8041 , n4475 , n5499 );
nand ( n8042 , n8040 , n8041 );
not ( n8043 , n5498 );
not ( n8044 , n4474 );
or ( n8045 , n8043 , n8044 );
or ( n8046 , n4474 , n5498 );
nand ( n8047 , n8045 , n8046 );
nand ( n8048 , n8042 , n8047 );
not ( n8049 , n5501 );
not ( n8050 , n4477 );
or ( n8051 , n8049 , n8050 );
or ( n8052 , n4477 , n5501 );
nand ( n8053 , n8051 , n8052 );
not ( n8054 , n5500 );
not ( n8055 , n4476 );
or ( n8056 , n8054 , n8055 );
or ( n8057 , n4476 , n5500 );
nand ( n8058 , n8056 , n8057 );
nand ( n8059 , n8053 , n8058 );
nor ( n8060 , n8048 , n8059 );
not ( n8061 , n5495 );
not ( n8062 , n4471 );
or ( n8063 , n8061 , n8062 );
or ( n8064 , n4471 , n5495 );
nand ( n8065 , n8063 , n8064 );
not ( n8066 , n5494 );
not ( n8067 , n4470 );
or ( n8068 , n8066 , n8067 );
or ( n8069 , n4470 , n5494 );
nand ( n8070 , n8068 , n8069 );
nand ( n8071 , n8065 , n8070 );
not ( n8072 , n5497 );
not ( n8073 , n4473 );
or ( n8074 , n8072 , n8073 );
or ( n8075 , n4473 , n5497 );
nand ( n8076 , n8074 , n8075 );
not ( n8077 , n5496 );
not ( n8078 , n4472 );
or ( n8079 , n8077 , n8078 );
or ( n8080 , n4472 , n5496 );
nand ( n8081 , n8079 , n8080 );
nand ( n8082 , n8076 , n8081 );
nor ( n8083 , n8071 , n8082 );
nand ( n8084 , n8014 , n8037 , n8060 , n8083 );
not ( n8085 , n5491 );
not ( n8086 , n4467 );
or ( n8087 , n8085 , n8086 );
or ( n8088 , n4467 , n5491 );
nand ( n8089 , n8087 , n8088 );
not ( n8090 , n5490 );
not ( n8091 , n4466 );
or ( n8092 , n8090 , n8091 );
or ( n8093 , n4466 , n5490 );
nand ( n8094 , n8092 , n8093 );
nand ( n8095 , n8089 , n8094 );
not ( n8096 , n5493 );
not ( n8097 , n4469 );
or ( n8098 , n8096 , n8097 );
or ( n8099 , n4469 , n5493 );
nand ( n8100 , n8098 , n8099 );
not ( n8101 , n5492 );
not ( n8102 , n4468 );
or ( n8103 , n8101 , n8102 );
or ( n8104 , n4468 , n5492 );
nand ( n8105 , n8103 , n8104 );
nand ( n8106 , n8100 , n8105 );
nor ( n8107 , n8095 , n8106 );
not ( n8108 , n5487 );
not ( n8109 , n4463 );
or ( n8110 , n8108 , n8109 );
or ( n8111 , n4463 , n5487 );
nand ( n8112 , n8110 , n8111 );
not ( n8113 , n5486 );
not ( n8114 , n4462 );
or ( n8115 , n8113 , n8114 );
or ( n8116 , n4462 , n5486 );
nand ( n8117 , n8115 , n8116 );
nand ( n8118 , n8112 , n8117 );
not ( n8119 , n5489 );
not ( n8120 , n4465 );
or ( n8121 , n8119 , n8120 );
or ( n8122 , n4465 , n5489 );
nand ( n8123 , n8121 , n8122 );
not ( n8124 , n5488 );
not ( n8125 , n4464 );
or ( n8126 , n8124 , n8125 );
or ( n8127 , n4464 , n5488 );
nand ( n8128 , n8126 , n8127 );
nand ( n8129 , n8123 , n8128 );
nor ( n8130 , n8118 , n8129 );
not ( n8131 , n5483 );
not ( n8132 , n4459 );
or ( n8133 , n8131 , n8132 );
or ( n8134 , n4459 , n5483 );
nand ( n8135 , n8133 , n8134 );
not ( n8136 , n5482 );
not ( n8137 , n4458 );
or ( n8138 , n8136 , n8137 );
or ( n8139 , n4458 , n5482 );
nand ( n8140 , n8138 , n8139 );
nand ( n8141 , n8135 , n8140 );
not ( n8142 , n5485 );
not ( n8143 , n4461 );
or ( n8144 , n8142 , n8143 );
or ( n8145 , n4461 , n5485 );
nand ( n8146 , n8144 , n8145 );
not ( n8147 , n5484 );
not ( n8148 , n4460 );
or ( n8149 , n8147 , n8148 );
or ( n8150 , n4460 , n5484 );
nand ( n8151 , n8149 , n8150 );
nand ( n8152 , n8146 , n8151 );
nor ( n8153 , n8141 , n8152 );
not ( n8154 , n5479 );
not ( n8155 , n4455 );
or ( n8156 , n8154 , n8155 );
or ( n8157 , n4455 , n5479 );
nand ( n8158 , n8156 , n8157 );
not ( n8159 , n5478 );
not ( n8160 , n4454 );
or ( n8161 , n8159 , n8160 );
or ( n8162 , n4454 , n5478 );
nand ( n8163 , n8161 , n8162 );
nand ( n8164 , n8158 , n8163 );
not ( n8165 , n5481 );
not ( n8166 , n4457 );
or ( n8167 , n8165 , n8166 );
or ( n8168 , n4457 , n5481 );
nand ( n8169 , n8167 , n8168 );
not ( n8170 , n5480 );
not ( n8171 , n4456 );
or ( n8172 , n8170 , n8171 );
or ( n8173 , n4456 , n5480 );
nand ( n8174 , n8172 , n8173 );
nand ( n8175 , n8169 , n8174 );
nor ( n8176 , n8164 , n8175 );
nand ( n8177 , n8107 , n8130 , n8153 , n8176 );
nor ( n8178 , n8084 , n8177 );
not ( n8179 , n5451 );
not ( n8180 , n4427 );
or ( n8181 , n8179 , n8180 );
or ( n8182 , n4427 , n5451 );
nand ( n8183 , n8181 , n8182 );
not ( n8184 , n5450 );
not ( n8185 , n4426 );
or ( n8186 , n8184 , n8185 );
or ( n8187 , n4426 , n5450 );
nand ( n8188 , n8186 , n8187 );
nand ( n8189 , n8183 , n8188 );
not ( n8190 , n5453 );
not ( n8191 , n4429 );
or ( n8192 , n8190 , n8191 );
or ( n8193 , n4429 , n5453 );
nand ( n8194 , n8192 , n8193 );
not ( n8195 , n5452 );
not ( n8196 , n4428 );
or ( n8197 , n8195 , n8196 );
or ( n8198 , n4428 , n5452 );
nand ( n8199 , n8197 , n8198 );
nand ( n8200 , n8194 , n8199 );
nor ( n8201 , n8189 , n8200 );
not ( n8202 , n5455 );
not ( n8203 , n4431 );
or ( n8204 , n8202 , n8203 );
or ( n8205 , n4431 , n5455 );
nand ( n8206 , n8204 , n8205 );
not ( n8207 , n5454 );
not ( n8208 , n4430 );
or ( n8209 , n8207 , n8208 );
or ( n8210 , n4430 , n5454 );
nand ( n8211 , n8209 , n8210 );
nand ( n8212 , n8206 , n8211 );
not ( n8213 , n5457 );
not ( n8214 , n4433 );
or ( n8215 , n8213 , n8214 );
or ( n8216 , n4433 , n5457 );
nand ( n8217 , n8215 , n8216 );
not ( n8218 , n5456 );
not ( n8219 , n4432 );
or ( n8220 , n8218 , n8219 );
or ( n8221 , n4432 , n5456 );
nand ( n8222 , n8220 , n8221 );
nand ( n8223 , n8217 , n8222 );
nor ( n8224 , n8212 , n8223 );
not ( n8225 , n5459 );
not ( n8226 , n4435 );
or ( n8227 , n8225 , n8226 );
or ( n8228 , n4435 , n5459 );
nand ( n8229 , n8227 , n8228 );
not ( n8230 , n5458 );
not ( n8231 , n4434 );
or ( n8232 , n8230 , n8231 );
or ( n8233 , n4434 , n5458 );
nand ( n8234 , n8232 , n8233 );
nand ( n8235 , n8229 , n8234 );
not ( n8236 , n5461 );
not ( n8237 , n4437 );
or ( n8238 , n8236 , n8237 );
or ( n8239 , n4437 , n5461 );
nand ( n8240 , n8238 , n8239 );
not ( n8241 , n5460 );
not ( n8242 , n4436 );
or ( n8243 , n8241 , n8242 );
or ( n8244 , n4436 , n5460 );
nand ( n8245 , n8243 , n8244 );
nand ( n8246 , n8240 , n8245 );
nor ( n8247 , n8235 , n8246 );
not ( n8248 , n5447 );
not ( n8249 , n4423 );
or ( n8250 , n8248 , n8249 );
or ( n8251 , n4423 , n5447 );
nand ( n8252 , n8250 , n8251 );
not ( n8253 , n5446 );
not ( n8254 , n4422 );
or ( n8255 , n8253 , n8254 );
or ( n8256 , n4422 , n5446 );
nand ( n8257 , n8255 , n8256 );
nand ( n8258 , n8252 , n8257 );
not ( n8259 , n5449 );
not ( n8260 , n4425 );
or ( n8261 , n8259 , n8260 );
or ( n8262 , n4425 , n5449 );
nand ( n8263 , n8261 , n8262 );
not ( n8264 , n5448 );
not ( n8265 , n4424 );
or ( n8266 , n8264 , n8265 );
or ( n8267 , n4424 , n5448 );
nand ( n8268 , n8266 , n8267 );
nand ( n8269 , n8263 , n8268 );
nor ( n8270 , n8258 , n8269 );
nand ( n8271 , n8201 , n8224 , n8247 , n8270 );
not ( n8272 , n5471 );
not ( n8273 , n4447 );
or ( n8274 , n8272 , n8273 );
or ( n8275 , n4447 , n5471 );
nand ( n8276 , n8274 , n8275 );
not ( n8277 , n5470 );
not ( n8278 , n4446 );
or ( n8279 , n8277 , n8278 );
or ( n8280 , n4446 , n5470 );
nand ( n8281 , n8279 , n8280 );
nand ( n8282 , n8276 , n8281 );
not ( n8283 , n5473 );
not ( n8284 , n4449 );
or ( n8285 , n8283 , n8284 );
or ( n8286 , n4449 , n5473 );
nand ( n8287 , n8285 , n8286 );
not ( n8288 , n5472 );
not ( n8289 , n4448 );
or ( n8290 , n8288 , n8289 );
or ( n8291 , n4448 , n5472 );
nand ( n8292 , n8290 , n8291 );
nand ( n8293 , n8287 , n8292 );
nor ( n8294 , n8282 , n8293 );
not ( n8295 , n5475 );
not ( n8296 , n4451 );
or ( n8297 , n8295 , n8296 );
or ( n8298 , n4451 , n5475 );
nand ( n8299 , n8297 , n8298 );
not ( n8300 , n5474 );
not ( n8301 , n4450 );
or ( n8302 , n8300 , n8301 );
or ( n8303 , n4450 , n5474 );
nand ( n8304 , n8302 , n8303 );
nand ( n8305 , n8299 , n8304 );
not ( n8306 , n5477 );
not ( n8307 , n4453 );
or ( n8308 , n8306 , n8307 );
or ( n8309 , n4453 , n5477 );
nand ( n8310 , n8308 , n8309 );
not ( n8311 , n5476 );
not ( n8312 , n4452 );
or ( n8313 , n8311 , n8312 );
or ( n8314 , n4452 , n5476 );
nand ( n8315 , n8313 , n8314 );
nand ( n8316 , n8310 , n8315 );
nor ( n8317 , n8305 , n8316 );
not ( n8318 , n5467 );
not ( n8319 , n4443 );
or ( n8320 , n8318 , n8319 );
or ( n8321 , n4443 , n5467 );
nand ( n8322 , n8320 , n8321 );
not ( n8323 , n5466 );
not ( n8324 , n4442 );
or ( n8325 , n8323 , n8324 );
or ( n8326 , n4442 , n5466 );
nand ( n8327 , n8325 , n8326 );
nand ( n8328 , n8322 , n8327 );
not ( n8329 , n5469 );
not ( n8330 , n4445 );
or ( n8331 , n8329 , n8330 );
or ( n8332 , n4445 , n5469 );
nand ( n8333 , n8331 , n8332 );
not ( n8334 , n5468 );
not ( n8335 , n4444 );
or ( n8336 , n8334 , n8335 );
or ( n8337 , n4444 , n5468 );
nand ( n8338 , n8336 , n8337 );
nand ( n8339 , n8333 , n8338 );
nor ( n8340 , n8328 , n8339 );
not ( n8341 , n5463 );
not ( n8342 , n4439 );
or ( n8343 , n8341 , n8342 );
or ( n8344 , n4439 , n5463 );
nand ( n8345 , n8343 , n8344 );
not ( n8346 , n5462 );
not ( n8347 , n4438 );
or ( n8348 , n8346 , n8347 );
or ( n8349 , n4438 , n5462 );
nand ( n8350 , n8348 , n8349 );
nand ( n8351 , n8345 , n8350 );
not ( n8352 , n5465 );
not ( n8353 , n4441 );
or ( n8354 , n8352 , n8353 );
or ( n8355 , n4441 , n5465 );
nand ( n8356 , n8354 , n8355 );
not ( n8357 , n5464 );
not ( n8358 , n4440 );
or ( n8359 , n8357 , n8358 );
or ( n8360 , n4440 , n5464 );
nand ( n8361 , n8359 , n8360 );
nand ( n8362 , n8356 , n8361 );
nor ( n8363 , n8351 , n8362 );
nand ( n8364 , n8294 , n8317 , n8340 , n8363 );
nor ( n8365 , n8271 , n8364 );
nand ( n8366 , n7806 , n7991 , n8178 , n8365 );
not ( n8367 , n5539 );
not ( n8368 , n4515 );
or ( n8369 , n8367 , n8368 );
or ( n8370 , n4515 , n5539 );
nand ( n8371 , n8369 , n8370 );
not ( n8372 , n5538 );
not ( n8373 , n4514 );
or ( n8374 , n8372 , n8373 );
or ( n8375 , n4514 , n5538 );
nand ( n8376 , n8374 , n8375 );
nand ( n8377 , n8371 , n8376 );
not ( n8378 , n5541 );
not ( n8379 , n4517 );
or ( n8380 , n8378 , n8379 );
or ( n8381 , n4517 , n5541 );
nand ( n8382 , n8380 , n8381 );
not ( n8383 , n5540 );
not ( n8384 , n4516 );
or ( n8385 , n8383 , n8384 );
or ( n8386 , n4516 , n5540 );
nand ( n8387 , n8385 , n8386 );
nand ( n8388 , n8382 , n8387 );
nor ( n8389 , n8377 , n8388 );
not ( n8390 , n5535 );
not ( n8391 , n4511 );
or ( n8392 , n8390 , n8391 );
or ( n8393 , n4511 , n5535 );
nand ( n8394 , n8392 , n8393 );
not ( n8395 , n5534 );
not ( n8396 , n4510 );
or ( n8397 , n8395 , n8396 );
or ( n8398 , n4510 , n5534 );
nand ( n8399 , n8397 , n8398 );
nand ( n8400 , n8394 , n8399 );
not ( n8401 , n5537 );
not ( n8402 , n4513 );
or ( n8403 , n8401 , n8402 );
or ( n8404 , n4513 , n5537 );
nand ( n8405 , n8403 , n8404 );
not ( n8406 , n5536 );
not ( n8407 , n4512 );
or ( n8408 , n8406 , n8407 );
or ( n8409 , n4512 , n5536 );
nand ( n8410 , n8408 , n8409 );
nand ( n8411 , n8405 , n8410 );
nor ( n8412 , n8400 , n8411 );
not ( n8413 , n5531 );
not ( n8414 , n4507 );
or ( n8415 , n8413 , n8414 );
or ( n8416 , n4507 , n5531 );
nand ( n8417 , n8415 , n8416 );
not ( n8418 , n5530 );
not ( n8419 , n4506 );
or ( n8420 , n8418 , n8419 );
or ( n8421 , n4506 , n5530 );
nand ( n8422 , n8420 , n8421 );
nand ( n8423 , n8417 , n8422 );
not ( n8424 , n5533 );
not ( n8425 , n4509 );
or ( n8426 , n8424 , n8425 );
or ( n8427 , n4509 , n5533 );
nand ( n8428 , n8426 , n8427 );
not ( n8429 , n5532 );
not ( n8430 , n4508 );
or ( n8431 , n8429 , n8430 );
or ( n8432 , n4508 , n5532 );
nand ( n8433 , n8431 , n8432 );
nand ( n8434 , n8428 , n8433 );
nor ( n8435 , n8423 , n8434 );
not ( n8436 , n5527 );
not ( n8437 , n4503 );
or ( n8438 , n8436 , n8437 );
or ( n8439 , n4503 , n5527 );
nand ( n8440 , n8438 , n8439 );
not ( n8441 , n5526 );
not ( n8442 , n4502 );
or ( n8443 , n8441 , n8442 );
or ( n8444 , n4502 , n5526 );
nand ( n8445 , n8443 , n8444 );
nand ( n8446 , n8440 , n8445 );
not ( n8447 , n5529 );
not ( n8448 , n4505 );
or ( n8449 , n8447 , n8448 );
or ( n8450 , n4505 , n5529 );
nand ( n8451 , n8449 , n8450 );
not ( n8452 , n5528 );
not ( n8453 , n4504 );
or ( n8454 , n8452 , n8453 );
or ( n8455 , n4504 , n5528 );
nand ( n8456 , n8454 , n8455 );
nand ( n8457 , n8451 , n8456 );
nor ( n8458 , n8446 , n8457 );
nand ( n8459 , n8389 , n8412 , n8435 , n8458 );
not ( n8460 , n5523 );
not ( n8461 , n4499 );
or ( n8462 , n8460 , n8461 );
or ( n8463 , n4499 , n5523 );
nand ( n8464 , n8462 , n8463 );
not ( n8465 , n5522 );
not ( n8466 , n4498 );
or ( n8467 , n8465 , n8466 );
or ( n8468 , n4498 , n5522 );
nand ( n8469 , n8467 , n8468 );
nand ( n8470 , n8464 , n8469 );
not ( n8471 , n5525 );
not ( n8472 , n4501 );
or ( n8473 , n8471 , n8472 );
or ( n8474 , n4501 , n5525 );
nand ( n8475 , n8473 , n8474 );
not ( n8476 , n5524 );
not ( n8477 , n4500 );
or ( n8478 , n8476 , n8477 );
or ( n8479 , n4500 , n5524 );
nand ( n8480 , n8478 , n8479 );
nand ( n8481 , n8475 , n8480 );
nor ( n8482 , n8470 , n8481 );
not ( n8483 , n5519 );
not ( n8484 , n4495 );
or ( n8485 , n8483 , n8484 );
or ( n8486 , n4495 , n5519 );
nand ( n8487 , n8485 , n8486 );
not ( n8488 , n5518 );
not ( n8489 , n4494 );
or ( n8490 , n8488 , n8489 );
or ( n8491 , n4494 , n5518 );
nand ( n8492 , n8490 , n8491 );
nand ( n8493 , n8487 , n8492 );
not ( n8494 , n5521 );
not ( n8495 , n4497 );
or ( n8496 , n8494 , n8495 );
or ( n8497 , n4497 , n5521 );
nand ( n8498 , n8496 , n8497 );
not ( n8499 , n5520 );
not ( n8500 , n4496 );
or ( n8501 , n8499 , n8500 );
or ( n8502 , n4496 , n5520 );
nand ( n8503 , n8501 , n8502 );
nand ( n8504 , n8498 , n8503 );
nor ( n8505 , n8493 , n8504 );
not ( n8506 , n5513 );
not ( n8507 , n4489 );
or ( n8508 , n8506 , n8507 );
or ( n8509 , n4489 , n5513 );
nand ( n8510 , n8508 , n8509 );
not ( n8511 , n5512 );
not ( n8512 , n4488 );
or ( n8513 , n8511 , n8512 );
or ( n8514 , n4488 , n5512 );
nand ( n8515 , n8513 , n8514 );
nand ( n8516 , n8510 , n8515 );
not ( n8517 , n5511 );
not ( n8518 , n4487 );
or ( n8519 , n8517 , n8518 );
or ( n8520 , n4487 , n5511 );
nand ( n8521 , n8519 , n8520 );
not ( n8522 , n5510 );
not ( n8523 , n4486 );
or ( n8524 , n8522 , n8523 );
or ( n8525 , n4486 , n5510 );
nand ( n8526 , n8524 , n8525 );
nand ( n8527 , n8521 , n8526 );
nor ( n8528 , n8516 , n8527 );
not ( n8529 , n5516 );
not ( n8530 , n4492 );
or ( n8531 , n8529 , n8530 );
or ( n8532 , n4492 , n5516 );
nand ( n8533 , n8531 , n8532 );
not ( n8534 , n5517 );
not ( n8535 , n4493 );
or ( n8536 , n8534 , n8535 );
or ( n8537 , n4493 , n5517 );
nand ( n8538 , n8536 , n8537 );
not ( n8539 , n5514 );
not ( n8540 , n4490 );
or ( n8541 , n8539 , n8540 );
or ( n8542 , n4490 , n5514 );
nand ( n8543 , n8541 , n8542 );
not ( n8544 , n5515 );
not ( n8545 , n4491 );
or ( n8546 , n8544 , n8545 );
or ( n8547 , n4491 , n5515 );
nand ( n8548 , n8546 , n8547 );
and ( n8549 , n8533 , n8538 , n8543 , n8548 );
nand ( n8550 , n8482 , n8505 , n8528 , n8549 );
nor ( n8551 , n8459 , n8550 );
not ( n8552 , n5555 );
not ( n8553 , n4531 );
or ( n8554 , n8552 , n8553 );
or ( n8555 , n4531 , n5555 );
nand ( n8556 , n8554 , n8555 );
not ( n8557 , n5554 );
not ( n8558 , n4530 );
or ( n8559 , n8557 , n8558 );
or ( n8560 , n4530 , n5554 );
nand ( n8561 , n8559 , n8560 );
nand ( n8562 , n8556 , n8561 );
not ( n8563 , n5557 );
not ( n8564 , n4533 );
or ( n8565 , n8563 , n8564 );
or ( n8566 , n4533 , n5557 );
nand ( n8567 , n8565 , n8566 );
not ( n8568 , n5556 );
not ( n8569 , n4532 );
or ( n8570 , n8568 , n8569 );
or ( n8571 , n4532 , n5556 );
nand ( n8572 , n8570 , n8571 );
nand ( n8573 , n8567 , n8572 );
nor ( n8574 , n8562 , n8573 );
not ( n8575 , n5551 );
not ( n8576 , n4527 );
or ( n8577 , n8575 , n8576 );
or ( n8578 , n4527 , n5551 );
nand ( n8579 , n8577 , n8578 );
not ( n8580 , n5550 );
not ( n8581 , n4526 );
or ( n8582 , n8580 , n8581 );
or ( n8583 , n4526 , n5550 );
nand ( n8584 , n8582 , n8583 );
nand ( n8585 , n8579 , n8584 );
not ( n8586 , n5553 );
not ( n8587 , n4529 );
or ( n8588 , n8586 , n8587 );
or ( n8589 , n4529 , n5553 );
nand ( n8590 , n8588 , n8589 );
not ( n8591 , n5552 );
not ( n8592 , n4528 );
or ( n8593 , n8591 , n8592 );
or ( n8594 , n4528 , n5552 );
nand ( n8595 , n8593 , n8594 );
nand ( n8596 , n8590 , n8595 );
nor ( n8597 , n8585 , n8596 );
not ( n8598 , n5547 );
not ( n8599 , n4523 );
or ( n8600 , n8598 , n8599 );
or ( n8601 , n4523 , n5547 );
nand ( n8602 , n8600 , n8601 );
not ( n8603 , n5546 );
not ( n8604 , n4522 );
or ( n8605 , n8603 , n8604 );
or ( n8606 , n4522 , n5546 );
nand ( n8607 , n8605 , n8606 );
nand ( n8608 , n8602 , n8607 );
not ( n8609 , n5549 );
not ( n8610 , n4525 );
or ( n8611 , n8609 , n8610 );
or ( n8612 , n4525 , n5549 );
nand ( n8613 , n8611 , n8612 );
not ( n8614 , n5548 );
not ( n8615 , n4524 );
or ( n8616 , n8614 , n8615 );
or ( n8617 , n4524 , n5548 );
nand ( n8618 , n8616 , n8617 );
nand ( n8619 , n8613 , n8618 );
nor ( n8620 , n8608 , n8619 );
not ( n8621 , n5543 );
not ( n8622 , n4519 );
or ( n8623 , n8621 , n8622 );
or ( n8624 , n4519 , n5543 );
nand ( n8625 , n8623 , n8624 );
not ( n8626 , n5542 );
not ( n8627 , n4518 );
or ( n8628 , n8626 , n8627 );
or ( n8629 , n4518 , n5542 );
nand ( n8630 , n8628 , n8629 );
nand ( n8631 , n8625 , n8630 );
not ( n8632 , n5545 );
not ( n8633 , n4521 );
or ( n8634 , n8632 , n8633 );
or ( n8635 , n4521 , n5545 );
nand ( n8636 , n8634 , n8635 );
not ( n8637 , n5544 );
not ( n8638 , n4520 );
or ( n8639 , n8637 , n8638 );
or ( n8640 , n4520 , n5544 );
nand ( n8641 , n8639 , n8640 );
nand ( n8642 , n8636 , n8641 );
nor ( n8643 , n8631 , n8642 );
nand ( n8644 , n8574 , n8597 , n8620 , n8643 );
not ( n8645 , n5571 );
not ( n8646 , n4547 );
or ( n8647 , n8645 , n8646 );
or ( n8648 , n4547 , n5571 );
nand ( n8649 , n8647 , n8648 );
not ( n8650 , n5570 );
not ( n8651 , n4546 );
or ( n8652 , n8650 , n8651 );
or ( n8653 , n4546 , n5570 );
nand ( n8654 , n8652 , n8653 );
nand ( n8655 , n8649 , n8654 );
not ( n8656 , n5573 );
not ( n8657 , n4549 );
or ( n8658 , n8656 , n8657 );
or ( n8659 , n4549 , n5573 );
nand ( n8660 , n8658 , n8659 );
not ( n8661 , n5572 );
not ( n8662 , n4548 );
or ( n8663 , n8661 , n8662 );
or ( n8664 , n4548 , n5572 );
nand ( n8665 , n8663 , n8664 );
nand ( n8666 , n8660 , n8665 );
nor ( n8667 , n8655 , n8666 );
not ( n8668 , n5567 );
not ( n8669 , n4543 );
or ( n8670 , n8668 , n8669 );
or ( n8671 , n4543 , n5567 );
nand ( n8672 , n8670 , n8671 );
not ( n8673 , n5566 );
not ( n8674 , n4542 );
or ( n8675 , n8673 , n8674 );
or ( n8676 , n4542 , n5566 );
nand ( n8677 , n8675 , n8676 );
nand ( n8678 , n8672 , n8677 );
not ( n8679 , n5569 );
not ( n8680 , n4545 );
or ( n8681 , n8679 , n8680 );
or ( n8682 , n4545 , n5569 );
nand ( n8683 , n8681 , n8682 );
not ( n8684 , n5568 );
not ( n8685 , n4544 );
or ( n8686 , n8684 , n8685 );
or ( n8687 , n4544 , n5568 );
nand ( n8688 , n8686 , n8687 );
nand ( n8689 , n8683 , n8688 );
nor ( n8690 , n8678 , n8689 );
not ( n8691 , n5563 );
not ( n8692 , n4539 );
or ( n8693 , n8691 , n8692 );
or ( n8694 , n4539 , n5563 );
nand ( n8695 , n8693 , n8694 );
not ( n8696 , n5562 );
not ( n8697 , n4538 );
or ( n8698 , n8696 , n8697 );
or ( n8699 , n4538 , n5562 );
nand ( n8700 , n8698 , n8699 );
nand ( n8701 , n8695 , n8700 );
not ( n8702 , n5565 );
not ( n8703 , n4541 );
or ( n8704 , n8702 , n8703 );
or ( n8705 , n4541 , n5565 );
nand ( n8706 , n8704 , n8705 );
not ( n8707 , n5564 );
not ( n8708 , n4540 );
or ( n8709 , n8707 , n8708 );
or ( n8710 , n4540 , n5564 );
nand ( n8711 , n8709 , n8710 );
nand ( n8712 , n8706 , n8711 );
nor ( n8713 , n8701 , n8712 );
not ( n8714 , n5559 );
not ( n8715 , n4535 );
or ( n8716 , n8714 , n8715 );
or ( n8717 , n4535 , n5559 );
nand ( n8718 , n8716 , n8717 );
not ( n8719 , n5558 );
not ( n8720 , n4534 );
or ( n8721 , n8719 , n8720 );
or ( n8722 , n4534 , n5558 );
nand ( n8723 , n8721 , n8722 );
nand ( n8724 , n8718 , n8723 );
not ( n8725 , n5561 );
not ( n8726 , n4537 );
or ( n8727 , n8725 , n8726 );
or ( n8728 , n4537 , n5561 );
nand ( n8729 , n8727 , n8728 );
not ( n8730 , n5560 );
not ( n8731 , n4536 );
or ( n8732 , n8730 , n8731 );
or ( n8733 , n4536 , n5560 );
nand ( n8734 , n8732 , n8733 );
nand ( n8735 , n8729 , n8734 );
nor ( n8736 , n8724 , n8735 );
nand ( n8737 , n8667 , n8690 , n8713 , n8736 );
nor ( n8738 , n8644 , n8737 );
not ( n8739 , n5583 );
not ( n8740 , n4559 );
or ( n8741 , n8739 , n8740 );
or ( n8742 , n4559 , n5583 );
nand ( n8743 , n8741 , n8742 );
not ( n8744 , n5582 );
not ( n8745 , n4558 );
or ( n8746 , n8744 , n8745 );
or ( n8747 , n4558 , n5582 );
nand ( n8748 , n8746 , n8747 );
nand ( n8749 , n8743 , n8748 );
not ( n8750 , n5585 );
not ( n8751 , n4561 );
or ( n8752 , n8750 , n8751 );
or ( n8753 , n4561 , n5585 );
nand ( n8754 , n8752 , n8753 );
not ( n8755 , n5584 );
not ( n8756 , n4560 );
or ( n8757 , n8755 , n8756 );
or ( n8758 , n4560 , n5584 );
nand ( n8759 , n8757 , n8758 );
nand ( n8760 , n8754 , n8759 );
nor ( n8761 , n8749 , n8760 );
not ( n8762 , n5587 );
not ( n8763 , n4563 );
or ( n8764 , n8762 , n8763 );
or ( n8765 , n4563 , n5587 );
nand ( n8766 , n8764 , n8765 );
not ( n8767 , n5586 );
not ( n8768 , n4562 );
or ( n8769 , n8767 , n8768 );
or ( n8770 , n4562 , n5586 );
nand ( n8771 , n8769 , n8770 );
nand ( n8772 , n8766 , n8771 );
not ( n8773 , n5589 );
not ( n8774 , n4565 );
or ( n8775 , n8773 , n8774 );
or ( n8776 , n4565 , n5589 );
nand ( n8777 , n8775 , n8776 );
not ( n8778 , n5588 );
not ( n8779 , n4564 );
or ( n8780 , n8778 , n8779 );
or ( n8781 , n4564 , n5588 );
nand ( n8782 , n8780 , n8781 );
nand ( n8783 , n8777 , n8782 );
nor ( n8784 , n8772 , n8783 );
not ( n8785 , n5579 );
not ( n8786 , n4555 );
or ( n8787 , n8785 , n8786 );
or ( n8788 , n4555 , n5579 );
nand ( n8789 , n8787 , n8788 );
not ( n8790 , n5578 );
not ( n8791 , n4554 );
or ( n8792 , n8790 , n8791 );
or ( n8793 , n4554 , n5578 );
nand ( n8794 , n8792 , n8793 );
nand ( n8795 , n8789 , n8794 );
not ( n8796 , n5581 );
not ( n8797 , n4557 );
or ( n8798 , n8796 , n8797 );
or ( n8799 , n4557 , n5581 );
nand ( n8800 , n8798 , n8799 );
not ( n8801 , n5580 );
not ( n8802 , n4556 );
or ( n8803 , n8801 , n8802 );
or ( n8804 , n4556 , n5580 );
nand ( n8805 , n8803 , n8804 );
nand ( n8806 , n8800 , n8805 );
nor ( n8807 , n8795 , n8806 );
not ( n8808 , n5575 );
not ( n8809 , n4551 );
or ( n8810 , n8808 , n8809 );
or ( n8811 , n4551 , n5575 );
nand ( n8812 , n8810 , n8811 );
not ( n8813 , n5574 );
not ( n8814 , n4550 );
or ( n8815 , n8813 , n8814 );
or ( n8816 , n4550 , n5574 );
nand ( n8817 , n8815 , n8816 );
nand ( n8818 , n8812 , n8817 );
not ( n8819 , n5577 );
not ( n8820 , n4553 );
or ( n8821 , n8819 , n8820 );
or ( n8822 , n4553 , n5577 );
nand ( n8823 , n8821 , n8822 );
not ( n8824 , n5576 );
not ( n8825 , n4552 );
or ( n8826 , n8824 , n8825 );
or ( n8827 , n4552 , n5576 );
nand ( n8828 , n8826 , n8827 );
nand ( n8829 , n8823 , n8828 );
nor ( n8830 , n8818 , n8829 );
nand ( n8831 , n8761 , n8784 , n8807 , n8830 );
not ( n8832 , n5603 );
not ( n8833 , n4579 );
or ( n8834 , n8832 , n8833 );
or ( n8835 , n4579 , n5603 );
nand ( n8836 , n8834 , n8835 );
not ( n8837 , n5602 );
not ( n8838 , n4578 );
or ( n8839 , n8837 , n8838 );
or ( n8840 , n4578 , n5602 );
nand ( n8841 , n8839 , n8840 );
nand ( n8842 , n8836 , n8841 );
not ( n8843 , n5605 );
not ( n8844 , n4581 );
or ( n8845 , n8843 , n8844 );
or ( n8846 , n4581 , n5605 );
nand ( n8847 , n8845 , n8846 );
not ( n8848 , n5604 );
not ( n8849 , n4580 );
or ( n8850 , n8848 , n8849 );
or ( n8851 , n4580 , n5604 );
nand ( n8852 , n8850 , n8851 );
nand ( n8853 , n8847 , n8852 );
nor ( n8854 , n8842 , n8853 );
not ( n8855 , n5599 );
not ( n8856 , n4575 );
or ( n8857 , n8855 , n8856 );
or ( n8858 , n4575 , n5599 );
nand ( n8859 , n8857 , n8858 );
not ( n8860 , n5598 );
not ( n8861 , n4574 );
or ( n8862 , n8860 , n8861 );
or ( n8863 , n4574 , n5598 );
nand ( n8864 , n8862 , n8863 );
nand ( n8865 , n8859 , n8864 );
not ( n8866 , n5601 );
not ( n8867 , n4577 );
or ( n8868 , n8866 , n8867 );
or ( n8869 , n4577 , n5601 );
nand ( n8870 , n8868 , n8869 );
not ( n8871 , n5600 );
not ( n8872 , n4576 );
or ( n8873 , n8871 , n8872 );
or ( n8874 , n4576 , n5600 );
nand ( n8875 , n8873 , n8874 );
nand ( n8876 , n8870 , n8875 );
nor ( n8877 , n8865 , n8876 );
not ( n8878 , n5595 );
not ( n8879 , n4571 );
or ( n8880 , n8878 , n8879 );
or ( n8881 , n4571 , n5595 );
nand ( n8882 , n8880 , n8881 );
not ( n8883 , n5594 );
not ( n8884 , n4570 );
or ( n8885 , n8883 , n8884 );
or ( n8886 , n4570 , n5594 );
nand ( n8887 , n8885 , n8886 );
nand ( n8888 , n8882 , n8887 );
not ( n8889 , n5597 );
not ( n8890 , n4573 );
or ( n8891 , n8889 , n8890 );
or ( n8892 , n4573 , n5597 );
nand ( n8893 , n8891 , n8892 );
not ( n8894 , n5596 );
not ( n8895 , n4572 );
or ( n8896 , n8894 , n8895 );
or ( n8897 , n4572 , n5596 );
nand ( n8898 , n8896 , n8897 );
nand ( n8899 , n8893 , n8898 );
nor ( n8900 , n8888 , n8899 );
not ( n8901 , n5591 );
not ( n8902 , n4567 );
or ( n8903 , n8901 , n8902 );
or ( n8904 , n4567 , n5591 );
nand ( n8905 , n8903 , n8904 );
not ( n8906 , n5590 );
not ( n8907 , n4566 );
or ( n8908 , n8906 , n8907 );
or ( n8909 , n4566 , n5590 );
nand ( n8910 , n8908 , n8909 );
nand ( n8911 , n8905 , n8910 );
not ( n8912 , n5593 );
not ( n8913 , n4569 );
or ( n8914 , n8912 , n8913 );
or ( n8915 , n4569 , n5593 );
nand ( n8916 , n8914 , n8915 );
not ( n8917 , n5592 );
not ( n8918 , n4568 );
or ( n8919 , n8917 , n8918 );
or ( n8920 , n4568 , n5592 );
nand ( n8921 , n8919 , n8920 );
nand ( n8922 , n8916 , n8921 );
nor ( n8923 , n8911 , n8922 );
nand ( n8924 , n8854 , n8877 , n8900 , n8923 );
nor ( n8925 , n8831 , n8924 );
not ( n8926 , n5619 );
not ( n8927 , n4595 );
or ( n8928 , n8926 , n8927 );
or ( n8929 , n4595 , n5619 );
nand ( n8930 , n8928 , n8929 );
not ( n8931 , n5618 );
not ( n8932 , n4594 );
or ( n8933 , n8931 , n8932 );
or ( n8934 , n4594 , n5618 );
nand ( n8935 , n8933 , n8934 );
nand ( n8936 , n8930 , n8935 );
not ( n8937 , n5621 );
not ( n8938 , n4597 );
or ( n8939 , n8937 , n8938 );
or ( n8940 , n4597 , n5621 );
nand ( n8941 , n8939 , n8940 );
not ( n8942 , n5620 );
not ( n8943 , n4596 );
or ( n8944 , n8942 , n8943 );
or ( n8945 , n4596 , n5620 );
nand ( n8946 , n8944 , n8945 );
nand ( n8947 , n8941 , n8946 );
nor ( n8948 , n8936 , n8947 );
not ( n8949 , n5615 );
not ( n8950 , n4591 );
or ( n8951 , n8949 , n8950 );
or ( n8952 , n4591 , n5615 );
nand ( n8953 , n8951 , n8952 );
not ( n8954 , n5614 );
not ( n8955 , n4590 );
or ( n8956 , n8954 , n8955 );
or ( n8957 , n4590 , n5614 );
nand ( n8958 , n8956 , n8957 );
nand ( n8959 , n8953 , n8958 );
not ( n8960 , n5617 );
not ( n8961 , n4593 );
or ( n8962 , n8960 , n8961 );
or ( n8963 , n4593 , n5617 );
nand ( n8964 , n8962 , n8963 );
not ( n8965 , n5616 );
not ( n8966 , n4592 );
or ( n8967 , n8965 , n8966 );
or ( n8968 , n4592 , n5616 );
nand ( n8969 , n8967 , n8968 );
nand ( n8970 , n8964 , n8969 );
nor ( n8971 , n8959 , n8970 );
not ( n8972 , n5611 );
not ( n8973 , n4587 );
or ( n8974 , n8972 , n8973 );
or ( n8975 , n4587 , n5611 );
nand ( n8976 , n8974 , n8975 );
not ( n8977 , n5610 );
not ( n8978 , n4586 );
or ( n8979 , n8977 , n8978 );
or ( n8980 , n4586 , n5610 );
nand ( n8981 , n8979 , n8980 );
nand ( n8982 , n8976 , n8981 );
not ( n8983 , n5613 );
not ( n8984 , n4589 );
or ( n8985 , n8983 , n8984 );
or ( n8986 , n4589 , n5613 );
nand ( n8987 , n8985 , n8986 );
not ( n8988 , n5612 );
not ( n8989 , n4588 );
or ( n8990 , n8988 , n8989 );
or ( n8991 , n4588 , n5612 );
nand ( n8992 , n8990 , n8991 );
nand ( n8993 , n8987 , n8992 );
nor ( n8994 , n8982 , n8993 );
not ( n8995 , n5607 );
not ( n8996 , n4583 );
or ( n8997 , n8995 , n8996 );
or ( n8998 , n4583 , n5607 );
nand ( n8999 , n8997 , n8998 );
not ( n9000 , n5606 );
not ( n9001 , n4582 );
or ( n9002 , n9000 , n9001 );
or ( n9003 , n4582 , n5606 );
nand ( n9004 , n9002 , n9003 );
nand ( n9005 , n8999 , n9004 );
not ( n9006 , n5609 );
not ( n9007 , n4585 );
or ( n9008 , n9006 , n9007 );
or ( n9009 , n4585 , n5609 );
nand ( n9010 , n9008 , n9009 );
not ( n9011 , n5608 );
not ( n9012 , n4584 );
or ( n9013 , n9011 , n9012 );
or ( n9014 , n4584 , n5608 );
nand ( n9015 , n9013 , n9014 );
nand ( n9016 , n9010 , n9015 );
nor ( n9017 , n9005 , n9016 );
nand ( n9018 , n8948 , n8971 , n8994 , n9017 );
not ( n9019 , n5635 );
not ( n9020 , n4611 );
or ( n9021 , n9019 , n9020 );
or ( n9022 , n4611 , n5635 );
nand ( n9023 , n9021 , n9022 );
not ( n9024 , n5634 );
not ( n9025 , n4610 );
or ( n9026 , n9024 , n9025 );
or ( n9027 , n4610 , n5634 );
nand ( n9028 , n9026 , n9027 );
nand ( n9029 , n9023 , n9028 );
not ( n9030 , n5637 );
not ( n9031 , n4613 );
or ( n9032 , n9030 , n9031 );
or ( n9033 , n4613 , n5637 );
nand ( n9034 , n9032 , n9033 );
not ( n9035 , n5636 );
not ( n9036 , n4612 );
or ( n9037 , n9035 , n9036 );
or ( n9038 , n4612 , n5636 );
nand ( n9039 , n9037 , n9038 );
nand ( n9040 , n9034 , n9039 );
nor ( n9041 , n9029 , n9040 );
not ( n9042 , n5631 );
not ( n9043 , n4607 );
or ( n9044 , n9042 , n9043 );
or ( n9045 , n4607 , n5631 );
nand ( n9046 , n9044 , n9045 );
not ( n9047 , n5630 );
not ( n9048 , n4606 );
or ( n9049 , n9047 , n9048 );
or ( n9050 , n4606 , n5630 );
nand ( n9051 , n9049 , n9050 );
nand ( n9052 , n9046 , n9051 );
not ( n9053 , n5633 );
not ( n9054 , n4609 );
or ( n9055 , n9053 , n9054 );
or ( n9056 , n4609 , n5633 );
nand ( n9057 , n9055 , n9056 );
not ( n9058 , n5632 );
not ( n9059 , n4608 );
or ( n9060 , n9058 , n9059 );
or ( n9061 , n4608 , n5632 );
nand ( n9062 , n9060 , n9061 );
nand ( n9063 , n9057 , n9062 );
nor ( n9064 , n9052 , n9063 );
not ( n9065 , n5627 );
not ( n9066 , n4603 );
or ( n9067 , n9065 , n9066 );
or ( n9068 , n4603 , n5627 );
nand ( n9069 , n9067 , n9068 );
not ( n9070 , n5626 );
not ( n9071 , n4602 );
or ( n9072 , n9070 , n9071 );
or ( n9073 , n4602 , n5626 );
nand ( n9074 , n9072 , n9073 );
nand ( n9075 , n9069 , n9074 );
not ( n9076 , n5629 );
not ( n9077 , n4605 );
or ( n9078 , n9076 , n9077 );
or ( n9079 , n4605 , n5629 );
nand ( n9080 , n9078 , n9079 );
not ( n9081 , n5628 );
not ( n9082 , n4604 );
or ( n9083 , n9081 , n9082 );
or ( n9084 , n4604 , n5628 );
nand ( n9085 , n9083 , n9084 );
nand ( n9086 , n9080 , n9085 );
nor ( n9087 , n9075 , n9086 );
not ( n9088 , n5623 );
not ( n9089 , n4599 );
or ( n9090 , n9088 , n9089 );
or ( n9091 , n4599 , n5623 );
nand ( n9092 , n9090 , n9091 );
not ( n9093 , n5622 );
not ( n9094 , n4598 );
or ( n9095 , n9093 , n9094 );
or ( n9096 , n4598 , n5622 );
nand ( n9097 , n9095 , n9096 );
nand ( n9098 , n9092 , n9097 );
not ( n9099 , n5625 );
not ( n9100 , n4601 );
or ( n9101 , n9099 , n9100 );
or ( n9102 , n4601 , n5625 );
nand ( n9103 , n9101 , n9102 );
not ( n9104 , n5624 );
not ( n9105 , n4600 );
or ( n9106 , n9104 , n9105 );
or ( n9107 , n4600 , n5624 );
nand ( n9108 , n9106 , n9107 );
nand ( n9109 , n9103 , n9108 );
nor ( n9110 , n9098 , n9109 );
nand ( n9111 , n9041 , n9064 , n9087 , n9110 );
nor ( n9112 , n9018 , n9111 );
nand ( n9113 , n8551 , n8738 , n8925 , n9112 );
nor ( n9114 , n8366 , n9113 );
not ( n9115 , n5651 );
not ( n9116 , n4627 );
or ( n9117 , n9115 , n9116 );
or ( n9118 , n4627 , n5651 );
nand ( n9119 , n9117 , n9118 );
not ( n9120 , n5650 );
not ( n9121 , n4626 );
or ( n9122 , n9120 , n9121 );
or ( n9123 , n4626 , n5650 );
nand ( n9124 , n9122 , n9123 );
nand ( n9125 , n9119 , n9124 );
not ( n9126 , n5653 );
not ( n9127 , n4629 );
or ( n9128 , n9126 , n9127 );
or ( n9129 , n4629 , n5653 );
nand ( n9130 , n9128 , n9129 );
not ( n9131 , n5652 );
not ( n9132 , n4628 );
or ( n9133 , n9131 , n9132 );
or ( n9134 , n4628 , n5652 );
nand ( n9135 , n9133 , n9134 );
nand ( n9136 , n9130 , n9135 );
nor ( n9137 , n9125 , n9136 );
not ( n9138 , n5647 );
not ( n9139 , n4623 );
or ( n9140 , n9138 , n9139 );
or ( n9141 , n4623 , n5647 );
nand ( n9142 , n9140 , n9141 );
not ( n9143 , n5646 );
not ( n9144 , n4622 );
or ( n9145 , n9143 , n9144 );
or ( n9146 , n4622 , n5646 );
nand ( n9147 , n9145 , n9146 );
nand ( n9148 , n9142 , n9147 );
not ( n9149 , n5649 );
not ( n9150 , n4625 );
or ( n9151 , n9149 , n9150 );
or ( n9152 , n4625 , n5649 );
nand ( n9153 , n9151 , n9152 );
not ( n9154 , n5648 );
not ( n9155 , n4624 );
or ( n9156 , n9154 , n9155 );
or ( n9157 , n4624 , n5648 );
nand ( n9158 , n9156 , n9157 );
nand ( n9159 , n9153 , n9158 );
nor ( n9160 , n9148 , n9159 );
not ( n9161 , n5641 );
not ( n9162 , n4617 );
or ( n9163 , n9161 , n9162 );
or ( n9164 , n4617 , n5641 );
nand ( n9165 , n9163 , n9164 );
not ( n9166 , n5640 );
not ( n9167 , n4616 );
or ( n9168 , n9166 , n9167 );
or ( n9169 , n4616 , n5640 );
nand ( n9170 , n9168 , n9169 );
nand ( n9171 , n9165 , n9170 );
not ( n9172 , n5639 );
not ( n9173 , n4615 );
or ( n9174 , n9172 , n9173 );
or ( n9175 , n4615 , n5639 );
nand ( n9176 , n9174 , n9175 );
not ( n9177 , n5638 );
not ( n9178 , n4614 );
or ( n9179 , n9177 , n9178 );
or ( n9180 , n4614 , n5638 );
nand ( n9181 , n9179 , n9180 );
nand ( n9182 , n9176 , n9181 );
nor ( n9183 , n9171 , n9182 );
not ( n9184 , n5644 );
not ( n9185 , n4620 );
or ( n9186 , n9184 , n9185 );
or ( n9187 , n4620 , n5644 );
nand ( n9188 , n9186 , n9187 );
not ( n9189 , n5645 );
not ( n9190 , n4621 );
or ( n9191 , n9189 , n9190 );
or ( n9192 , n4621 , n5645 );
nand ( n9193 , n9191 , n9192 );
not ( n9194 , n5642 );
not ( n9195 , n4618 );
or ( n9196 , n9194 , n9195 );
or ( n9197 , n4618 , n5642 );
nand ( n9198 , n9196 , n9197 );
not ( n9199 , n5643 );
not ( n9200 , n4619 );
or ( n9201 , n9199 , n9200 );
or ( n9202 , n4619 , n5643 );
nand ( n9203 , n9201 , n9202 );
and ( n9204 , n9188 , n9193 , n9198 , n9203 );
nand ( n9205 , n9137 , n9160 , n9183 , n9204 );
not ( n9206 , n5667 );
not ( n9207 , n4643 );
or ( n9208 , n9206 , n9207 );
or ( n9209 , n4643 , n5667 );
nand ( n9210 , n9208 , n9209 );
not ( n9211 , n5666 );
not ( n9212 , n4642 );
or ( n9213 , n9211 , n9212 );
or ( n9214 , n4642 , n5666 );
nand ( n9215 , n9213 , n9214 );
nand ( n9216 , n9210 , n9215 );
not ( n9217 , n5669 );
not ( n9218 , n4645 );
or ( n9219 , n9217 , n9218 );
or ( n9220 , n4645 , n5669 );
nand ( n9221 , n9219 , n9220 );
not ( n9222 , n5668 );
not ( n9223 , n4644 );
or ( n9224 , n9222 , n9223 );
or ( n9225 , n4644 , n5668 );
nand ( n9226 , n9224 , n9225 );
nand ( n9227 , n9221 , n9226 );
nor ( n9228 , n9216 , n9227 );
not ( n9229 , n5663 );
not ( n9230 , n4639 );
or ( n9231 , n9229 , n9230 );
or ( n9232 , n4639 , n5663 );
nand ( n9233 , n9231 , n9232 );
not ( n9234 , n5662 );
not ( n9235 , n4638 );
or ( n9236 , n9234 , n9235 );
or ( n9237 , n4638 , n5662 );
nand ( n9238 , n9236 , n9237 );
nand ( n9239 , n9233 , n9238 );
not ( n9240 , n5665 );
not ( n9241 , n4641 );
or ( n9242 , n9240 , n9241 );
or ( n9243 , n4641 , n5665 );
nand ( n9244 , n9242 , n9243 );
not ( n9245 , n5664 );
not ( n9246 , n4640 );
or ( n9247 , n9245 , n9246 );
or ( n9248 , n4640 , n5664 );
nand ( n9249 , n9247 , n9248 );
nand ( n9250 , n9244 , n9249 );
nor ( n9251 , n9239 , n9250 );
not ( n9252 , n5659 );
not ( n9253 , n4635 );
or ( n9254 , n9252 , n9253 );
or ( n9255 , n4635 , n5659 );
nand ( n9256 , n9254 , n9255 );
not ( n9257 , n5658 );
not ( n9258 , n4634 );
or ( n9259 , n9257 , n9258 );
or ( n9260 , n4634 , n5658 );
nand ( n9261 , n9259 , n9260 );
nand ( n9262 , n9256 , n9261 );
not ( n9263 , n5661 );
not ( n9264 , n4637 );
or ( n9265 , n9263 , n9264 );
or ( n9266 , n4637 , n5661 );
nand ( n9267 , n9265 , n9266 );
not ( n9268 , n5660 );
not ( n9269 , n4636 );
or ( n9270 , n9268 , n9269 );
or ( n9271 , n4636 , n5660 );
nand ( n9272 , n9270 , n9271 );
nand ( n9273 , n9267 , n9272 );
nor ( n9274 , n9262 , n9273 );
not ( n9275 , n5655 );
not ( n9276 , n4631 );
or ( n9277 , n9275 , n9276 );
or ( n9278 , n4631 , n5655 );
nand ( n9279 , n9277 , n9278 );
not ( n9280 , n5654 );
not ( n9281 , n4630 );
or ( n9282 , n9280 , n9281 );
or ( n9283 , n4630 , n5654 );
nand ( n9284 , n9282 , n9283 );
nand ( n9285 , n9279 , n9284 );
not ( n9286 , n5657 );
not ( n9287 , n4633 );
or ( n9288 , n9286 , n9287 );
or ( n9289 , n4633 , n5657 );
nand ( n9290 , n9288 , n9289 );
not ( n9291 , n5656 );
not ( n9292 , n4632 );
or ( n9293 , n9291 , n9292 );
or ( n9294 , n4632 , n5656 );
nand ( n9295 , n9293 , n9294 );
nand ( n9296 , n9290 , n9295 );
nor ( n9297 , n9285 , n9296 );
nand ( n9298 , n9228 , n9251 , n9274 , n9297 );
nor ( n9299 , n9205 , n9298 );
not ( n9300 , n5679 );
not ( n9301 , n4655 );
or ( n9302 , n9300 , n9301 );
or ( n9303 , n4655 , n5679 );
nand ( n9304 , n9302 , n9303 );
not ( n9305 , n5681 );
not ( n9306 , n4657 );
or ( n9307 , n9305 , n9306 );
or ( n9308 , n4657 , n5681 );
nand ( n9309 , n9307 , n9308 );
not ( n9310 , n5678 );
not ( n9311 , n4654 );
or ( n9312 , n9310 , n9311 );
or ( n9313 , n4654 , n5678 );
nand ( n9314 , n9312 , n9313 );
not ( n9315 , n5680 );
not ( n9316 , n4656 );
or ( n9317 , n9315 , n9316 );
or ( n9318 , n4656 , n5680 );
nand ( n9319 , n9317 , n9318 );
nand ( n9320 , n9304 , n9309 , n9314 , n9319 );
not ( n9321 , n9320 );
not ( n9322 , n5675 );
not ( n9323 , n4651 );
or ( n9324 , n9322 , n9323 );
or ( n9325 , n4651 , n5675 );
nand ( n9326 , n9324 , n9325 );
not ( n9327 , n5674 );
not ( n9328 , n4650 );
or ( n9329 , n9327 , n9328 );
or ( n9330 , n4650 , n5674 );
nand ( n9331 , n9329 , n9330 );
nand ( n9332 , n9326 , n9331 );
not ( n9333 , n5677 );
not ( n9334 , n4653 );
or ( n9335 , n9333 , n9334 );
or ( n9336 , n4653 , n5677 );
nand ( n9337 , n9335 , n9336 );
not ( n9338 , n5676 );
not ( n9339 , n4652 );
or ( n9340 , n9338 , n9339 );
or ( n9341 , n4652 , n5676 );
nand ( n9342 , n9340 , n9341 );
nand ( n9343 , n9337 , n9342 );
nor ( n9344 , n9332 , n9343 );
not ( n9345 , n5683 );
not ( n9346 , n4659 );
or ( n9347 , n9345 , n9346 );
or ( n9348 , n4659 , n5683 );
nand ( n9349 , n9347 , n9348 );
not ( n9350 , n5682 );
not ( n9351 , n4658 );
or ( n9352 , n9350 , n9351 );
or ( n9353 , n4658 , n5682 );
nand ( n9354 , n9352 , n9353 );
nand ( n9355 , n9349 , n9354 );
not ( n9356 , n5685 );
not ( n9357 , n4661 );
or ( n9358 , n9356 , n9357 );
or ( n9359 , n4661 , n5685 );
nand ( n9360 , n9358 , n9359 );
not ( n9361 , n5684 );
not ( n9362 , n4660 );
or ( n9363 , n9361 , n9362 );
or ( n9364 , n4660 , n5684 );
nand ( n9365 , n9363 , n9364 );
nand ( n9366 , n9360 , n9365 );
nor ( n9367 , n9355 , n9366 );
not ( n9368 , n5671 );
not ( n9369 , n4647 );
or ( n9370 , n9368 , n9369 );
or ( n9371 , n4647 , n5671 );
nand ( n9372 , n9370 , n9371 );
not ( n9373 , n5670 );
not ( n9374 , n4646 );
or ( n9375 , n9373 , n9374 );
or ( n9376 , n4646 , n5670 );
nand ( n9377 , n9375 , n9376 );
nand ( n9378 , n9372 , n9377 );
not ( n9379 , n5673 );
not ( n9380 , n4649 );
or ( n9381 , n9379 , n9380 );
or ( n9382 , n4649 , n5673 );
nand ( n9383 , n9381 , n9382 );
not ( n9384 , n5672 );
not ( n9385 , n4648 );
or ( n9386 , n9384 , n9385 );
or ( n9387 , n4648 , n5672 );
nand ( n9388 , n9386 , n9387 );
nand ( n9389 , n9383 , n9388 );
nor ( n9390 , n9378 , n9389 );
nand ( n9391 , n9321 , n9344 , n9367 , n9390 );
not ( n9392 , n5695 );
not ( n9393 , n4671 );
or ( n9394 , n9392 , n9393 );
or ( n9395 , n4671 , n5695 );
nand ( n9396 , n9394 , n9395 );
not ( n9397 , n5694 );
not ( n9398 , n4670 );
or ( n9399 , n9397 , n9398 );
or ( n9400 , n4670 , n5694 );
nand ( n9401 , n9399 , n9400 );
nand ( n9402 , n9396 , n9401 );
not ( n9403 , n5697 );
not ( n9404 , n4673 );
or ( n9405 , n9403 , n9404 );
or ( n9406 , n4673 , n5697 );
nand ( n9407 , n9405 , n9406 );
not ( n9408 , n5696 );
not ( n9409 , n4672 );
or ( n9410 , n9408 , n9409 );
or ( n9411 , n4672 , n5696 );
nand ( n9412 , n9410 , n9411 );
nand ( n9413 , n9407 , n9412 );
nor ( n9414 , n9402 , n9413 );
not ( n9415 , n5699 );
not ( n9416 , n4675 );
or ( n9417 , n9415 , n9416 );
or ( n9418 , n4675 , n5699 );
nand ( n9419 , n9417 , n9418 );
not ( n9420 , n5698 );
not ( n9421 , n4674 );
or ( n9422 , n9420 , n9421 );
or ( n9423 , n4674 , n5698 );
nand ( n9424 , n9422 , n9423 );
nand ( n9425 , n9419 , n9424 );
not ( n9426 , n5701 );
not ( n9427 , n4677 );
or ( n9428 , n9426 , n9427 );
or ( n9429 , n4677 , n5701 );
nand ( n9430 , n9428 , n9429 );
not ( n9431 , n5700 );
not ( n9432 , n4676 );
or ( n9433 , n9431 , n9432 );
or ( n9434 , n4676 , n5700 );
nand ( n9435 , n9433 , n9434 );
nand ( n9436 , n9430 , n9435 );
nor ( n9437 , n9425 , n9436 );
not ( n9438 , n5691 );
not ( n9439 , n4667 );
or ( n9440 , n9438 , n9439 );
or ( n9441 , n4667 , n5691 );
nand ( n9442 , n9440 , n9441 );
not ( n9443 , n5690 );
not ( n9444 , n4666 );
or ( n9445 , n9443 , n9444 );
or ( n9446 , n4666 , n5690 );
nand ( n9447 , n9445 , n9446 );
nand ( n9448 , n9442 , n9447 );
not ( n9449 , n5693 );
not ( n9450 , n4669 );
or ( n9451 , n9449 , n9450 );
or ( n9452 , n4669 , n5693 );
nand ( n9453 , n9451 , n9452 );
not ( n9454 , n5692 );
not ( n9455 , n4668 );
or ( n9456 , n9454 , n9455 );
or ( n9457 , n4668 , n5692 );
nand ( n9458 , n9456 , n9457 );
nand ( n9459 , n9453 , n9458 );
nor ( n9460 , n9448 , n9459 );
not ( n9461 , n5687 );
not ( n9462 , n4663 );
or ( n9463 , n9461 , n9462 );
or ( n9464 , n4663 , n5687 );
nand ( n9465 , n9463 , n9464 );
not ( n9466 , n5686 );
not ( n9467 , n4662 );
or ( n9468 , n9466 , n9467 );
or ( n9469 , n4662 , n5686 );
nand ( n9470 , n9468 , n9469 );
nand ( n9471 , n9465 , n9470 );
not ( n9472 , n5689 );
not ( n9473 , n4665 );
or ( n9474 , n9472 , n9473 );
or ( n9475 , n4665 , n5689 );
nand ( n9476 , n9474 , n9475 );
not ( n9477 , n5688 );
not ( n9478 , n4664 );
or ( n9479 , n9477 , n9478 );
or ( n9480 , n4664 , n5688 );
nand ( n9481 , n9479 , n9480 );
nand ( n9482 , n9476 , n9481 );
nor ( n9483 , n9471 , n9482 );
nand ( n9484 , n9414 , n9437 , n9460 , n9483 );
nor ( n9485 , n9391 , n9484 );
not ( n9486 , n5711 );
not ( n9487 , n4687 );
or ( n9488 , n9486 , n9487 );
or ( n9489 , n4687 , n5711 );
nand ( n9490 , n9488 , n9489 );
not ( n9491 , n5710 );
not ( n9492 , n4686 );
or ( n9493 , n9491 , n9492 );
or ( n9494 , n4686 , n5710 );
nand ( n9495 , n9493 , n9494 );
nand ( n9496 , n9490 , n9495 );
not ( n9497 , n5713 );
not ( n9498 , n4689 );
or ( n9499 , n9497 , n9498 );
or ( n9500 , n4689 , n5713 );
nand ( n9501 , n9499 , n9500 );
not ( n9502 , n5712 );
not ( n9503 , n4688 );
or ( n9504 , n9502 , n9503 );
or ( n9505 , n4688 , n5712 );
nand ( n9506 , n9504 , n9505 );
nand ( n9507 , n9501 , n9506 );
nor ( n9508 , n9496 , n9507 );
not ( n9509 , n5716 );
not ( n9510 , n4692 );
or ( n9511 , n9509 , n9510 );
or ( n9512 , n4692 , n5716 );
nand ( n9513 , n9511 , n9512 );
not ( n9514 , n5717 );
not ( n9515 , n4693 );
or ( n9516 , n9514 , n9515 );
or ( n9517 , n4693 , n5717 );
nand ( n9518 , n9516 , n9517 );
not ( n9519 , n5714 );
not ( n9520 , n4690 );
or ( n9521 , n9519 , n9520 );
or ( n9522 , n4690 , n5714 );
nand ( n9523 , n9521 , n9522 );
not ( n9524 , n5715 );
not ( n9525 , n4691 );
or ( n9526 , n9524 , n9525 );
or ( n9527 , n4691 , n5715 );
nand ( n9528 , n9526 , n9527 );
and ( n9529 , n9513 , n9518 , n9523 , n9528 );
not ( n9530 , n5703 );
not ( n9531 , n4679 );
or ( n9532 , n9530 , n9531 );
or ( n9533 , n4679 , n5703 );
nand ( n9534 , n9532 , n9533 );
not ( n9535 , n5702 );
not ( n9536 , n4678 );
or ( n9537 , n9535 , n9536 );
or ( n9538 , n4678 , n5702 );
nand ( n9539 , n9537 , n9538 );
nand ( n9540 , n9534 , n9539 );
not ( n9541 , n5705 );
not ( n9542 , n4681 );
or ( n9543 , n9541 , n9542 );
or ( n9544 , n4681 , n5705 );
nand ( n9545 , n9543 , n9544 );
not ( n9546 , n5704 );
not ( n9547 , n4680 );
or ( n9548 , n9546 , n9547 );
or ( n9549 , n4680 , n5704 );
nand ( n9550 , n9548 , n9549 );
nand ( n9551 , n9545 , n9550 );
nor ( n9552 , n9540 , n9551 );
not ( n9553 , n5709 );
not ( n9554 , n4685 );
or ( n9555 , n9553 , n9554 );
or ( n9556 , n4685 , n5709 );
nand ( n9557 , n9555 , n9556 );
not ( n9558 , n5708 );
not ( n9559 , n4684 );
or ( n9560 , n9558 , n9559 );
or ( n9561 , n4684 , n5708 );
nand ( n9562 , n9560 , n9561 );
nand ( n9563 , n9557 , n9562 );
not ( n9564 , n5707 );
not ( n9565 , n4683 );
or ( n9566 , n9564 , n9565 );
or ( n9567 , n4683 , n5707 );
nand ( n9568 , n9566 , n9567 );
not ( n9569 , n5706 );
not ( n9570 , n4682 );
or ( n9571 , n9569 , n9570 );
or ( n9572 , n4682 , n5706 );
nand ( n9573 , n9571 , n9572 );
nand ( n9574 , n9568 , n9573 );
nor ( n9575 , n9563 , n9574 );
nand ( n9576 , n9508 , n9529 , n9552 , n9575 );
not ( n9577 , n5727 );
not ( n9578 , n4703 );
or ( n9579 , n9577 , n9578 );
or ( n9580 , n4703 , n5727 );
nand ( n9581 , n9579 , n9580 );
not ( n9582 , n5726 );
not ( n9583 , n4702 );
or ( n9584 , n9582 , n9583 );
or ( n9585 , n4702 , n5726 );
nand ( n9586 , n9584 , n9585 );
nand ( n9587 , n9581 , n9586 );
not ( n9588 , n5729 );
not ( n9589 , n4705 );
or ( n9590 , n9588 , n9589 );
or ( n9591 , n4705 , n5729 );
nand ( n9592 , n9590 , n9591 );
not ( n9593 , n5728 );
not ( n9594 , n4704 );
or ( n9595 , n9593 , n9594 );
or ( n9596 , n4704 , n5728 );
nand ( n9597 , n9595 , n9596 );
nand ( n9598 , n9592 , n9597 );
nor ( n9599 , n9587 , n9598 );
not ( n9600 , n5732 );
not ( n9601 , n4708 );
or ( n9602 , n9600 , n9601 );
or ( n9603 , n4708 , n5732 );
nand ( n9604 , n9602 , n9603 );
not ( n9605 , n5733 );
not ( n9606 , n4709 );
or ( n9607 , n9605 , n9606 );
or ( n9608 , n4709 , n5733 );
nand ( n9609 , n9607 , n9608 );
not ( n9610 , n5730 );
not ( n9611 , n4706 );
or ( n9612 , n9610 , n9611 );
or ( n9613 , n4706 , n5730 );
nand ( n9614 , n9612 , n9613 );
not ( n9615 , n5731 );
not ( n9616 , n4707 );
or ( n9617 , n9615 , n9616 );
or ( n9618 , n4707 , n5731 );
nand ( n9619 , n9617 , n9618 );
and ( n9620 , n9604 , n9609 , n9614 , n9619 );
not ( n9621 , n5719 );
not ( n9622 , n4695 );
or ( n9623 , n9621 , n9622 );
or ( n9624 , n4695 , n5719 );
nand ( n9625 , n9623 , n9624 );
not ( n9626 , n5718 );
not ( n9627 , n4694 );
or ( n9628 , n9626 , n9627 );
or ( n9629 , n4694 , n5718 );
nand ( n9630 , n9628 , n9629 );
nand ( n9631 , n9625 , n9630 );
not ( n9632 , n5721 );
not ( n9633 , n4697 );
or ( n9634 , n9632 , n9633 );
or ( n9635 , n4697 , n5721 );
nand ( n9636 , n9634 , n9635 );
not ( n9637 , n5720 );
not ( n9638 , n4696 );
or ( n9639 , n9637 , n9638 );
or ( n9640 , n4696 , n5720 );
nand ( n9641 , n9639 , n9640 );
nand ( n9642 , n9636 , n9641 );
nor ( n9643 , n9631 , n9642 );
not ( n9644 , n5725 );
not ( n9645 , n4701 );
or ( n9646 , n9644 , n9645 );
or ( n9647 , n4701 , n5725 );
nand ( n9648 , n9646 , n9647 );
not ( n9649 , n5724 );
not ( n9650 , n4700 );
or ( n9651 , n9649 , n9650 );
or ( n9652 , n4700 , n5724 );
nand ( n9653 , n9651 , n9652 );
nand ( n9654 , n9648 , n9653 );
not ( n9655 , n5723 );
not ( n9656 , n4699 );
or ( n9657 , n9655 , n9656 );
or ( n9658 , n4699 , n5723 );
nand ( n9659 , n9657 , n9658 );
not ( n9660 , n5722 );
not ( n9661 , n4698 );
or ( n9662 , n9660 , n9661 );
or ( n9663 , n4698 , n5722 );
nand ( n9664 , n9662 , n9663 );
nand ( n9665 , n9659 , n9664 );
nor ( n9666 , n9654 , n9665 );
nand ( n9667 , n9599 , n9620 , n9643 , n9666 );
nor ( n9668 , n9576 , n9667 );
not ( n9669 , n5747 );
not ( n9670 , n4723 );
or ( n9671 , n9669 , n9670 );
or ( n9672 , n4723 , n5747 );
nand ( n9673 , n9671 , n9672 );
not ( n9674 , n5746 );
not ( n9675 , n4722 );
or ( n9676 , n9674 , n9675 );
or ( n9677 , n4722 , n5746 );
nand ( n9678 , n9676 , n9677 );
nand ( n9679 , n9673 , n9678 );
not ( n9680 , n5749 );
not ( n9681 , n4725 );
or ( n9682 , n9680 , n9681 );
or ( n9683 , n4725 , n5749 );
nand ( n9684 , n9682 , n9683 );
not ( n9685 , n5748 );
not ( n9686 , n4724 );
or ( n9687 , n9685 , n9686 );
or ( n9688 , n4724 , n5748 );
nand ( n9689 , n9687 , n9688 );
nand ( n9690 , n9684 , n9689 );
nor ( n9691 , n9679 , n9690 );
not ( n9692 , n5743 );
not ( n9693 , n4719 );
or ( n9694 , n9692 , n9693 );
or ( n9695 , n4719 , n5743 );
nand ( n9696 , n9694 , n9695 );
not ( n9697 , n5742 );
not ( n9698 , n4718 );
or ( n9699 , n9697 , n9698 );
or ( n9700 , n4718 , n5742 );
nand ( n9701 , n9699 , n9700 );
nand ( n9702 , n9696 , n9701 );
not ( n9703 , n5745 );
not ( n9704 , n4721 );
or ( n9705 , n9703 , n9704 );
or ( n9706 , n4721 , n5745 );
nand ( n9707 , n9705 , n9706 );
not ( n9708 , n5744 );
not ( n9709 , n4720 );
or ( n9710 , n9708 , n9709 );
or ( n9711 , n4720 , n5744 );
nand ( n9712 , n9710 , n9711 );
nand ( n9713 , n9707 , n9712 );
nor ( n9714 , n9702 , n9713 );
not ( n9715 , n5736 );
not ( n9716 , n4712 );
or ( n9717 , n9715 , n9716 );
or ( n9718 , n4712 , n5736 );
nand ( n9719 , n9717 , n9718 );
not ( n9720 , n5737 );
not ( n9721 , n4713 );
or ( n9722 , n9720 , n9721 );
or ( n9723 , n4713 , n5737 );
nand ( n9724 , n9722 , n9723 );
not ( n9725 , n5734 );
not ( n9726 , n4710 );
or ( n9727 , n9725 , n9726 );
or ( n9728 , n4710 , n5734 );
nand ( n9729 , n9727 , n9728 );
not ( n9730 , n5735 );
not ( n9731 , n4711 );
or ( n9732 , n9730 , n9731 );
or ( n9733 , n4711 , n5735 );
nand ( n9734 , n9732 , n9733 );
nand ( n9735 , n9719 , n9724 , n9729 , n9734 );
not ( n9736 , n9735 );
not ( n9737 , n5739 );
not ( n9738 , n4715 );
or ( n9739 , n9737 , n9738 );
or ( n9740 , n4715 , n5739 );
nand ( n9741 , n9739 , n9740 );
not ( n9742 , n5738 );
not ( n9743 , n4714 );
or ( n9744 , n9742 , n9743 );
or ( n9745 , n4714 , n5738 );
nand ( n9746 , n9744 , n9745 );
nand ( n9747 , n9741 , n9746 );
not ( n9748 , n5741 );
not ( n9749 , n4717 );
or ( n9750 , n9748 , n9749 );
or ( n9751 , n4717 , n5741 );
nand ( n9752 , n9750 , n9751 );
not ( n9753 , n5740 );
not ( n9754 , n4716 );
or ( n9755 , n9753 , n9754 );
or ( n9756 , n4716 , n5740 );
nand ( n9757 , n9755 , n9756 );
nand ( n9758 , n9752 , n9757 );
nor ( n9759 , n9747 , n9758 );
nand ( n9760 , n9691 , n9714 , n9736 , n9759 );
not ( n9761 , n5763 );
not ( n9762 , n4739 );
or ( n9763 , n9761 , n9762 );
or ( n9764 , n4739 , n5763 );
nand ( n9765 , n9763 , n9764 );
not ( n9766 , n5762 );
not ( n9767 , n4738 );
or ( n9768 , n9766 , n9767 );
or ( n9769 , n4738 , n5762 );
nand ( n9770 , n9768 , n9769 );
nand ( n9771 , n9765 , n9770 );
not ( n9772 , n5765 );
not ( n9773 , n4741 );
or ( n9774 , n9772 , n9773 );
or ( n9775 , n4741 , n5765 );
nand ( n9776 , n9774 , n9775 );
not ( n9777 , n5764 );
not ( n9778 , n4740 );
or ( n9779 , n9777 , n9778 );
or ( n9780 , n4740 , n5764 );
nand ( n9781 , n9779 , n9780 );
nand ( n9782 , n9776 , n9781 );
nor ( n9783 , n9771 , n9782 );
not ( n9784 , n5752 );
not ( n9785 , n4728 );
or ( n9786 , n9784 , n9785 );
or ( n9787 , n4728 , n5752 );
nand ( n9788 , n9786 , n9787 );
not ( n9789 , n5753 );
not ( n9790 , n4729 );
or ( n9791 , n9789 , n9790 );
or ( n9792 , n4729 , n5753 );
nand ( n9793 , n9791 , n9792 );
not ( n9794 , n5750 );
not ( n9795 , n4726 );
or ( n9796 , n9794 , n9795 );
or ( n9797 , n4726 , n5750 );
nand ( n9798 , n9796 , n9797 );
not ( n9799 , n5751 );
not ( n9800 , n4727 );
or ( n9801 , n9799 , n9800 );
or ( n9802 , n4727 , n5751 );
nand ( n9803 , n9801 , n9802 );
nand ( n9804 , n9788 , n9793 , n9798 , n9803 );
not ( n9805 , n9804 );
not ( n9806 , n5755 );
not ( n9807 , n4731 );
or ( n9808 , n9806 , n9807 );
or ( n9809 , n4731 , n5755 );
nand ( n9810 , n9808 , n9809 );
not ( n9811 , n5754 );
not ( n9812 , n4730 );
or ( n9813 , n9811 , n9812 );
or ( n9814 , n4730 , n5754 );
nand ( n9815 , n9813 , n9814 );
nand ( n9816 , n9810 , n9815 );
not ( n9817 , n5757 );
not ( n9818 , n4733 );
or ( n9819 , n9817 , n9818 );
or ( n9820 , n4733 , n5757 );
nand ( n9821 , n9819 , n9820 );
not ( n9822 , n5756 );
not ( n9823 , n4732 );
or ( n9824 , n9822 , n9823 );
or ( n9825 , n4732 , n5756 );
nand ( n9826 , n9824 , n9825 );
nand ( n9827 , n9821 , n9826 );
nor ( n9828 , n9816 , n9827 );
not ( n9829 , n5760 );
not ( n9830 , n4736 );
or ( n9831 , n9829 , n9830 );
or ( n9832 , n4736 , n5760 );
nand ( n9833 , n9831 , n9832 );
not ( n9834 , n5761 );
not ( n9835 , n4737 );
or ( n9836 , n9834 , n9835 );
or ( n9837 , n4737 , n5761 );
nand ( n9838 , n9836 , n9837 );
not ( n9839 , n4734 );
not ( n9840 , n5758 );
or ( n9841 , n9839 , n9840 );
or ( n9842 , n5758 , n4734 );
nand ( n9843 , n9841 , n9842 );
not ( n9844 , n4735 );
and ( n9845 , n5759 , n9844 );
not ( n9846 , n5759 );
and ( n9847 , n9846 , n4735 );
nor ( n9848 , n9845 , n9847 );
nand ( n9849 , n9833 , n9838 , n9843 , n9848 );
not ( n9850 , n9849 );
nand ( n9851 , n9783 , n9805 , n9828 , n9850 );
nor ( n9852 , n9760 , n9851 );
nand ( n9853 , n9299 , n9485 , n9668 , n9852 );
not ( n9854 , n5771 );
not ( n9855 , n4747 );
or ( n9856 , n9854 , n9855 );
or ( n9857 , n4747 , n5771 );
nand ( n9858 , n9856 , n9857 );
not ( n9859 , n5770 );
not ( n9860 , n4746 );
or ( n9861 , n9859 , n9860 );
or ( n9862 , n4746 , n5770 );
nand ( n9863 , n9861 , n9862 );
nand ( n9864 , n9858 , n9863 );
not ( n9865 , n5773 );
not ( n9866 , n4749 );
or ( n9867 , n9865 , n9866 );
or ( n9868 , n4749 , n5773 );
nand ( n9869 , n9867 , n9868 );
not ( n9870 , n5772 );
not ( n9871 , n4748 );
or ( n9872 , n9870 , n9871 );
or ( n9873 , n4748 , n5772 );
nand ( n9874 , n9872 , n9873 );
nand ( n9875 , n9869 , n9874 );
nor ( n9876 , n9864 , n9875 );
not ( n9877 , n5779 );
not ( n9878 , n4755 );
or ( n9879 , n9877 , n9878 );
or ( n9880 , n4755 , n5779 );
nand ( n9881 , n9879 , n9880 );
not ( n9882 , n5778 );
not ( n9883 , n4754 );
or ( n9884 , n9882 , n9883 );
or ( n9885 , n4754 , n5778 );
nand ( n9886 , n9884 , n9885 );
nand ( n9887 , n9881 , n9886 );
not ( n9888 , n5781 );
not ( n9889 , n4757 );
or ( n9890 , n9888 , n9889 );
or ( n9891 , n4757 , n5781 );
nand ( n9892 , n9890 , n9891 );
not ( n9893 , n5780 );
not ( n9894 , n4756 );
or ( n9895 , n9893 , n9894 );
or ( n9896 , n4756 , n5780 );
nand ( n9897 , n9895 , n9896 );
nand ( n9898 , n9892 , n9897 );
nor ( n9899 , n9887 , n9898 );
not ( n9900 , n5767 );
not ( n9901 , n4743 );
or ( n9902 , n9900 , n9901 );
or ( n9903 , n4743 , n5767 );
nand ( n9904 , n9902 , n9903 );
not ( n9905 , n5766 );
not ( n9906 , n4742 );
or ( n9907 , n9905 , n9906 );
or ( n9908 , n4742 , n5766 );
nand ( n9909 , n9907 , n9908 );
nand ( n9910 , n9904 , n9909 );
not ( n9911 , n5769 );
not ( n9912 , n4745 );
or ( n9913 , n9911 , n9912 );
or ( n9914 , n4745 , n5769 );
nand ( n9915 , n9913 , n9914 );
not ( n9916 , n5768 );
not ( n9917 , n4744 );
or ( n9918 , n9916 , n9917 );
or ( n9919 , n4744 , n5768 );
nand ( n9920 , n9918 , n9919 );
nand ( n9921 , n9915 , n9920 );
nor ( n9922 , n9910 , n9921 );
not ( n9923 , n5775 );
not ( n9924 , n4751 );
or ( n9925 , n9923 , n9924 );
or ( n9926 , n4751 , n5775 );
nand ( n9927 , n9925 , n9926 );
not ( n9928 , n5777 );
not ( n9929 , n4753 );
or ( n9930 , n9928 , n9929 );
or ( n9931 , n4753 , n5777 );
nand ( n9932 , n9930 , n9931 );
not ( n9933 , n5774 );
not ( n9934 , n4750 );
or ( n9935 , n9933 , n9934 );
or ( n9936 , n4750 , n5774 );
nand ( n9937 , n9935 , n9936 );
not ( n9938 , n5776 );
not ( n9939 , n4752 );
or ( n9940 , n9938 , n9939 );
or ( n9941 , n4752 , n5776 );
nand ( n9942 , n9940 , n9941 );
and ( n9943 , n9927 , n9932 , n9937 , n9942 );
nand ( n9944 , n9876 , n9899 , n9922 , n9943 );
not ( n9945 , n5795 );
not ( n9946 , n4771 );
or ( n9947 , n9945 , n9946 );
or ( n9948 , n4771 , n5795 );
nand ( n9949 , n9947 , n9948 );
not ( n9950 , n5794 );
not ( n9951 , n4770 );
or ( n9952 , n9950 , n9951 );
or ( n9953 , n4770 , n5794 );
nand ( n9954 , n9952 , n9953 );
nand ( n9955 , n9949 , n9954 );
not ( n9956 , n5797 );
not ( n9957 , n4773 );
or ( n9958 , n9956 , n9957 );
or ( n9959 , n4773 , n5797 );
nand ( n9960 , n9958 , n9959 );
not ( n9961 , n5796 );
not ( n9962 , n4772 );
or ( n9963 , n9961 , n9962 );
or ( n9964 , n4772 , n5796 );
nand ( n9965 , n9963 , n9964 );
nand ( n9966 , n9960 , n9965 );
nor ( n9967 , n9955 , n9966 );
not ( n9968 , n5791 );
not ( n9969 , n4767 );
or ( n9970 , n9968 , n9969 );
or ( n9971 , n4767 , n5791 );
nand ( n9972 , n9970 , n9971 );
not ( n9973 , n5790 );
not ( n9974 , n4766 );
or ( n9975 , n9973 , n9974 );
or ( n9976 , n4766 , n5790 );
nand ( n9977 , n9975 , n9976 );
nand ( n9978 , n9972 , n9977 );
not ( n9979 , n5793 );
not ( n9980 , n4769 );
or ( n9981 , n9979 , n9980 );
or ( n9982 , n4769 , n5793 );
nand ( n9983 , n9981 , n9982 );
not ( n9984 , n5792 );
not ( n9985 , n4768 );
or ( n9986 , n9984 , n9985 );
or ( n9987 , n4768 , n5792 );
nand ( n9988 , n9986 , n9987 );
nand ( n9989 , n9983 , n9988 );
nor ( n9990 , n9978 , n9989 );
not ( n9991 , n5787 );
not ( n9992 , n4763 );
or ( n9993 , n9991 , n9992 );
or ( n9994 , n4763 , n5787 );
nand ( n9995 , n9993 , n9994 );
not ( n9996 , n5786 );
not ( n9997 , n4762 );
or ( n9998 , n9996 , n9997 );
or ( n9999 , n4762 , n5786 );
nand ( n10000 , n9998 , n9999 );
nand ( n10001 , n9995 , n10000 );
not ( n10002 , n5789 );
not ( n10003 , n4765 );
or ( n10004 , n10002 , n10003 );
or ( n10005 , n4765 , n5789 );
nand ( n10006 , n10004 , n10005 );
not ( n10007 , n5788 );
not ( n10008 , n4764 );
or ( n10009 , n10007 , n10008 );
or ( n10010 , n4764 , n5788 );
nand ( n10011 , n10009 , n10010 );
nand ( n10012 , n10006 , n10011 );
nor ( n10013 , n10001 , n10012 );
not ( n10014 , n5783 );
not ( n10015 , n4759 );
or ( n10016 , n10014 , n10015 );
or ( n10017 , n4759 , n5783 );
nand ( n10018 , n10016 , n10017 );
not ( n10019 , n5782 );
not ( n10020 , n4758 );
or ( n10021 , n10019 , n10020 );
or ( n10022 , n4758 , n5782 );
nand ( n10023 , n10021 , n10022 );
nand ( n10024 , n10018 , n10023 );
not ( n10025 , n5785 );
not ( n10026 , n4761 );
or ( n10027 , n10025 , n10026 );
or ( n10028 , n4761 , n5785 );
nand ( n10029 , n10027 , n10028 );
not ( n10030 , n5784 );
not ( n10031 , n4760 );
or ( n10032 , n10030 , n10031 );
or ( n10033 , n4760 , n5784 );
nand ( n10034 , n10032 , n10033 );
nand ( n10035 , n10029 , n10034 );
nor ( n10036 , n10024 , n10035 );
nand ( n10037 , n9967 , n9990 , n10013 , n10036 );
nor ( n10038 , n9944 , n10037 );
not ( n10039 , n5803 );
not ( n10040 , n4779 );
or ( n10041 , n10039 , n10040 );
or ( n10042 , n4779 , n5803 );
nand ( n10043 , n10041 , n10042 );
not ( n10044 , n5805 );
not ( n10045 , n4781 );
or ( n10046 , n10044 , n10045 );
or ( n10047 , n4781 , n5805 );
nand ( n10048 , n10046 , n10047 );
not ( n10049 , n5802 );
not ( n10050 , n4778 );
or ( n10051 , n10049 , n10050 );
or ( n10052 , n4778 , n5802 );
nand ( n10053 , n10051 , n10052 );
not ( n10054 , n5804 );
not ( n10055 , n4780 );
or ( n10056 , n10054 , n10055 );
or ( n10057 , n4780 , n5804 );
nand ( n10058 , n10056 , n10057 );
nand ( n10059 , n10043 , n10048 , n10053 , n10058 );
not ( n10060 , n5798 );
not ( n10061 , n4774 );
or ( n10062 , n10060 , n10061 );
or ( n10063 , n4774 , n5798 );
nand ( n10064 , n10062 , n10063 );
not ( n10065 , n5799 );
not ( n10066 , n4775 );
or ( n10067 , n10065 , n10066 );
or ( n10068 , n4775 , n5799 );
nand ( n10069 , n10067 , n10068 );
not ( n10070 , n5800 );
not ( n10071 , n4776 );
or ( n10072 , n10070 , n10071 );
or ( n10073 , n4776 , n5800 );
nand ( n10074 , n10072 , n10073 );
not ( n10075 , n5801 );
not ( n10076 , n4777 );
or ( n10077 , n10075 , n10076 );
or ( n10078 , n4777 , n5801 );
nand ( n10079 , n10077 , n10078 );
nand ( n10080 , n10064 , n10069 , n10074 , n10079 );
nor ( n10081 , n10059 , n10080 );
not ( n10082 , n5808 );
not ( n10083 , n4784 );
or ( n10084 , n10082 , n10083 );
or ( n10085 , n4784 , n5808 );
nand ( n10086 , n10084 , n10085 );
not ( n10087 , n5809 );
not ( n10088 , n4785 );
or ( n10089 , n10087 , n10088 );
or ( n10090 , n4785 , n5809 );
nand ( n10091 , n10089 , n10090 );
not ( n10092 , n5806 );
not ( n10093 , n4782 );
or ( n10094 , n10092 , n10093 );
or ( n10095 , n4782 , n5806 );
nand ( n10096 , n10094 , n10095 );
not ( n10097 , n5807 );
not ( n10098 , n4783 );
or ( n10099 , n10097 , n10098 );
or ( n10100 , n4783 , n5807 );
nand ( n10101 , n10099 , n10100 );
nand ( n10102 , n10086 , n10091 , n10096 , n10101 );
not ( n10103 , n4787 );
not ( n10104 , n5811 );
or ( n10105 , n10103 , n10104 );
or ( n10106 , n5811 , n4787 );
nand ( n10107 , n10105 , n10106 );
not ( n10108 , n4786 );
not ( n10109 , n5810 );
or ( n10110 , n10108 , n10109 );
or ( n10111 , n5810 , n4786 );
nand ( n10112 , n10110 , n10111 );
not ( n10113 , n4789 );
not ( n10114 , n5813 );
or ( n10115 , n10113 , n10114 );
or ( n10116 , n5813 , n4789 );
nand ( n10117 , n10115 , n10116 );
not ( n10118 , n4788 );
not ( n10119 , n5812 );
or ( n10120 , n10118 , n10119 );
or ( n10121 , n5812 , n4788 );
nand ( n10122 , n10120 , n10121 );
nand ( n10123 , n10107 , n10112 , n10117 , n10122 );
nor ( n10124 , n10102 , n10123 );
nand ( n10125 , n10081 , n10124 );
not ( n10126 , n5828 );
not ( n10127 , n4804 );
or ( n10128 , n10126 , n10127 );
or ( n10129 , n4804 , n5828 );
nand ( n10130 , n10128 , n10129 );
not ( n10131 , n5829 );
not ( n10132 , n4805 );
or ( n10133 , n10131 , n10132 );
or ( n10134 , n4805 , n5829 );
nand ( n10135 , n10133 , n10134 );
not ( n10136 , n5826 );
not ( n10137 , n4802 );
or ( n10138 , n10136 , n10137 );
or ( n10139 , n4802 , n5826 );
nand ( n10140 , n10138 , n10139 );
not ( n10141 , n5827 );
not ( n10142 , n4803 );
or ( n10143 , n10141 , n10142 );
or ( n10144 , n4803 , n5827 );
nand ( n10145 , n10143 , n10144 );
nand ( n10146 , n10130 , n10135 , n10140 , n10145 );
not ( n10147 , n10146 );
not ( n10148 , n5823 );
not ( n10149 , n4799 );
or ( n10150 , n10148 , n10149 );
or ( n10151 , n4799 , n5823 );
nand ( n10152 , n10150 , n10151 );
not ( n10153 , n5822 );
not ( n10154 , n4798 );
or ( n10155 , n10153 , n10154 );
or ( n10156 , n4798 , n5822 );
nand ( n10157 , n10155 , n10156 );
nand ( n10158 , n10152 , n10157 );
not ( n10159 , n5825 );
not ( n10160 , n4801 );
or ( n10161 , n10159 , n10160 );
or ( n10162 , n4801 , n5825 );
nand ( n10163 , n10161 , n10162 );
not ( n10164 , n5824 );
not ( n10165 , n4800 );
or ( n10166 , n10164 , n10165 );
or ( n10167 , n4800 , n5824 );
nand ( n10168 , n10166 , n10167 );
nand ( n10169 , n10163 , n10168 );
nor ( n10170 , n10158 , n10169 );
not ( n10171 , n5819 );
not ( n10172 , n4795 );
or ( n10173 , n10171 , n10172 );
or ( n10174 , n4795 , n5819 );
nand ( n10175 , n10173 , n10174 );
not ( n10176 , n5818 );
not ( n10177 , n4794 );
or ( n10178 , n10176 , n10177 );
or ( n10179 , n4794 , n5818 );
nand ( n10180 , n10178 , n10179 );
nand ( n10181 , n10175 , n10180 );
not ( n10182 , n5821 );
not ( n10183 , n4797 );
or ( n10184 , n10182 , n10183 );
or ( n10185 , n4797 , n5821 );
nand ( n10186 , n10184 , n10185 );
not ( n10187 , n5820 );
not ( n10188 , n4796 );
or ( n10189 , n10187 , n10188 );
or ( n10190 , n4796 , n5820 );
nand ( n10191 , n10189 , n10190 );
nand ( n10192 , n10186 , n10191 );
nor ( n10193 , n10181 , n10192 );
not ( n10194 , n5817 );
not ( n10195 , n4793 );
or ( n10196 , n10194 , n10195 );
or ( n10197 , n4793 , n5817 );
nand ( n10198 , n10196 , n10197 );
not ( n10199 , n5816 );
not ( n10200 , n4792 );
or ( n10201 , n10199 , n10200 );
or ( n10202 , n4792 , n5816 );
nand ( n10203 , n10201 , n10202 );
nand ( n10204 , n10198 , n10203 );
not ( n10205 , n5815 );
not ( n10206 , n4791 );
or ( n10207 , n10205 , n10206 );
or ( n10208 , n4791 , n5815 );
nand ( n10209 , n10207 , n10208 );
not ( n10210 , n5814 );
not ( n10211 , n4790 );
or ( n10212 , n10210 , n10211 );
or ( n10213 , n4790 , n5814 );
nand ( n10214 , n10212 , n10213 );
nand ( n10215 , n10209 , n10214 );
nor ( n10216 , n10204 , n10215 );
nand ( n10217 , n10147 , n10170 , n10193 , n10216 );
nor ( n10218 , n10125 , n10217 );
not ( n10219 , n5859 );
not ( n10220 , n4835 );
or ( n10221 , n10219 , n10220 );
or ( n10222 , n4835 , n5859 );
nand ( n10223 , n10221 , n10222 );
not ( n10224 , n5858 );
not ( n10225 , n4834 );
or ( n10226 , n10224 , n10225 );
or ( n10227 , n4834 , n5858 );
nand ( n10228 , n10226 , n10227 );
nand ( n10229 , n10223 , n10228 );
not ( n10230 , n5861 );
not ( n10231 , n4837 );
or ( n10232 , n10230 , n10231 );
or ( n10233 , n4837 , n5861 );
nand ( n10234 , n10232 , n10233 );
not ( n10235 , n5860 );
not ( n10236 , n4836 );
or ( n10237 , n10235 , n10236 );
or ( n10238 , n4836 , n5860 );
nand ( n10239 , n10237 , n10238 );
nand ( n10240 , n10234 , n10239 );
nor ( n10241 , n10229 , n10240 );
not ( n10242 , n5855 );
not ( n10243 , n4831 );
or ( n10244 , n10242 , n10243 );
or ( n10245 , n4831 , n5855 );
nand ( n10246 , n10244 , n10245 );
not ( n10247 , n5854 );
not ( n10248 , n4830 );
or ( n10249 , n10247 , n10248 );
or ( n10250 , n4830 , n5854 );
nand ( n10251 , n10249 , n10250 );
nand ( n10252 , n10246 , n10251 );
not ( n10253 , n5857 );
not ( n10254 , n4833 );
or ( n10255 , n10253 , n10254 );
or ( n10256 , n4833 , n5857 );
nand ( n10257 , n10255 , n10256 );
not ( n10258 , n5856 );
not ( n10259 , n4832 );
or ( n10260 , n10258 , n10259 );
or ( n10261 , n4832 , n5856 );
nand ( n10262 , n10260 , n10261 );
nand ( n10263 , n10257 , n10262 );
nor ( n10264 , n10252 , n10263 );
not ( n10265 , n5848 );
not ( n10266 , n4824 );
or ( n10267 , n10265 , n10266 );
or ( n10268 , n4824 , n5848 );
nand ( n10269 , n10267 , n10268 );
not ( n10270 , n5849 );
not ( n10271 , n4825 );
or ( n10272 , n10270 , n10271 );
or ( n10273 , n4825 , n5849 );
nand ( n10274 , n10272 , n10273 );
not ( n10275 , n5846 );
not ( n10276 , n4822 );
or ( n10277 , n10275 , n10276 );
or ( n10278 , n4822 , n5846 );
nand ( n10279 , n10277 , n10278 );
not ( n10280 , n5847 );
not ( n10281 , n4823 );
or ( n10282 , n10280 , n10281 );
or ( n10283 , n4823 , n5847 );
nand ( n10284 , n10282 , n10283 );
nand ( n10285 , n10269 , n10274 , n10279 , n10284 );
not ( n10286 , n10285 );
not ( n10287 , n5853 );
not ( n10288 , n4829 );
or ( n10289 , n10287 , n10288 );
or ( n10290 , n4829 , n5853 );
nand ( n10291 , n10289 , n10290 );
not ( n10292 , n5852 );
not ( n10293 , n4828 );
or ( n10294 , n10292 , n10293 );
or ( n10295 , n4828 , n5852 );
nand ( n10296 , n10294 , n10295 );
nand ( n10297 , n10291 , n10296 );
not ( n10298 , n5851 );
not ( n10299 , n4827 );
or ( n10300 , n10298 , n10299 );
or ( n10301 , n4827 , n5851 );
nand ( n10302 , n10300 , n10301 );
not ( n10303 , n5850 );
not ( n10304 , n4826 );
or ( n10305 , n10303 , n10304 );
or ( n10306 , n4826 , n5850 );
nand ( n10307 , n10305 , n10306 );
nand ( n10308 , n10302 , n10307 );
nor ( n10309 , n10297 , n10308 );
nand ( n10310 , n10241 , n10264 , n10286 , n10309 );
not ( n10311 , n5843 );
not ( n10312 , n4819 );
or ( n10313 , n10311 , n10312 );
or ( n10314 , n4819 , n5843 );
nand ( n10315 , n10313 , n10314 );
not ( n10316 , n5842 );
not ( n10317 , n4818 );
or ( n10318 , n10316 , n10317 );
or ( n10319 , n4818 , n5842 );
nand ( n10320 , n10318 , n10319 );
nand ( n10321 , n10315 , n10320 );
not ( n10322 , n5845 );
not ( n10323 , n4821 );
or ( n10324 , n10322 , n10323 );
or ( n10325 , n4821 , n5845 );
nand ( n10326 , n10324 , n10325 );
not ( n10327 , n5844 );
not ( n10328 , n4820 );
or ( n10329 , n10327 , n10328 );
or ( n10330 , n4820 , n5844 );
nand ( n10331 , n10329 , n10330 );
nand ( n10332 , n10326 , n10331 );
nor ( n10333 , n10321 , n10332 );
not ( n10334 , n5839 );
not ( n10335 , n4815 );
or ( n10336 , n10334 , n10335 );
or ( n10337 , n4815 , n5839 );
nand ( n10338 , n10336 , n10337 );
not ( n10339 , n5838 );
not ( n10340 , n4814 );
or ( n10341 , n10339 , n10340 );
or ( n10342 , n4814 , n5838 );
nand ( n10343 , n10341 , n10342 );
nand ( n10344 , n10338 , n10343 );
not ( n10345 , n5841 );
not ( n10346 , n4817 );
or ( n10347 , n10345 , n10346 );
or ( n10348 , n4817 , n5841 );
nand ( n10349 , n10347 , n10348 );
not ( n10350 , n5840 );
not ( n10351 , n4816 );
or ( n10352 , n10350 , n10351 );
or ( n10353 , n4816 , n5840 );
nand ( n10354 , n10352 , n10353 );
nand ( n10355 , n10349 , n10354 );
nor ( n10356 , n10344 , n10355 );
not ( n10357 , n5832 );
not ( n10358 , n4808 );
or ( n10359 , n10357 , n10358 );
or ( n10360 , n4808 , n5832 );
nand ( n10361 , n10359 , n10360 );
not ( n10362 , n5833 );
not ( n10363 , n4809 );
or ( n10364 , n10362 , n10363 );
or ( n10365 , n4809 , n5833 );
nand ( n10366 , n10364 , n10365 );
not ( n10367 , n5830 );
not ( n10368 , n4806 );
or ( n10369 , n10367 , n10368 );
or ( n10370 , n4806 , n5830 );
nand ( n10371 , n10369 , n10370 );
not ( n10372 , n5831 );
not ( n10373 , n4807 );
or ( n10374 , n10372 , n10373 );
or ( n10375 , n4807 , n5831 );
nand ( n10376 , n10374 , n10375 );
nand ( n10377 , n10361 , n10366 , n10371 , n10376 );
not ( n10378 , n10377 );
not ( n10379 , n5836 );
not ( n10380 , n4812 );
or ( n10381 , n10379 , n10380 );
or ( n10382 , n4812 , n5836 );
nand ( n10383 , n10381 , n10382 );
not ( n10384 , n5837 );
not ( n10385 , n4813 );
or ( n10386 , n10384 , n10385 );
or ( n10387 , n4813 , n5837 );
nand ( n10388 , n10386 , n10387 );
not ( n10389 , n4810 );
not ( n10390 , n5834 );
or ( n10391 , n10389 , n10390 );
or ( n10392 , n5834 , n4810 );
nand ( n10393 , n10391 , n10392 );
not ( n10394 , n4811 );
and ( n10395 , n5835 , n10394 );
not ( n10396 , n5835 );
and ( n10397 , n10396 , n4811 );
nor ( n10398 , n10395 , n10397 );
nand ( n10399 , n10383 , n10388 , n10393 , n10398 );
not ( n10400 , n10399 );
nand ( n10401 , n10333 , n10356 , n10378 , n10400 );
nor ( n10402 , n10310 , n10401 );
not ( n10403 , n5875 );
not ( n10404 , n4851 );
or ( n10405 , n10403 , n10404 );
or ( n10406 , n4851 , n5875 );
nand ( n10407 , n10405 , n10406 );
not ( n10408 , n5874 );
not ( n10409 , n4850 );
or ( n10410 , n10408 , n10409 );
or ( n10411 , n4850 , n5874 );
nand ( n10412 , n10410 , n10411 );
nand ( n10413 , n10407 , n10412 );
not ( n10414 , n5877 );
not ( n10415 , n4853 );
or ( n10416 , n10414 , n10415 );
or ( n10417 , n4853 , n5877 );
nand ( n10418 , n10416 , n10417 );
not ( n10419 , n5876 );
not ( n10420 , n4852 );
or ( n10421 , n10419 , n10420 );
or ( n10422 , n4852 , n5876 );
nand ( n10423 , n10421 , n10422 );
nand ( n10424 , n10418 , n10423 );
nor ( n10425 , n10413 , n10424 );
not ( n10426 , n5864 );
not ( n10427 , n4840 );
or ( n10428 , n10426 , n10427 );
or ( n10429 , n4840 , n5864 );
nand ( n10430 , n10428 , n10429 );
not ( n10431 , n5865 );
not ( n10432 , n4841 );
or ( n10433 , n10431 , n10432 );
or ( n10434 , n4841 , n5865 );
nand ( n10435 , n10433 , n10434 );
nand ( n10436 , n10430 , n10435 );
not ( n10437 , n5863 );
not ( n10438 , n4839 );
or ( n10439 , n10437 , n10438 );
or ( n10440 , n4839 , n5863 );
nand ( n10441 , n10439 , n10440 );
not ( n10442 , n5862 );
not ( n10443 , n4838 );
or ( n10444 , n10442 , n10443 );
or ( n10445 , n4838 , n5862 );
nand ( n10446 , n10444 , n10445 );
nand ( n10447 , n10441 , n10446 );
nor ( n10448 , n10436 , n10447 );
not ( n10449 , n5867 );
not ( n10450 , n4843 );
or ( n10451 , n10449 , n10450 );
or ( n10452 , n4843 , n5867 );
nand ( n10453 , n10451 , n10452 );
not ( n10454 , n5866 );
not ( n10455 , n4842 );
or ( n10456 , n10454 , n10455 );
or ( n10457 , n4842 , n5866 );
nand ( n10458 , n10456 , n10457 );
nand ( n10459 , n10453 , n10458 );
not ( n10460 , n5869 );
not ( n10461 , n4845 );
or ( n10462 , n10460 , n10461 );
or ( n10463 , n4845 , n5869 );
nand ( n10464 , n10462 , n10463 );
not ( n10465 , n5868 );
not ( n10466 , n4844 );
or ( n10467 , n10465 , n10466 );
or ( n10468 , n4844 , n5868 );
nand ( n10469 , n10467 , n10468 );
nand ( n10470 , n10464 , n10469 );
nor ( n10471 , n10459 , n10470 );
not ( n10472 , n5870 );
not ( n10473 , n4846 );
or ( n10474 , n10472 , n10473 );
or ( n10475 , n4846 , n5870 );
nand ( n10476 , n10474 , n10475 );
not ( n10477 , n5871 );
not ( n10478 , n4847 );
or ( n10479 , n10477 , n10478 );
or ( n10480 , n4847 , n5871 );
nand ( n10481 , n10479 , n10480 );
not ( n10482 , n4848 );
not ( n10483 , n5872 );
or ( n10484 , n10482 , n10483 );
or ( n10485 , n5872 , n4848 );
nand ( n10486 , n10484 , n10485 );
not ( n10487 , n4849 );
and ( n10488 , n5873 , n10487 );
not ( n10489 , n5873 );
and ( n10490 , n10489 , n4849 );
nor ( n10491 , n10488 , n10490 );
nand ( n10492 , n10476 , n10481 , n10486 , n10491 );
not ( n10493 , n10492 );
nand ( n10494 , n10425 , n10448 , n10471 , n10493 );
not ( n10495 , n5891 );
not ( n10496 , n4867 );
or ( n10497 , n10495 , n10496 );
or ( n10498 , n4867 , n5891 );
nand ( n10499 , n10497 , n10498 );
not ( n10500 , n5890 );
not ( n10501 , n4866 );
or ( n10502 , n10500 , n10501 );
or ( n10503 , n4866 , n5890 );
nand ( n10504 , n10502 , n10503 );
nand ( n10505 , n10499 , n10504 );
not ( n10506 , n4869 );
not ( n10507 , n5893 );
or ( n10508 , n10506 , n10507 );
or ( n10509 , n5893 , n4869 );
nand ( n10510 , n10508 , n10509 );
not ( n10511 , n4868 );
not ( n10512 , n5892 );
or ( n10513 , n10511 , n10512 );
or ( n10514 , n5892 , n4868 );
nand ( n10515 , n10513 , n10514 );
nand ( n10516 , n10510 , n10515 );
nor ( n10517 , n10505 , n10516 );
not ( n10518 , n5887 );
not ( n10519 , n4863 );
or ( n10520 , n10518 , n10519 );
or ( n10521 , n4863 , n5887 );
nand ( n10522 , n10520 , n10521 );
not ( n10523 , n5886 );
not ( n10524 , n4862 );
or ( n10525 , n10523 , n10524 );
or ( n10526 , n4862 , n5886 );
nand ( n10527 , n10525 , n10526 );
nand ( n10528 , n10522 , n10527 );
not ( n10529 , n5889 );
not ( n10530 , n4865 );
or ( n10531 , n10529 , n10530 );
or ( n10532 , n4865 , n5889 );
nand ( n10533 , n10531 , n10532 );
not ( n10534 , n5888 );
not ( n10535 , n4864 );
or ( n10536 , n10534 , n10535 );
or ( n10537 , n4864 , n5888 );
nand ( n10538 , n10536 , n10537 );
nand ( n10539 , n10533 , n10538 );
nor ( n10540 , n10528 , n10539 );
not ( n10541 , n5882 );
not ( n10542 , n4858 );
or ( n10543 , n10541 , n10542 );
or ( n10544 , n4858 , n5882 );
nand ( n10545 , n10543 , n10544 );
not ( n10546 , n5883 );
not ( n10547 , n4859 );
or ( n10548 , n10546 , n10547 );
or ( n10549 , n4859 , n5883 );
nand ( n10550 , n10548 , n10549 );
not ( n10551 , n4860 );
not ( n10552 , n5884 );
or ( n10553 , n10551 , n10552 );
or ( n10554 , n5884 , n4860 );
nand ( n10555 , n10553 , n10554 );
not ( n10556 , n4861 );
and ( n10557 , n5885 , n10556 );
not ( n10558 , n5885 );
and ( n10559 , n10558 , n4861 );
nor ( n10560 , n10557 , n10559 );
nand ( n10561 , n10545 , n10550 , n10555 , n10560 );
not ( n10562 , n10561 );
not ( n10563 , n5880 );
not ( n10564 , n4856 );
or ( n10565 , n10563 , n10564 );
or ( n10566 , n4856 , n5880 );
nand ( n10567 , n10565 , n10566 );
not ( n10568 , n4854 );
not ( n10569 , n5878 );
or ( n10570 , n10568 , n10569 );
or ( n10571 , n5878 , n4854 );
nand ( n10572 , n10570 , n10571 );
not ( n10573 , n4857 );
and ( n10574 , n5881 , n10573 );
not ( n10575 , n5881 );
and ( n10576 , n10575 , n4857 );
nor ( n10577 , n10574 , n10576 );
not ( n10578 , n4855 );
and ( n10579 , n5879 , n10578 );
not ( n10580 , n5879 );
and ( n10581 , n10580 , n4855 );
nor ( n10582 , n10579 , n10581 );
nand ( n10583 , n10567 , n10572 , n10577 , n10582 );
not ( n10584 , n10583 );
nand ( n10585 , n10517 , n10540 , n10562 , n10584 );
nor ( n10586 , n10494 , n10585 );
nand ( n10587 , n10038 , n10218 , n10402 , n10586 );
nor ( n10588 , n9853 , n10587 );
not ( n10589 , n5899 );
not ( n10590 , n4875 );
or ( n10591 , n10589 , n10590 );
or ( n10592 , n4875 , n5899 );
nand ( n10593 , n10591 , n10592 );
not ( n10594 , n5898 );
not ( n10595 , n4874 );
or ( n10596 , n10594 , n10595 );
or ( n10597 , n4874 , n5898 );
nand ( n10598 , n10596 , n10597 );
nand ( n10599 , n10593 , n10598 );
not ( n10600 , n5901 );
not ( n10601 , n4877 );
or ( n10602 , n10600 , n10601 );
or ( n10603 , n4877 , n5901 );
nand ( n10604 , n10602 , n10603 );
not ( n10605 , n5900 );
not ( n10606 , n4876 );
or ( n10607 , n10605 , n10606 );
or ( n10608 , n4876 , n5900 );
nand ( n10609 , n10607 , n10608 );
nand ( n10610 , n10604 , n10609 );
nor ( n10611 , n10599 , n10610 );
not ( n10612 , n5907 );
not ( n10613 , n4883 );
or ( n10614 , n10612 , n10613 );
or ( n10615 , n4883 , n5907 );
nand ( n10616 , n10614 , n10615 );
not ( n10617 , n5906 );
not ( n10618 , n4882 );
or ( n10619 , n10617 , n10618 );
or ( n10620 , n4882 , n5906 );
nand ( n10621 , n10619 , n10620 );
nand ( n10622 , n10616 , n10621 );
not ( n10623 , n5909 );
not ( n10624 , n4885 );
or ( n10625 , n10623 , n10624 );
or ( n10626 , n4885 , n5909 );
nand ( n10627 , n10625 , n10626 );
not ( n10628 , n5908 );
not ( n10629 , n4884 );
or ( n10630 , n10628 , n10629 );
or ( n10631 , n4884 , n5908 );
nand ( n10632 , n10630 , n10631 );
nand ( n10633 , n10627 , n10632 );
nor ( n10634 , n10622 , n10633 );
not ( n10635 , n5895 );
not ( n10636 , n4871 );
or ( n10637 , n10635 , n10636 );
or ( n10638 , n4871 , n5895 );
nand ( n10639 , n10637 , n10638 );
not ( n10640 , n5894 );
not ( n10641 , n4870 );
or ( n10642 , n10640 , n10641 );
or ( n10643 , n4870 , n5894 );
nand ( n10644 , n10642 , n10643 );
nand ( n10645 , n10639 , n10644 );
not ( n10646 , n5897 );
not ( n10647 , n4873 );
or ( n10648 , n10646 , n10647 );
or ( n10649 , n4873 , n5897 );
nand ( n10650 , n10648 , n10649 );
not ( n10651 , n5896 );
not ( n10652 , n4872 );
or ( n10653 , n10651 , n10652 );
or ( n10654 , n4872 , n5896 );
nand ( n10655 , n10653 , n10654 );
nand ( n10656 , n10650 , n10655 );
nor ( n10657 , n10645 , n10656 );
not ( n10658 , n5904 );
not ( n10659 , n4880 );
or ( n10660 , n10658 , n10659 );
or ( n10661 , n4880 , n5904 );
nand ( n10662 , n10660 , n10661 );
not ( n10663 , n5905 );
not ( n10664 , n4881 );
or ( n10665 , n10663 , n10664 );
or ( n10666 , n4881 , n5905 );
nand ( n10667 , n10665 , n10666 );
not ( n10668 , n5902 );
not ( n10669 , n4878 );
or ( n10670 , n10668 , n10669 );
or ( n10671 , n4878 , n5902 );
nand ( n10672 , n10670 , n10671 );
not ( n10673 , n5903 );
not ( n10674 , n4879 );
or ( n10675 , n10673 , n10674 );
or ( n10676 , n4879 , n5903 );
nand ( n10677 , n10675 , n10676 );
and ( n10678 , n10662 , n10667 , n10672 , n10677 );
nand ( n10679 , n10611 , n10634 , n10657 , n10678 );
not ( n10680 , n5923 );
not ( n10681 , n4899 );
or ( n10682 , n10680 , n10681 );
or ( n10683 , n4899 , n5923 );
nand ( n10684 , n10682 , n10683 );
not ( n10685 , n5922 );
not ( n10686 , n4898 );
or ( n10687 , n10685 , n10686 );
or ( n10688 , n4898 , n5922 );
nand ( n10689 , n10687 , n10688 );
nand ( n10690 , n10684 , n10689 );
not ( n10691 , n5925 );
not ( n10692 , n4901 );
or ( n10693 , n10691 , n10692 );
or ( n10694 , n4901 , n5925 );
nand ( n10695 , n10693 , n10694 );
not ( n10696 , n5924 );
not ( n10697 , n4900 );
or ( n10698 , n10696 , n10697 );
or ( n10699 , n4900 , n5924 );
nand ( n10700 , n10698 , n10699 );
nand ( n10701 , n10695 , n10700 );
nor ( n10702 , n10690 , n10701 );
not ( n10703 , n5919 );
not ( n10704 , n4895 );
or ( n10705 , n10703 , n10704 );
or ( n10706 , n4895 , n5919 );
nand ( n10707 , n10705 , n10706 );
not ( n10708 , n5918 );
not ( n10709 , n4894 );
or ( n10710 , n10708 , n10709 );
or ( n10711 , n4894 , n5918 );
nand ( n10712 , n10710 , n10711 );
nand ( n10713 , n10707 , n10712 );
not ( n10714 , n5921 );
not ( n10715 , n4897 );
or ( n10716 , n10714 , n10715 );
or ( n10717 , n4897 , n5921 );
nand ( n10718 , n10716 , n10717 );
not ( n10719 , n5920 );
not ( n10720 , n4896 );
or ( n10721 , n10719 , n10720 );
or ( n10722 , n4896 , n5920 );
nand ( n10723 , n10721 , n10722 );
nand ( n10724 , n10718 , n10723 );
nor ( n10725 , n10713 , n10724 );
not ( n10726 , n5915 );
not ( n10727 , n4891 );
or ( n10728 , n10726 , n10727 );
or ( n10729 , n4891 , n5915 );
nand ( n10730 , n10728 , n10729 );
not ( n10731 , n5914 );
not ( n10732 , n4890 );
or ( n10733 , n10731 , n10732 );
or ( n10734 , n4890 , n5914 );
nand ( n10735 , n10733 , n10734 );
nand ( n10736 , n10730 , n10735 );
not ( n10737 , n5917 );
not ( n10738 , n4893 );
or ( n10739 , n10737 , n10738 );
or ( n10740 , n4893 , n5917 );
nand ( n10741 , n10739 , n10740 );
not ( n10742 , n5916 );
not ( n10743 , n4892 );
or ( n10744 , n10742 , n10743 );
or ( n10745 , n4892 , n5916 );
nand ( n10746 , n10744 , n10745 );
nand ( n10747 , n10741 , n10746 );
nor ( n10748 , n10736 , n10747 );
not ( n10749 , n5911 );
not ( n10750 , n4887 );
or ( n10751 , n10749 , n10750 );
or ( n10752 , n4887 , n5911 );
nand ( n10753 , n10751 , n10752 );
not ( n10754 , n5910 );
not ( n10755 , n4886 );
or ( n10756 , n10754 , n10755 );
or ( n10757 , n4886 , n5910 );
nand ( n10758 , n10756 , n10757 );
nand ( n10759 , n10753 , n10758 );
not ( n10760 , n5913 );
not ( n10761 , n4889 );
or ( n10762 , n10760 , n10761 );
or ( n10763 , n4889 , n5913 );
nand ( n10764 , n10762 , n10763 );
not ( n10765 , n5912 );
not ( n10766 , n4888 );
or ( n10767 , n10765 , n10766 );
or ( n10768 , n4888 , n5912 );
nand ( n10769 , n10767 , n10768 );
nand ( n10770 , n10764 , n10769 );
nor ( n10771 , n10759 , n10770 );
nand ( n10772 , n10702 , n10725 , n10748 , n10771 );
nor ( n10773 , n10679 , n10772 );
not ( n10774 , n5971 );
not ( n10775 , n4947 );
or ( n10776 , n10774 , n10775 );
or ( n10777 , n4947 , n5971 );
nand ( n10778 , n10776 , n10777 );
not ( n10779 , n5970 );
not ( n10780 , n4946 );
or ( n10781 , n10779 , n10780 );
or ( n10782 , n4946 , n5970 );
nand ( n10783 , n10781 , n10782 );
nand ( n10784 , n10778 , n10783 );
not ( n10785 , n5973 );
not ( n10786 , n4949 );
or ( n10787 , n10785 , n10786 );
or ( n10788 , n4949 , n5973 );
nand ( n10789 , n10787 , n10788 );
not ( n10790 , n5972 );
not ( n10791 , n4948 );
or ( n10792 , n10790 , n10791 );
or ( n10793 , n4948 , n5972 );
nand ( n10794 , n10792 , n10793 );
nand ( n10795 , n10789 , n10794 );
nor ( n10796 , n10784 , n10795 );
not ( n10797 , n5967 );
not ( n10798 , n4943 );
or ( n10799 , n10797 , n10798 );
or ( n10800 , n4943 , n5967 );
nand ( n10801 , n10799 , n10800 );
not ( n10802 , n5966 );
not ( n10803 , n4942 );
or ( n10804 , n10802 , n10803 );
or ( n10805 , n4942 , n5966 );
nand ( n10806 , n10804 , n10805 );
nand ( n10807 , n10801 , n10806 );
not ( n10808 , n5969 );
not ( n10809 , n4945 );
or ( n10810 , n10808 , n10809 );
or ( n10811 , n4945 , n5969 );
nand ( n10812 , n10810 , n10811 );
not ( n10813 , n5968 );
not ( n10814 , n4944 );
or ( n10815 , n10813 , n10814 );
or ( n10816 , n4944 , n5968 );
nand ( n10817 , n10815 , n10816 );
nand ( n10818 , n10812 , n10817 );
nor ( n10819 , n10807 , n10818 );
not ( n10820 , n5960 );
not ( n10821 , n4936 );
or ( n10822 , n10820 , n10821 );
or ( n10823 , n4936 , n5960 );
nand ( n10824 , n10822 , n10823 );
not ( n10825 , n5961 );
not ( n10826 , n4937 );
or ( n10827 , n10825 , n10826 );
or ( n10828 , n4937 , n5961 );
nand ( n10829 , n10827 , n10828 );
not ( n10830 , n5958 );
not ( n10831 , n4934 );
or ( n10832 , n10830 , n10831 );
or ( n10833 , n4934 , n5958 );
nand ( n10834 , n10832 , n10833 );
not ( n10835 , n5959 );
not ( n10836 , n4935 );
or ( n10837 , n10835 , n10836 );
or ( n10838 , n4935 , n5959 );
nand ( n10839 , n10837 , n10838 );
and ( n10840 , n10824 , n10829 , n10834 , n10839 );
not ( n10841 , n5963 );
not ( n10842 , n4939 );
or ( n10843 , n10841 , n10842 );
or ( n10844 , n4939 , n5963 );
nand ( n10845 , n10843 , n10844 );
not ( n10846 , n5962 );
not ( n10847 , n4938 );
or ( n10848 , n10846 , n10847 );
or ( n10849 , n4938 , n5962 );
nand ( n10850 , n10848 , n10849 );
nand ( n10851 , n10845 , n10850 );
not ( n10852 , n5965 );
not ( n10853 , n4941 );
or ( n10854 , n10852 , n10853 );
or ( n10855 , n4941 , n5965 );
nand ( n10856 , n10854 , n10855 );
not ( n10857 , n5964 );
not ( n10858 , n4940 );
or ( n10859 , n10857 , n10858 );
or ( n10860 , n4940 , n5964 );
nand ( n10861 , n10859 , n10860 );
nand ( n10862 , n10856 , n10861 );
nor ( n10863 , n10851 , n10862 );
nand ( n10864 , n10796 , n10819 , n10840 , n10863 );
not ( n10865 , n5987 );
not ( n10866 , n4963 );
or ( n10867 , n10865 , n10866 );
or ( n10868 , n4963 , n5987 );
nand ( n10869 , n10867 , n10868 );
not ( n10870 , n5986 );
not ( n10871 , n4962 );
or ( n10872 , n10870 , n10871 );
or ( n10873 , n4962 , n5986 );
nand ( n10874 , n10872 , n10873 );
nand ( n10875 , n10869 , n10874 );
not ( n10876 , n5989 );
not ( n10877 , n4965 );
or ( n10878 , n10876 , n10877 );
or ( n10879 , n4965 , n5989 );
nand ( n10880 , n10878 , n10879 );
not ( n10881 , n5988 );
not ( n10882 , n4964 );
or ( n10883 , n10881 , n10882 );
or ( n10884 , n4964 , n5988 );
nand ( n10885 , n10883 , n10884 );
nand ( n10886 , n10880 , n10885 );
nor ( n10887 , n10875 , n10886 );
not ( n10888 , n5976 );
not ( n10889 , n4952 );
or ( n10890 , n10888 , n10889 );
or ( n10891 , n4952 , n5976 );
nand ( n10892 , n10890 , n10891 );
not ( n10893 , n5977 );
not ( n10894 , n4953 );
or ( n10895 , n10893 , n10894 );
or ( n10896 , n4953 , n5977 );
nand ( n10897 , n10895 , n10896 );
not ( n10898 , n5974 );
not ( n10899 , n4950 );
or ( n10900 , n10898 , n10899 );
or ( n10901 , n4950 , n5974 );
nand ( n10902 , n10900 , n10901 );
not ( n10903 , n5975 );
not ( n10904 , n4951 );
or ( n10905 , n10903 , n10904 );
or ( n10906 , n4951 , n5975 );
nand ( n10907 , n10905 , n10906 );
and ( n10908 , n10892 , n10897 , n10902 , n10907 );
not ( n10909 , n5979 );
not ( n10910 , n4955 );
or ( n10911 , n10909 , n10910 );
or ( n10912 , n4955 , n5979 );
nand ( n10913 , n10911 , n10912 );
not ( n10914 , n5978 );
not ( n10915 , n4954 );
or ( n10916 , n10914 , n10915 );
or ( n10917 , n4954 , n5978 );
nand ( n10918 , n10916 , n10917 );
nand ( n10919 , n10913 , n10918 );
not ( n10920 , n5981 );
not ( n10921 , n4957 );
or ( n10922 , n10920 , n10921 );
or ( n10923 , n4957 , n5981 );
nand ( n10924 , n10922 , n10923 );
not ( n10925 , n5980 );
not ( n10926 , n4956 );
or ( n10927 , n10925 , n10926 );
or ( n10928 , n4956 , n5980 );
nand ( n10929 , n10927 , n10928 );
nand ( n10930 , n10924 , n10929 );
nor ( n10931 , n10919 , n10930 );
not ( n10932 , n5985 );
not ( n10933 , n4961 );
or ( n10934 , n10932 , n10933 );
or ( n10935 , n4961 , n5985 );
nand ( n10936 , n10934 , n10935 );
not ( n10937 , n5984 );
not ( n10938 , n4960 );
or ( n10939 , n10937 , n10938 );
or ( n10940 , n4960 , n5984 );
nand ( n10941 , n10939 , n10940 );
nand ( n10942 , n10936 , n10941 );
not ( n10943 , n5983 );
not ( n10944 , n4959 );
or ( n10945 , n10943 , n10944 );
or ( n10946 , n4959 , n5983 );
nand ( n10947 , n10945 , n10946 );
not ( n10948 , n5982 );
not ( n10949 , n4958 );
or ( n10950 , n10948 , n10949 );
or ( n10951 , n4958 , n5982 );
nand ( n10952 , n10950 , n10951 );
nand ( n10953 , n10947 , n10952 );
nor ( n10954 , n10942 , n10953 );
nand ( n10955 , n10887 , n10908 , n10931 , n10954 );
nor ( n10956 , n10864 , n10955 );
not ( n10957 , n5935 );
not ( n10958 , n4911 );
or ( n10959 , n10957 , n10958 );
or ( n10960 , n4911 , n5935 );
nand ( n10961 , n10959 , n10960 );
not ( n10962 , n5934 );
not ( n10963 , n4910 );
or ( n10964 , n10962 , n10963 );
or ( n10965 , n4910 , n5934 );
nand ( n10966 , n10964 , n10965 );
nand ( n10967 , n10961 , n10966 );
not ( n10968 , n5937 );
not ( n10969 , n4913 );
or ( n10970 , n10968 , n10969 );
or ( n10971 , n4913 , n5937 );
nand ( n10972 , n10970 , n10971 );
not ( n10973 , n5936 );
not ( n10974 , n4912 );
or ( n10975 , n10973 , n10974 );
or ( n10976 , n4912 , n5936 );
nand ( n10977 , n10975 , n10976 );
nand ( n10978 , n10972 , n10977 );
nor ( n10979 , n10967 , n10978 );
not ( n10980 , n5931 );
not ( n10981 , n4907 );
or ( n10982 , n10980 , n10981 );
or ( n10983 , n4907 , n5931 );
nand ( n10984 , n10982 , n10983 );
not ( n10985 , n5930 );
not ( n10986 , n4906 );
or ( n10987 , n10985 , n10986 );
or ( n10988 , n4906 , n5930 );
nand ( n10989 , n10987 , n10988 );
nand ( n10990 , n10984 , n10989 );
not ( n10991 , n5933 );
not ( n10992 , n4909 );
or ( n10993 , n10991 , n10992 );
or ( n10994 , n4909 , n5933 );
nand ( n10995 , n10993 , n10994 );
not ( n10996 , n5932 );
not ( n10997 , n4908 );
or ( n10998 , n10996 , n10997 );
or ( n10999 , n4908 , n5932 );
nand ( n11000 , n10998 , n10999 );
nand ( n11001 , n10995 , n11000 );
nor ( n11002 , n10990 , n11001 );
not ( n11003 , n5940 );
not ( n11004 , n4916 );
or ( n11005 , n11003 , n11004 );
or ( n11006 , n4916 , n5940 );
nand ( n11007 , n11005 , n11006 );
not ( n11008 , n5941 );
not ( n11009 , n4917 );
or ( n11010 , n11008 , n11009 );
or ( n11011 , n4917 , n5941 );
nand ( n11012 , n11010 , n11011 );
not ( n11013 , n5938 );
not ( n11014 , n4914 );
or ( n11015 , n11013 , n11014 );
or ( n11016 , n4914 , n5938 );
nand ( n11017 , n11015 , n11016 );
not ( n11018 , n5939 );
not ( n11019 , n4915 );
or ( n11020 , n11018 , n11019 );
or ( n11021 , n4915 , n5939 );
nand ( n11022 , n11020 , n11021 );
nand ( n11023 , n11007 , n11012 , n11017 , n11022 );
not ( n11024 , n11023 );
not ( n11025 , n5927 );
not ( n11026 , n4903 );
or ( n11027 , n11025 , n11026 );
or ( n11028 , n4903 , n5927 );
nand ( n11029 , n11027 , n11028 );
not ( n11030 , n5926 );
not ( n11031 , n4902 );
or ( n11032 , n11030 , n11031 );
or ( n11033 , n4902 , n5926 );
nand ( n11034 , n11032 , n11033 );
nand ( n11035 , n11029 , n11034 );
not ( n11036 , n5929 );
not ( n11037 , n4905 );
or ( n11038 , n11036 , n11037 );
or ( n11039 , n4905 , n5929 );
nand ( n11040 , n11038 , n11039 );
not ( n11041 , n5928 );
not ( n11042 , n4904 );
or ( n11043 , n11041 , n11042 );
or ( n11044 , n4904 , n5928 );
nand ( n11045 , n11043 , n11044 );
nand ( n11046 , n11040 , n11045 );
nor ( n11047 , n11035 , n11046 );
nand ( n11048 , n10979 , n11002 , n11024 , n11047 );
not ( n11049 , n5944 );
not ( n11050 , n4920 );
or ( n11051 , n11049 , n11050 );
or ( n11052 , n4920 , n5944 );
nand ( n11053 , n11051 , n11052 );
not ( n11054 , n5945 );
not ( n11055 , n4921 );
or ( n11056 , n11054 , n11055 );
or ( n11057 , n4921 , n5945 );
nand ( n11058 , n11056 , n11057 );
not ( n11059 , n5942 );
not ( n11060 , n4918 );
or ( n11061 , n11059 , n11060 );
or ( n11062 , n4918 , n5942 );
nand ( n11063 , n11061 , n11062 );
not ( n11064 , n5943 );
not ( n11065 , n4919 );
or ( n11066 , n11064 , n11065 );
or ( n11067 , n4919 , n5943 );
nand ( n11068 , n11066 , n11067 );
and ( n11069 , n11053 , n11058 , n11063 , n11068 );
not ( n11070 , n5952 );
not ( n11071 , n4928 );
or ( n11072 , n11070 , n11071 );
or ( n11073 , n4928 , n5952 );
nand ( n11074 , n11072 , n11073 );
not ( n11075 , n5953 );
not ( n11076 , n4929 );
or ( n11077 , n11075 , n11076 );
or ( n11078 , n4929 , n5953 );
nand ( n11079 , n11077 , n11078 );
not ( n11080 , n5950 );
not ( n11081 , n4926 );
or ( n11082 , n11080 , n11081 );
or ( n11083 , n4926 , n5950 );
nand ( n11084 , n11082 , n11083 );
not ( n11085 , n5951 );
not ( n11086 , n4927 );
or ( n11087 , n11085 , n11086 );
or ( n11088 , n4927 , n5951 );
nand ( n11089 , n11087 , n11088 );
nand ( n11090 , n11074 , n11079 , n11084 , n11089 );
not ( n11091 , n11090 );
not ( n11092 , n4924 );
not ( n11093 , n5948 );
or ( n11094 , n11092 , n11093 );
or ( n11095 , n5948 , n4924 );
nand ( n11096 , n11094 , n11095 );
not ( n11097 , n4925 );
not ( n11098 , n5949 );
or ( n11099 , n11097 , n11098 );
or ( n11100 , n5949 , n4925 );
nand ( n11101 , n11099 , n11100 );
nand ( n11102 , n11096 , n11101 );
not ( n11103 , n4922 );
not ( n11104 , n5946 );
or ( n11105 , n11103 , n11104 );
or ( n11106 , n5946 , n4922 );
nand ( n11107 , n11105 , n11106 );
not ( n11108 , n4923 );
not ( n11109 , n5947 );
or ( n11110 , n11108 , n11109 );
or ( n11111 , n5947 , n4923 );
nand ( n11112 , n11110 , n11111 );
nand ( n11113 , n11107 , n11112 );
nor ( n11114 , n11102 , n11113 );
not ( n11115 , n4933 );
not ( n11116 , n5957 );
or ( n11117 , n11115 , n11116 );
or ( n11118 , n5957 , n4933 );
nand ( n11119 , n11117 , n11118 );
not ( n11120 , n4932 );
not ( n11121 , n5956 );
or ( n11122 , n11120 , n11121 );
or ( n11123 , n5956 , n4932 );
nand ( n11124 , n11122 , n11123 );
nand ( n11125 , n11119 , n11124 );
not ( n11126 , n4931 );
not ( n11127 , n5955 );
or ( n11128 , n11126 , n11127 );
or ( n11129 , n5955 , n4931 );
nand ( n11130 , n11128 , n11129 );
not ( n11131 , n4930 );
not ( n11132 , n5954 );
or ( n11133 , n11131 , n11132 );
or ( n11134 , n5954 , n4930 );
nand ( n11135 , n11133 , n11134 );
nand ( n11136 , n11130 , n11135 );
nor ( n11137 , n11125 , n11136 );
nand ( n11138 , n11069 , n11091 , n11114 , n11137 );
nor ( n11139 , n11048 , n11138 );
not ( n11140 , n6003 );
not ( n11141 , n4979 );
or ( n11142 , n11140 , n11141 );
or ( n11143 , n4979 , n6003 );
nand ( n11144 , n11142 , n11143 );
not ( n11145 , n6002 );
not ( n11146 , n4978 );
or ( n11147 , n11145 , n11146 );
or ( n11148 , n4978 , n6002 );
nand ( n11149 , n11147 , n11148 );
nand ( n11150 , n11144 , n11149 );
not ( n11151 , n6005 );
not ( n11152 , n4981 );
or ( n11153 , n11151 , n11152 );
or ( n11154 , n4981 , n6005 );
nand ( n11155 , n11153 , n11154 );
not ( n11156 , n6004 );
not ( n11157 , n4980 );
or ( n11158 , n11156 , n11157 );
or ( n11159 , n4980 , n6004 );
nand ( n11160 , n11158 , n11159 );
nand ( n11161 , n11155 , n11160 );
nor ( n11162 , n11150 , n11161 );
not ( n11163 , n5991 );
not ( n11164 , n4967 );
or ( n11165 , n11163 , n11164 );
or ( n11166 , n4967 , n5991 );
nand ( n11167 , n11165 , n11166 );
not ( n11168 , n5990 );
not ( n11169 , n4966 );
or ( n11170 , n11168 , n11169 );
or ( n11171 , n4966 , n5990 );
nand ( n11172 , n11170 , n11171 );
not ( n11173 , n5993 );
not ( n11174 , n4969 );
or ( n11175 , n11173 , n11174 );
or ( n11176 , n4969 , n5993 );
nand ( n11177 , n11175 , n11176 );
not ( n11178 , n5992 );
not ( n11179 , n4968 );
or ( n11180 , n11178 , n11179 );
or ( n11181 , n4968 , n5992 );
nand ( n11182 , n11180 , n11181 );
nand ( n11183 , n11167 , n11172 , n11177 , n11182 );
not ( n11184 , n11183 );
not ( n11185 , n5997 );
not ( n11186 , n4973 );
or ( n11187 , n11185 , n11186 );
or ( n11188 , n4973 , n5997 );
nand ( n11189 , n11187 , n11188 );
not ( n11190 , n5996 );
not ( n11191 , n4972 );
or ( n11192 , n11190 , n11191 );
or ( n11193 , n4972 , n5996 );
nand ( n11194 , n11192 , n11193 );
nand ( n11195 , n11189 , n11194 );
not ( n11196 , n5995 );
not ( n11197 , n4971 );
or ( n11198 , n11196 , n11197 );
or ( n11199 , n4971 , n5995 );
nand ( n11200 , n11198 , n11199 );
not ( n11201 , n5994 );
not ( n11202 , n4970 );
or ( n11203 , n11201 , n11202 );
or ( n11204 , n4970 , n5994 );
nand ( n11205 , n11203 , n11204 );
nand ( n11206 , n11200 , n11205 );
nor ( n11207 , n11195 , n11206 );
not ( n11208 , n6000 );
not ( n11209 , n4976 );
or ( n11210 , n11208 , n11209 );
or ( n11211 , n4976 , n6000 );
nand ( n11212 , n11210 , n11211 );
not ( n11213 , n6001 );
not ( n11214 , n4977 );
or ( n11215 , n11213 , n11214 );
or ( n11216 , n4977 , n6001 );
nand ( n11217 , n11215 , n11216 );
not ( n11218 , n4974 );
not ( n11219 , n5998 );
or ( n11220 , n11218 , n11219 );
or ( n11221 , n5998 , n4974 );
nand ( n11222 , n11220 , n11221 );
not ( n11223 , n4975 );
and ( n11224 , n5999 , n11223 );
not ( n11225 , n5999 );
and ( n11226 , n11225 , n4975 );
nor ( n11227 , n11224 , n11226 );
nand ( n11228 , n11212 , n11217 , n11222 , n11227 );
not ( n11229 , n11228 );
nand ( n11230 , n11162 , n11184 , n11207 , n11229 );
not ( n11231 , n4994 );
not ( n11232 , n6018 );
or ( n11233 , n11231 , n11232 );
or ( n11234 , n6018 , n4994 );
nand ( n11235 , n11233 , n11234 );
not ( n11236 , n4995 );
not ( n11237 , n6019 );
or ( n11238 , n11236 , n11237 );
or ( n11239 , n6019 , n4995 );
nand ( n11240 , n11238 , n11239 );
nand ( n11241 , n11235 , n11240 );
not ( n11242 , n6021 );
not ( n11243 , n4997 );
or ( n11244 , n11242 , n11243 );
or ( n11245 , n4997 , n6021 );
nand ( n11246 , n11244 , n11245 );
not ( n11247 , n6020 );
not ( n11248 , n4996 );
or ( n11249 , n11247 , n11248 );
or ( n11250 , n4996 , n6020 );
nand ( n11251 , n11249 , n11250 );
nand ( n11252 , n11246 , n11251 );
nor ( n11253 , n11241 , n11252 );
not ( n11254 , n6015 );
not ( n11255 , n4991 );
or ( n11256 , n11254 , n11255 );
or ( n11257 , n4991 , n6015 );
nand ( n11258 , n11256 , n11257 );
not ( n11259 , n6014 );
not ( n11260 , n4990 );
or ( n11261 , n11259 , n11260 );
or ( n11262 , n4990 , n6014 );
nand ( n11263 , n11261 , n11262 );
nand ( n11264 , n11258 , n11263 );
not ( n11265 , n6017 );
not ( n11266 , n4993 );
or ( n11267 , n11265 , n11266 );
or ( n11268 , n4993 , n6017 );
nand ( n11269 , n11267 , n11268 );
not ( n11270 , n6016 );
not ( n11271 , n4992 );
or ( n11272 , n11270 , n11271 );
or ( n11273 , n4992 , n6016 );
nand ( n11274 , n11272 , n11273 );
nand ( n11275 , n11269 , n11274 );
nor ( n11276 , n11264 , n11275 );
not ( n11277 , n6011 );
not ( n11278 , n4987 );
or ( n11279 , n11277 , n11278 );
or ( n11280 , n4987 , n6011 );
nand ( n11281 , n11279 , n11280 );
not ( n11282 , n6010 );
not ( n11283 , n4986 );
or ( n11284 , n11282 , n11283 );
or ( n11285 , n4986 , n6010 );
nand ( n11286 , n11284 , n11285 );
nand ( n11287 , n11281 , n11286 );
not ( n11288 , n6013 );
not ( n11289 , n4989 );
or ( n11290 , n11288 , n11289 );
or ( n11291 , n4989 , n6013 );
nand ( n11292 , n11290 , n11291 );
not ( n11293 , n6012 );
not ( n11294 , n4988 );
or ( n11295 , n11293 , n11294 );
or ( n11296 , n4988 , n6012 );
nand ( n11297 , n11295 , n11296 );
nand ( n11298 , n11292 , n11297 );
nor ( n11299 , n11287 , n11298 );
not ( n11300 , n6008 );
not ( n11301 , n4984 );
or ( n11302 , n11300 , n11301 );
or ( n11303 , n4984 , n6008 );
nand ( n11304 , n11302 , n11303 );
not ( n11305 , n4982 );
not ( n11306 , n6006 );
or ( n11307 , n11305 , n11306 );
or ( n11308 , n6006 , n4982 );
nand ( n11309 , n11307 , n11308 );
not ( n11310 , n4985 );
and ( n11311 , n6009 , n11310 );
not ( n11312 , n6009 );
and ( n11313 , n11312 , n4985 );
nor ( n11314 , n11311 , n11313 );
not ( n11315 , n4983 );
and ( n11316 , n6007 , n11315 );
not ( n11317 , n6007 );
and ( n11318 , n11317 , n4983 );
nor ( n11319 , n11316 , n11318 );
nand ( n11320 , n11304 , n11309 , n11314 , n11319 );
not ( n11321 , n11320 );
nand ( n11322 , n11253 , n11276 , n11299 , n11321 );
nor ( n11323 , n11230 , n11322 );
nand ( n11324 , n10773 , n10956 , n11139 , n11323 );
not ( n11325 , n6031 );
not ( n11326 , n5007 );
or ( n11327 , n11325 , n11326 );
or ( n11328 , n5007 , n6031 );
nand ( n11329 , n11327 , n11328 );
not ( n11330 , n6033 );
not ( n11331 , n5009 );
or ( n11332 , n11330 , n11331 );
or ( n11333 , n5009 , n6033 );
nand ( n11334 , n11332 , n11333 );
not ( n11335 , n6030 );
not ( n11336 , n5006 );
or ( n11337 , n11335 , n11336 );
or ( n11338 , n5006 , n6030 );
nand ( n11339 , n11337 , n11338 );
not ( n11340 , n6032 );
not ( n11341 , n5008 );
or ( n11342 , n11340 , n11341 );
or ( n11343 , n5008 , n6032 );
nand ( n11344 , n11342 , n11343 );
nand ( n11345 , n11329 , n11334 , n11339 , n11344 );
not ( n11346 , n11345 );
not ( n11347 , n6027 );
not ( n11348 , n5003 );
or ( n11349 , n11347 , n11348 );
or ( n11350 , n5003 , n6027 );
nand ( n11351 , n11349 , n11350 );
not ( n11352 , n6026 );
not ( n11353 , n5002 );
or ( n11354 , n11352 , n11353 );
or ( n11355 , n5002 , n6026 );
nand ( n11356 , n11354 , n11355 );
nand ( n11357 , n11351 , n11356 );
not ( n11358 , n6029 );
not ( n11359 , n5005 );
or ( n11360 , n11358 , n11359 );
or ( n11361 , n5005 , n6029 );
nand ( n11362 , n11360 , n11361 );
not ( n11363 , n6028 );
not ( n11364 , n5004 );
or ( n11365 , n11363 , n11364 );
or ( n11366 , n5004 , n6028 );
nand ( n11367 , n11365 , n11366 );
nand ( n11368 , n11362 , n11367 );
nor ( n11369 , n11357 , n11368 );
not ( n11370 , n6035 );
not ( n11371 , n5011 );
or ( n11372 , n11370 , n11371 );
or ( n11373 , n5011 , n6035 );
nand ( n11374 , n11372 , n11373 );
not ( n11375 , n6034 );
not ( n11376 , n5010 );
or ( n11377 , n11375 , n11376 );
or ( n11378 , n5010 , n6034 );
nand ( n11379 , n11377 , n11378 );
nand ( n11380 , n11374 , n11379 );
not ( n11381 , n6037 );
not ( n11382 , n5013 );
or ( n11383 , n11381 , n11382 );
or ( n11384 , n5013 , n6037 );
nand ( n11385 , n11383 , n11384 );
not ( n11386 , n6036 );
not ( n11387 , n5012 );
or ( n11388 , n11386 , n11387 );
or ( n11389 , n5012 , n6036 );
nand ( n11390 , n11388 , n11389 );
nand ( n11391 , n11385 , n11390 );
nor ( n11392 , n11380 , n11391 );
not ( n11393 , n6023 );
not ( n11394 , n4999 );
or ( n11395 , n11393 , n11394 );
or ( n11396 , n4999 , n6023 );
nand ( n11397 , n11395 , n11396 );
not ( n11398 , n6022 );
not ( n11399 , n4998 );
or ( n11400 , n11398 , n11399 );
or ( n11401 , n4998 , n6022 );
nand ( n11402 , n11400 , n11401 );
nand ( n11403 , n11397 , n11402 );
not ( n11404 , n6025 );
not ( n11405 , n5001 );
or ( n11406 , n11404 , n11405 );
or ( n11407 , n5001 , n6025 );
nand ( n11408 , n11406 , n11407 );
not ( n11409 , n6024 );
not ( n11410 , n5000 );
or ( n11411 , n11409 , n11410 );
or ( n11412 , n5000 , n6024 );
nand ( n11413 , n11411 , n11412 );
nand ( n11414 , n11408 , n11413 );
nor ( n11415 , n11403 , n11414 );
nand ( n11416 , n11346 , n11369 , n11392 , n11415 );
not ( n11417 , n6047 );
not ( n11418 , n5023 );
or ( n11419 , n11417 , n11418 );
or ( n11420 , n5023 , n6047 );
nand ( n11421 , n11419 , n11420 );
not ( n11422 , n6046 );
not ( n11423 , n5022 );
or ( n11424 , n11422 , n11423 );
or ( n11425 , n5022 , n6046 );
nand ( n11426 , n11424 , n11425 );
nand ( n11427 , n11421 , n11426 );
not ( n11428 , n6049 );
not ( n11429 , n5025 );
or ( n11430 , n11428 , n11429 );
or ( n11431 , n5025 , n6049 );
nand ( n11432 , n11430 , n11431 );
not ( n11433 , n6048 );
not ( n11434 , n5024 );
or ( n11435 , n11433 , n11434 );
or ( n11436 , n5024 , n6048 );
nand ( n11437 , n11435 , n11436 );
nand ( n11438 , n11432 , n11437 );
nor ( n11439 , n11427 , n11438 );
not ( n11440 , n6051 );
not ( n11441 , n5027 );
or ( n11442 , n11440 , n11441 );
or ( n11443 , n5027 , n6051 );
nand ( n11444 , n11442 , n11443 );
not ( n11445 , n6050 );
not ( n11446 , n5026 );
or ( n11447 , n11445 , n11446 );
or ( n11448 , n5026 , n6050 );
nand ( n11449 , n11447 , n11448 );
nand ( n11450 , n11444 , n11449 );
not ( n11451 , n6053 );
not ( n11452 , n5029 );
or ( n11453 , n11451 , n11452 );
or ( n11454 , n5029 , n6053 );
nand ( n11455 , n11453 , n11454 );
not ( n11456 , n6052 );
not ( n11457 , n5028 );
or ( n11458 , n11456 , n11457 );
or ( n11459 , n5028 , n6052 );
nand ( n11460 , n11458 , n11459 );
nand ( n11461 , n11455 , n11460 );
nor ( n11462 , n11450 , n11461 );
not ( n11463 , n6039 );
not ( n11464 , n5015 );
or ( n11465 , n11463 , n11464 );
or ( n11466 , n5015 , n6039 );
nand ( n11467 , n11465 , n11466 );
not ( n11468 , n6038 );
not ( n11469 , n5014 );
or ( n11470 , n11468 , n11469 );
or ( n11471 , n5014 , n6038 );
nand ( n11472 , n11470 , n11471 );
nand ( n11473 , n11467 , n11472 );
not ( n11474 , n6041 );
not ( n11475 , n5017 );
or ( n11476 , n11474 , n11475 );
or ( n11477 , n5017 , n6041 );
nand ( n11478 , n11476 , n11477 );
not ( n11479 , n6040 );
not ( n11480 , n5016 );
or ( n11481 , n11479 , n11480 );
or ( n11482 , n5016 , n6040 );
nand ( n11483 , n11481 , n11482 );
nand ( n11484 , n11478 , n11483 );
nor ( n11485 , n11473 , n11484 );
not ( n11486 , n6043 );
not ( n11487 , n5019 );
or ( n11488 , n11486 , n11487 );
or ( n11489 , n5019 , n6043 );
nand ( n11490 , n11488 , n11489 );
not ( n11491 , n6045 );
not ( n11492 , n5021 );
or ( n11493 , n11491 , n11492 );
or ( n11494 , n5021 , n6045 );
nand ( n11495 , n11493 , n11494 );
not ( n11496 , n6042 );
not ( n11497 , n5018 );
or ( n11498 , n11496 , n11497 );
or ( n11499 , n5018 , n6042 );
nand ( n11500 , n11498 , n11499 );
not ( n11501 , n6044 );
not ( n11502 , n5020 );
or ( n11503 , n11501 , n11502 );
or ( n11504 , n5020 , n6044 );
nand ( n11505 , n11503 , n11504 );
nand ( n11506 , n11490 , n11495 , n11500 , n11505 );
not ( n11507 , n11506 );
nand ( n11508 , n11439 , n11462 , n11485 , n11507 );
nor ( n11509 , n11416 , n11508 );
not ( n11510 , n6072 );
not ( n11511 , n5048 );
or ( n11512 , n11510 , n11511 );
or ( n11513 , n5048 , n6072 );
nand ( n11514 , n11512 , n11513 );
not ( n11515 , n6073 );
not ( n11516 , n5049 );
or ( n11517 , n11515 , n11516 );
or ( n11518 , n5049 , n6073 );
nand ( n11519 , n11517 , n11518 );
not ( n11520 , n6070 );
not ( n11521 , n5046 );
or ( n11522 , n11520 , n11521 );
or ( n11523 , n5046 , n6070 );
nand ( n11524 , n11522 , n11523 );
not ( n11525 , n6071 );
not ( n11526 , n5047 );
or ( n11527 , n11525 , n11526 );
or ( n11528 , n5047 , n6071 );
nand ( n11529 , n11527 , n11528 );
nand ( n11530 , n11514 , n11519 , n11524 , n11529 );
not ( n11531 , n11530 );
not ( n11532 , n6083 );
not ( n11533 , n5059 );
or ( n11534 , n11532 , n11533 );
or ( n11535 , n5059 , n6083 );
nand ( n11536 , n11534 , n11535 );
not ( n11537 , n6082 );
not ( n11538 , n5058 );
or ( n11539 , n11537 , n11538 );
or ( n11540 , n5058 , n6082 );
nand ( n11541 , n11539 , n11540 );
nand ( n11542 , n11536 , n11541 );
not ( n11543 , n6085 );
not ( n11544 , n5061 );
or ( n11545 , n11543 , n11544 );
or ( n11546 , n5061 , n6085 );
nand ( n11547 , n11545 , n11546 );
not ( n11548 , n6084 );
not ( n11549 , n5060 );
or ( n11550 , n11548 , n11549 );
or ( n11551 , n5060 , n6084 );
nand ( n11552 , n11550 , n11551 );
nand ( n11553 , n11547 , n11552 );
nor ( n11554 , n11542 , n11553 );
not ( n11555 , n6079 );
not ( n11556 , n5055 );
or ( n11557 , n11555 , n11556 );
or ( n11558 , n5055 , n6079 );
nand ( n11559 , n11557 , n11558 );
not ( n11560 , n6078 );
not ( n11561 , n5054 );
or ( n11562 , n11560 , n11561 );
or ( n11563 , n5054 , n6078 );
nand ( n11564 , n11562 , n11563 );
nand ( n11565 , n11559 , n11564 );
not ( n11566 , n6081 );
not ( n11567 , n5057 );
or ( n11568 , n11566 , n11567 );
or ( n11569 , n5057 , n6081 );
nand ( n11570 , n11568 , n11569 );
not ( n11571 , n6080 );
not ( n11572 , n5056 );
or ( n11573 , n11571 , n11572 );
or ( n11574 , n5056 , n6080 );
nand ( n11575 , n11573 , n11574 );
nand ( n11576 , n11570 , n11575 );
nor ( n11577 , n11565 , n11576 );
not ( n11578 , n6075 );
not ( n11579 , n5051 );
or ( n11580 , n11578 , n11579 );
or ( n11581 , n5051 , n6075 );
nand ( n11582 , n11580 , n11581 );
not ( n11583 , n6074 );
not ( n11584 , n5050 );
or ( n11585 , n11583 , n11584 );
or ( n11586 , n5050 , n6074 );
nand ( n11587 , n11585 , n11586 );
nand ( n11588 , n11582 , n11587 );
not ( n11589 , n6077 );
not ( n11590 , n5053 );
or ( n11591 , n11589 , n11590 );
or ( n11592 , n5053 , n6077 );
nand ( n11593 , n11591 , n11592 );
not ( n11594 , n6076 );
not ( n11595 , n5052 );
or ( n11596 , n11594 , n11595 );
or ( n11597 , n5052 , n6076 );
nand ( n11598 , n11596 , n11597 );
nand ( n11599 , n11593 , n11598 );
nor ( n11600 , n11588 , n11599 );
nand ( n11601 , n11531 , n11554 , n11577 , n11600 );
not ( n11602 , n6063 );
not ( n11603 , n5039 );
or ( n11604 , n11602 , n11603 );
or ( n11605 , n5039 , n6063 );
nand ( n11606 , n11604 , n11605 );
not ( n11607 , n6062 );
not ( n11608 , n5038 );
or ( n11609 , n11607 , n11608 );
or ( n11610 , n5038 , n6062 );
nand ( n11611 , n11609 , n11610 );
nand ( n11612 , n11606 , n11611 );
not ( n11613 , n6065 );
not ( n11614 , n5041 );
or ( n11615 , n11613 , n11614 );
or ( n11616 , n5041 , n6065 );
nand ( n11617 , n11615 , n11616 );
not ( n11618 , n6064 );
not ( n11619 , n5040 );
or ( n11620 , n11618 , n11619 );
or ( n11621 , n5040 , n6064 );
nand ( n11622 , n11620 , n11621 );
nand ( n11623 , n11617 , n11622 );
nor ( n11624 , n11612 , n11623 );
not ( n11625 , n6068 );
not ( n11626 , n5044 );
or ( n11627 , n11625 , n11626 );
or ( n11628 , n5044 , n6068 );
nand ( n11629 , n11627 , n11628 );
not ( n11630 , n6069 );
not ( n11631 , n5045 );
or ( n11632 , n11630 , n11631 );
or ( n11633 , n5045 , n6069 );
nand ( n11634 , n11632 , n11633 );
not ( n11635 , n6066 );
not ( n11636 , n5042 );
or ( n11637 , n11635 , n11636 );
or ( n11638 , n5042 , n6066 );
nand ( n11639 , n11637 , n11638 );
not ( n11640 , n6067 );
not ( n11641 , n5043 );
or ( n11642 , n11640 , n11641 );
or ( n11643 , n5043 , n6067 );
nand ( n11644 , n11642 , n11643 );
nand ( n11645 , n11629 , n11634 , n11639 , n11644 );
not ( n11646 , n11645 );
not ( n11647 , n6055 );
not ( n11648 , n5031 );
or ( n11649 , n11647 , n11648 );
or ( n11650 , n5031 , n6055 );
nand ( n11651 , n11649 , n11650 );
not ( n11652 , n6054 );
not ( n11653 , n5030 );
or ( n11654 , n11652 , n11653 );
or ( n11655 , n5030 , n6054 );
nand ( n11656 , n11654 , n11655 );
nand ( n11657 , n11651 , n11656 );
not ( n11658 , n6057 );
not ( n11659 , n5033 );
or ( n11660 , n11658 , n11659 );
or ( n11661 , n5033 , n6057 );
nand ( n11662 , n11660 , n11661 );
not ( n11663 , n6056 );
not ( n11664 , n5032 );
or ( n11665 , n11663 , n11664 );
or ( n11666 , n5032 , n6056 );
nand ( n11667 , n11665 , n11666 );
nand ( n11668 , n11662 , n11667 );
nor ( n11669 , n11657 , n11668 );
not ( n11670 , n6061 );
not ( n11671 , n5037 );
or ( n11672 , n11670 , n11671 );
or ( n11673 , n5037 , n6061 );
nand ( n11674 , n11672 , n11673 );
not ( n11675 , n6060 );
not ( n11676 , n5036 );
or ( n11677 , n11675 , n11676 );
or ( n11678 , n5036 , n6060 );
nand ( n11679 , n11677 , n11678 );
nand ( n11680 , n11674 , n11679 );
not ( n11681 , n6059 );
not ( n11682 , n5035 );
or ( n11683 , n11681 , n11682 );
or ( n11684 , n5035 , n6059 );
nand ( n11685 , n11683 , n11684 );
not ( n11686 , n6058 );
not ( n11687 , n5034 );
or ( n11688 , n11686 , n11687 );
or ( n11689 , n5034 , n6058 );
nand ( n11690 , n11688 , n11689 );
nand ( n11691 , n11685 , n11690 );
nor ( n11692 , n11680 , n11691 );
nand ( n11693 , n11624 , n11646 , n11669 , n11692 );
nor ( n11694 , n11601 , n11693 );
not ( n11695 , n6099 );
not ( n11696 , n5075 );
or ( n11697 , n11695 , n11696 );
or ( n11698 , n5075 , n6099 );
nand ( n11699 , n11697 , n11698 );
not ( n11700 , n6098 );
not ( n11701 , n5074 );
or ( n11702 , n11700 , n11701 );
or ( n11703 , n5074 , n6098 );
nand ( n11704 , n11702 , n11703 );
nand ( n11705 , n11699 , n11704 );
not ( n11706 , n6101 );
not ( n11707 , n5077 );
or ( n11708 , n11706 , n11707 );
or ( n11709 , n5077 , n6101 );
nand ( n11710 , n11708 , n11709 );
not ( n11711 , n6100 );
not ( n11712 , n5076 );
or ( n11713 , n11711 , n11712 );
or ( n11714 , n5076 , n6100 );
nand ( n11715 , n11713 , n11714 );
nand ( n11716 , n11710 , n11715 );
nor ( n11717 , n11705 , n11716 );
not ( n11718 , n6088 );
not ( n11719 , n5064 );
or ( n11720 , n11718 , n11719 );
or ( n11721 , n5064 , n6088 );
nand ( n11722 , n11720 , n11721 );
not ( n11723 , n6089 );
not ( n11724 , n5065 );
or ( n11725 , n11723 , n11724 );
or ( n11726 , n5065 , n6089 );
nand ( n11727 , n11725 , n11726 );
not ( n11728 , n6086 );
not ( n11729 , n5062 );
or ( n11730 , n11728 , n11729 );
or ( n11731 , n5062 , n6086 );
nand ( n11732 , n11730 , n11731 );
not ( n11733 , n6087 );
not ( n11734 , n5063 );
or ( n11735 , n11733 , n11734 );
or ( n11736 , n5063 , n6087 );
nand ( n11737 , n11735 , n11736 );
nand ( n11738 , n11722 , n11727 , n11732 , n11737 );
not ( n11739 , n11738 );
not ( n11740 , n6091 );
not ( n11741 , n5067 );
or ( n11742 , n11740 , n11741 );
or ( n11743 , n5067 , n6091 );
nand ( n11744 , n11742 , n11743 );
not ( n11745 , n6090 );
not ( n11746 , n5066 );
or ( n11747 , n11745 , n11746 );
or ( n11748 , n5066 , n6090 );
nand ( n11749 , n11747 , n11748 );
nand ( n11750 , n11744 , n11749 );
not ( n11751 , n6093 );
not ( n11752 , n5069 );
or ( n11753 , n11751 , n11752 );
or ( n11754 , n5069 , n6093 );
nand ( n11755 , n11753 , n11754 );
not ( n11756 , n6092 );
not ( n11757 , n5068 );
or ( n11758 , n11756 , n11757 );
or ( n11759 , n5068 , n6092 );
nand ( n11760 , n11758 , n11759 );
nand ( n11761 , n11755 , n11760 );
nor ( n11762 , n11750 , n11761 );
not ( n11763 , n6096 );
not ( n11764 , n5072 );
or ( n11765 , n11763 , n11764 );
or ( n11766 , n5072 , n6096 );
nand ( n11767 , n11765 , n11766 );
not ( n11768 , n6097 );
not ( n11769 , n5073 );
or ( n11770 , n11768 , n11769 );
or ( n11771 , n5073 , n6097 );
nand ( n11772 , n11770 , n11771 );
not ( n11773 , n5070 );
not ( n11774 , n6094 );
or ( n11775 , n11773 , n11774 );
or ( n11776 , n6094 , n5070 );
nand ( n11777 , n11775 , n11776 );
not ( n11778 , n5071 );
and ( n11779 , n6095 , n11778 );
not ( n11780 , n6095 );
and ( n11781 , n11780 , n5071 );
nor ( n11782 , n11779 , n11781 );
nand ( n11783 , n11767 , n11772 , n11777 , n11782 );
not ( n11784 , n11783 );
nand ( n11785 , n11717 , n11739 , n11762 , n11784 );
not ( n11786 , n6115 );
not ( n11787 , n5091 );
or ( n11788 , n11786 , n11787 );
or ( n11789 , n5091 , n6115 );
nand ( n11790 , n11788 , n11789 );
not ( n11791 , n6114 );
not ( n11792 , n5090 );
or ( n11793 , n11791 , n11792 );
or ( n11794 , n5090 , n6114 );
nand ( n11795 , n11793 , n11794 );
nand ( n11796 , n11790 , n11795 );
not ( n11797 , n6117 );
not ( n11798 , n5093 );
or ( n11799 , n11797 , n11798 );
or ( n11800 , n5093 , n6117 );
nand ( n11801 , n11799 , n11800 );
not ( n11802 , n6116 );
not ( n11803 , n5092 );
or ( n11804 , n11802 , n11803 );
or ( n11805 , n5092 , n6116 );
nand ( n11806 , n11804 , n11805 );
nand ( n11807 , n11801 , n11806 );
nor ( n11808 , n11796 , n11807 );
not ( n11809 , n6107 );
not ( n11810 , n5083 );
or ( n11811 , n11809 , n11810 );
or ( n11812 , n5083 , n6107 );
nand ( n11813 , n11811 , n11812 );
not ( n11814 , n6106 );
not ( n11815 , n5082 );
or ( n11816 , n11814 , n11815 );
or ( n11817 , n5082 , n6106 );
nand ( n11818 , n11816 , n11817 );
nand ( n11819 , n11813 , n11818 );
not ( n11820 , n6109 );
not ( n11821 , n5085 );
or ( n11822 , n11820 , n11821 );
or ( n11823 , n5085 , n6109 );
nand ( n11824 , n11822 , n11823 );
not ( n11825 , n6108 );
not ( n11826 , n5084 );
or ( n11827 , n11825 , n11826 );
or ( n11828 , n5084 , n6108 );
nand ( n11829 , n11827 , n11828 );
nand ( n11830 , n11824 , n11829 );
nor ( n11831 , n11819 , n11830 );
not ( n11832 , n6111 );
not ( n11833 , n5087 );
or ( n11834 , n11832 , n11833 );
or ( n11835 , n5087 , n6111 );
nand ( n11836 , n11834 , n11835 );
not ( n11837 , n6110 );
not ( n11838 , n5086 );
or ( n11839 , n11837 , n11838 );
or ( n11840 , n5086 , n6110 );
nand ( n11841 , n11839 , n11840 );
nand ( n11842 , n11836 , n11841 );
not ( n11843 , n6113 );
not ( n11844 , n5089 );
or ( n11845 , n11843 , n11844 );
or ( n11846 , n5089 , n6113 );
nand ( n11847 , n11845 , n11846 );
not ( n11848 , n6112 );
not ( n11849 , n5088 );
or ( n11850 , n11848 , n11849 );
or ( n11851 , n5088 , n6112 );
nand ( n11852 , n11850 , n11851 );
nand ( n11853 , n11847 , n11852 );
nor ( n11854 , n11842 , n11853 );
not ( n11855 , n6102 );
not ( n11856 , n5078 );
or ( n11857 , n11855 , n11856 );
or ( n11858 , n5078 , n6102 );
nand ( n11859 , n11857 , n11858 );
not ( n11860 , n6103 );
not ( n11861 , n5079 );
or ( n11862 , n11860 , n11861 );
or ( n11863 , n5079 , n6103 );
nand ( n11864 , n11862 , n11863 );
not ( n11865 , n5080 );
and ( n11866 , n6104 , n11865 );
not ( n11867 , n6104 );
and ( n11868 , n11867 , n5080 );
nor ( n11869 , n11866 , n11868 );
not ( n11870 , n5081 );
and ( n11871 , n6105 , n11870 );
not ( n11872 , n6105 );
and ( n11873 , n11872 , n5081 );
nor ( n11874 , n11871 , n11873 );
nand ( n11875 , n11859 , n11864 , n11869 , n11874 );
not ( n11876 , n11875 );
nand ( n11877 , n11808 , n11831 , n11854 , n11876 );
nor ( n11878 , n11785 , n11877 );
not ( n11879 , n6131 );
not ( n11880 , n5107 );
or ( n11881 , n11879 , n11880 );
or ( n11882 , n5107 , n6131 );
nand ( n11883 , n11881 , n11882 );
not ( n11884 , n6130 );
not ( n11885 , n5106 );
or ( n11886 , n11884 , n11885 );
or ( n11887 , n5106 , n6130 );
nand ( n11888 , n11886 , n11887 );
nand ( n11889 , n11883 , n11888 );
not ( n11890 , n6133 );
not ( n11891 , n5109 );
or ( n11892 , n11890 , n11891 );
or ( n11893 , n5109 , n6133 );
nand ( n11894 , n11892 , n11893 );
not ( n11895 , n6132 );
not ( n11896 , n5108 );
or ( n11897 , n11895 , n11896 );
or ( n11898 , n5108 , n6132 );
nand ( n11899 , n11897 , n11898 );
nand ( n11900 , n11894 , n11899 );
nor ( n11901 , n11889 , n11900 );
not ( n11902 , n5105 );
not ( n11903 , n6129 );
or ( n11904 , n11902 , n11903 );
or ( n11905 , n6129 , n5105 );
nand ( n11906 , n11904 , n11905 );
not ( n11907 , n5104 );
not ( n11908 , n6128 );
or ( n11909 , n11907 , n11908 );
or ( n11910 , n6128 , n5104 );
nand ( n11911 , n11909 , n11910 );
nand ( n11912 , n11906 , n11911 );
not ( n11913 , n6127 );
not ( n11914 , n5103 );
or ( n11915 , n11913 , n11914 );
or ( n11916 , n5103 , n6127 );
nand ( n11917 , n11915 , n11916 );
not ( n11918 , n6126 );
not ( n11919 , n5102 );
or ( n11920 , n11918 , n11919 );
or ( n11921 , n5102 , n6126 );
nand ( n11922 , n11920 , n11921 );
nand ( n11923 , n11917 , n11922 );
nor ( n11924 , n11912 , n11923 );
not ( n11925 , n6123 );
not ( n11926 , n5099 );
or ( n11927 , n11925 , n11926 );
or ( n11928 , n5099 , n6123 );
nand ( n11929 , n11927 , n11928 );
not ( n11930 , n6122 );
not ( n11931 , n5098 );
or ( n11932 , n11930 , n11931 );
or ( n11933 , n5098 , n6122 );
nand ( n11934 , n11932 , n11933 );
nand ( n11935 , n11929 , n11934 );
not ( n11936 , n6125 );
not ( n11937 , n5101 );
or ( n11938 , n11936 , n11937 );
or ( n11939 , n5101 , n6125 );
nand ( n11940 , n11938 , n11939 );
not ( n11941 , n6124 );
not ( n11942 , n5100 );
or ( n11943 , n11941 , n11942 );
or ( n11944 , n5100 , n6124 );
nand ( n11945 , n11943 , n11944 );
nand ( n11946 , n11940 , n11945 );
nor ( n11947 , n11935 , n11946 );
not ( n11948 , n6118 );
not ( n11949 , n5094 );
or ( n11950 , n11948 , n11949 );
or ( n11951 , n5094 , n6118 );
nand ( n11952 , n11950 , n11951 );
not ( n11953 , n6119 );
not ( n11954 , n5095 );
or ( n11955 , n11953 , n11954 );
or ( n11956 , n5095 , n6119 );
nand ( n11957 , n11955 , n11956 );
not ( n11958 , n5096 );
and ( n11959 , n6120 , n11958 );
not ( n11960 , n6120 );
and ( n11961 , n11960 , n5096 );
nor ( n11962 , n11959 , n11961 );
not ( n11963 , n5097 );
and ( n11964 , n6121 , n11963 );
not ( n11965 , n6121 );
and ( n11966 , n11965 , n5097 );
nor ( n11967 , n11964 , n11966 );
nand ( n11968 , n11952 , n11957 , n11962 , n11967 );
not ( n11969 , n11968 );
nand ( n11970 , n11901 , n11924 , n11947 , n11969 );
not ( n11971 , n6136 );
not ( n11972 , n5112 );
or ( n11973 , n11971 , n11972 );
or ( n11974 , n5112 , n6136 );
nand ( n11975 , n11973 , n11974 );
not ( n11976 , n6137 );
not ( n11977 , n5113 );
or ( n11978 , n11976 , n11977 );
or ( n11979 , n5113 , n6137 );
nand ( n11980 , n11978 , n11979 );
not ( n11981 , n6134 );
not ( n11982 , n5110 );
or ( n11983 , n11981 , n11982 );
or ( n11984 , n5110 , n6134 );
nand ( n11985 , n11983 , n11984 );
not ( n11986 , n6135 );
not ( n11987 , n5111 );
or ( n11988 , n11986 , n11987 );
or ( n11989 , n5111 , n6135 );
nand ( n11990 , n11988 , n11989 );
nand ( n11991 , n11975 , n11980 , n11985 , n11990 );
not ( n11992 , n11991 );
not ( n11993 , n6143 );
not ( n11994 , n5119 );
or ( n11995 , n11993 , n11994 );
or ( n11996 , n5119 , n6143 );
nand ( n11997 , n11995 , n11996 );
not ( n11998 , n6142 );
not ( n11999 , n5118 );
or ( n12000 , n11998 , n11999 );
or ( n12001 , n5118 , n6142 );
nand ( n12002 , n12000 , n12001 );
not ( n12003 , n6145 );
not ( n12004 , n5121 );
or ( n12005 , n12003 , n12004 );
or ( n12006 , n5121 , n6145 );
nand ( n12007 , n12005 , n12006 );
not ( n12008 , n6144 );
not ( n12009 , n5120 );
or ( n12010 , n12008 , n12009 );
or ( n12011 , n5120 , n6144 );
nand ( n12012 , n12010 , n12011 );
nand ( n12013 , n11997 , n12002 , n12007 , n12012 );
not ( n12014 , n12013 );
not ( n12015 , n5117 );
and ( n12016 , n6141 , n12015 );
not ( n12017 , n6141 );
and ( n12018 , n12017 , n5117 );
nor ( n12019 , n12016 , n12018 );
not ( n12020 , n5116 );
and ( n12021 , n6140 , n12020 );
not ( n12022 , n6140 );
and ( n12023 , n12022 , n5116 );
nor ( n12024 , n12021 , n12023 );
not ( n12025 , n5115 );
and ( n12026 , n6139 , n12025 );
not ( n12027 , n6139 );
and ( n12028 , n12027 , n5115 );
nor ( n12029 , n12026 , n12028 );
not ( n12030 , n5114 );
and ( n12031 , n6138 , n12030 );
not ( n12032 , n6138 );
and ( n12033 , n12032 , n5114 );
nor ( n12034 , n12031 , n12033 );
nand ( n12035 , n12019 , n12024 , n12029 , n12034 );
not ( n12036 , n12035 );
not ( n12037 , n6146 );
not ( n12038 , n5122 );
or ( n12039 , n12037 , n12038 );
or ( n12040 , n5122 , n6146 );
nand ( n12041 , n12039 , n12040 );
not ( n12042 , n6147 );
and ( n12043 , n5123 , n12042 );
not ( n12044 , n5123 );
and ( n12045 , n12044 , n6147 );
nor ( n12046 , n12043 , n12045 );
not ( n12047 , n6148 );
and ( n12048 , n5124 , n12047 );
not ( n12049 , n5124 );
and ( n12050 , n12049 , n6148 );
nor ( n12051 , n12048 , n12050 );
not ( n12052 , n6149 );
and ( n12053 , n5125 , n12052 );
not ( n12054 , n5125 );
and ( n12055 , n12054 , n6149 );
nor ( n12056 , n12053 , n12055 );
nand ( n12057 , n12041 , n12046 , n12051 , n12056 );
not ( n12058 , n12057 );
nand ( n12059 , n11992 , n12014 , n12036 , n12058 );
nor ( n12060 , n11970 , n12059 );
nand ( n12061 , n11509 , n11694 , n11878 , n12060 );
nor ( n12062 , n11324 , n12061 );
nand ( n12063 , n7621 , n9114 , n10588 , n12062 );
buf ( n12064 , n12063 );
buf ( n12065 , n12064 );
not ( n12066 , n12063 );
buf ( n12067 , n12066 );
buf ( n12068 , n12067 );
endmodule

