//
// Conformal-LEC Version 16.10-d005 ( 21-Apr-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
output n36 , n37 , n38 , n39 , n40 , n41 , n42 ;

wire n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , 
     n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , 
     n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , 
     n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , 
     n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , 
     n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , 
     n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , 
     n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , 
     n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , 
     n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , 
     n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , 
     n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , 
     n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , 
     n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , 
     n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , 
     n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , 
     n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , 
     n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , 
     n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , 
     n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , 
     n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , 
     n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , 
     n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , 
     n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , 
     n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , 
     n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , 
     n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , 
     n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , 
     n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , 
     n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , 
     n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , 
     n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , 
     n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , 
     n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , 
     n425 , n426 , n427 , n428 , n429 , n430 , n431 ;
buf ( n41 , n149 );
buf ( n37 , n235 );
buf ( n36 , n325 );
buf ( n40 , n395 );
buf ( n39 , n412 );
buf ( n42 , n422 );
buf ( n38 , n431 );
buf ( n88 , n18 );
buf ( n89 , n15 );
buf ( n90 , n13 );
buf ( n91 , n9 );
buf ( n92 , n22 );
buf ( n93 , n20 );
buf ( n94 , n29 );
buf ( n95 , n16 );
buf ( n96 , n21 );
buf ( n97 , n23 );
buf ( n98 , n24 );
buf ( n99 , n14 );
buf ( n100 , n6 );
buf ( n101 , n11 );
buf ( n102 , n0 );
buf ( n103 , n7 );
buf ( n104 , n28 );
buf ( n105 , n3 );
buf ( n106 , n1 );
buf ( n107 , n31 );
buf ( n108 , n33 );
buf ( n109 , n12 );
buf ( n110 , n25 );
buf ( n111 , n30 );
buf ( n112 , n27 );
buf ( n113 , n2 );
buf ( n114 , n34 );
buf ( n115 , n35 );
buf ( n116 , n32 );
buf ( n117 , n10 );
buf ( n118 , n8 );
buf ( n119 , n26 );
buf ( n120 , n17 );
buf ( n121 , n4 );
buf ( n122 , n19 );
buf ( n123 , n5 );
not ( n124 , n111 );
nand ( n125 , n124 , n113 );
not ( n126 , n103 );
nand ( n127 , n126 , n105 );
not ( n128 , n119 );
nand ( n129 , n128 , n121 );
not ( n130 , n88 );
nand ( n131 , n130 , n89 );
nand ( n132 , n125 , n127 , n129 , n131 );
not ( n133 , n132 );
not ( n134 , n107 );
nand ( n135 , n134 , n109 );
not ( n136 , n95 );
nand ( n137 , n136 , n97 );
not ( n138 , n91 );
nand ( n139 , n138 , n93 );
nand ( n140 , n135 , n137 , n139 );
not ( n141 , n99 );
nand ( n142 , n141 , n101 );
not ( n143 , n115 );
nand ( n144 , n143 , n117 );
nand ( n145 , n142 , n144 );
nor ( n146 , n140 , n145 );
nand ( n147 , n133 , n146 );
buf ( n148 , n147 );
buf ( n149 , n148 );
not ( n150 , n110 );
not ( n151 , n150 );
not ( n152 , n107 );
nand ( n153 , n152 , n109 );
not ( n154 , n153 );
nand ( n155 , n133 , n146 );
not ( n156 , n155 );
or ( n157 , n154 , n156 );
nand ( n158 , n157 , n109 );
not ( n159 , n158 );
not ( n160 , n159 );
or ( n161 , n151 , n160 );
not ( n162 , n99 );
nand ( n163 , n162 , n101 );
not ( n164 , n163 );
not ( n165 , n155 );
or ( n166 , n164 , n165 );
nand ( n167 , n166 , n101 );
not ( n168 , n167 );
not ( n169 , n102 );
nand ( n170 , n168 , n169 );
nand ( n171 , n161 , n170 );
not ( n172 , n115 );
nand ( n173 , n172 , n117 );
nand ( n174 , n147 , n173 );
not ( n175 , n117 );
nor ( n176 , n175 , n118 );
nand ( n177 , n174 , n176 );
not ( n178 , n91 );
not ( n179 , n95 );
nand ( n180 , n179 , n97 );
not ( n181 , n91 );
nand ( n182 , n181 , n93 );
nand ( n183 , n134 , n109 );
nand ( n184 , n180 , n182 , n183 );
nand ( n185 , n142 , n144 );
nor ( n186 , n184 , n185 );
nand ( n187 , n133 , n186 );
not ( n188 , n187 );
or ( n189 , n178 , n188 );
not ( n190 , n93 );
nor ( n191 , n190 , n94 );
nand ( n192 , n189 , n191 );
not ( n193 , n186 );
not ( n194 , n133 );
or ( n195 , n193 , n194 );
nand ( n196 , n195 , n88 );
not ( n197 , n90 );
and ( n198 , n197 , n89 );
nand ( n199 , n196 , n198 );
nand ( n200 , n177 , n192 , n199 );
nor ( n201 , n171 , n200 );
not ( n202 , n113 );
nor ( n203 , n202 , n114 );
not ( n204 , n203 );
nand ( n205 , n147 , n125 );
not ( n206 , n205 );
or ( n207 , n204 , n206 );
nand ( n208 , n128 , n121 );
not ( n209 , n208 );
not ( n210 , n147 );
or ( n211 , n209 , n210 );
not ( n212 , n121 );
nor ( n213 , n212 , n122 );
nand ( n214 , n211 , n213 );
nand ( n215 , n207 , n214 );
not ( n216 , n97 );
nor ( n217 , n216 , n98 );
not ( n218 , n217 );
nand ( n219 , n187 , n95 );
not ( n220 , n219 );
or ( n221 , n218 , n220 );
buf ( n222 , n127 );
not ( n223 , n222 );
not ( n224 , n187 );
or ( n225 , n223 , n224 );
not ( n226 , n105 );
nor ( n227 , n226 , n106 );
nand ( n228 , n225 , n227 );
nand ( n229 , n221 , n228 );
nor ( n230 , n215 , n229 );
nand ( n231 , n201 , n230 );
not ( n232 , n231 );
not ( n233 , n232 );
buf ( n234 , n233 );
buf ( n235 , n234 );
not ( n236 , n168 );
or ( n237 , n236 , n104 );
not ( n238 , n187 );
not ( n239 , n222 );
or ( n240 , n238 , n239 );
not ( n241 , n105 );
nor ( n242 , n241 , n108 );
nand ( n243 , n240 , n242 );
nand ( n244 , n237 , n243 );
not ( n245 , n97 );
nor ( n246 , n245 , n100 );
not ( n247 , n246 );
not ( n248 , n219 );
or ( n249 , n247 , n248 );
not ( n250 , n89 );
nor ( n251 , n250 , n92 );
nand ( n252 , n196 , n251 );
nand ( n253 , n249 , n252 );
nor ( n254 , n244 , n253 );
not ( n255 , n91 );
not ( n256 , n187 );
or ( n257 , n255 , n256 );
nand ( n258 , n257 , n93 );
not ( n259 , n258 );
not ( n260 , n96 );
and ( n261 , n259 , n260 );
not ( n262 , n173 );
not ( n263 , n147 );
or ( n264 , n262 , n263 );
not ( n265 , n117 );
nor ( n266 , n265 , n120 );
nand ( n267 , n264 , n266 );
not ( n268 , n208 );
not ( n269 , n147 );
or ( n270 , n268 , n269 );
not ( n271 , n121 );
nor ( n272 , n271 , n123 );
nand ( n273 , n270 , n272 );
nand ( n274 , n267 , n273 );
nor ( n275 , n261 , n274 );
not ( n276 , n112 );
nand ( n277 , n159 , n276 );
not ( n278 , n277 );
not ( n279 , n113 );
nor ( n280 , n279 , n116 );
and ( n281 , n205 , n280 );
nor ( n282 , n278 , n281 );
nand ( n283 , n254 , n275 , n282 );
not ( n284 , n283 );
not ( n285 , n232 );
or ( n286 , n284 , n285 );
nor ( n287 , n110 , n158 );
nand ( n288 , n278 , n287 );
not ( n289 , n243 );
not ( n290 , n228 );
and ( n291 , n289 , n290 );
and ( n292 , n280 , n203 );
and ( n293 , n205 , n292 );
nor ( n294 , n291 , n293 );
not ( n295 , n236 );
buf ( n296 , n155 );
and ( n297 , n296 , n163 );
nand ( n298 , n101 , n169 );
nor ( n299 , n297 , n298 );
not ( n300 , n104 );
nand ( n301 , n295 , n299 , n300 );
nand ( n302 , n288 , n294 , n301 );
nand ( n303 , n219 , n217 );
not ( n304 , n303 );
nand ( n305 , n219 , n246 );
not ( n306 , n305 );
and ( n307 , n304 , n306 );
nand ( n308 , n196 , n89 );
nor ( n309 , n308 , n92 );
not ( n310 , n199 );
and ( n311 , n309 , n310 );
nor ( n312 , n307 , n311 );
not ( n313 , n192 );
nor ( n314 , n258 , n96 );
nand ( n315 , n313 , n314 );
nand ( n316 , n174 , n176 );
nor ( n317 , n316 , n267 );
not ( n318 , n317 );
nor ( n319 , n273 , n214 );
not ( n320 , n319 );
nand ( n321 , n312 , n315 , n318 , n320 );
nor ( n322 , n302 , n321 );
nand ( n323 , n286 , n322 );
buf ( n324 , n323 );
buf ( n325 , n324 );
and ( n326 , n323 , n120 );
not ( n327 , n326 );
buf ( n328 , n148 );
nand ( n329 , n328 , n115 );
nand ( n330 , n233 , n118 );
nand ( n331 , n329 , n330 , n117 );
not ( n332 , n331 );
and ( n333 , n327 , n332 );
not ( n334 , n100 );
not ( n335 , n283 );
not ( n336 , n232 );
or ( n337 , n335 , n336 );
nand ( n338 , n337 , n322 );
not ( n339 , n338 );
or ( n340 , n334 , n339 );
and ( n341 , n233 , n98 );
nand ( n342 , n219 , n97 );
nor ( n343 , n341 , n342 );
nand ( n344 , n340 , n343 );
not ( n345 , n344 );
nor ( n346 , n333 , n345 );
not ( n347 , n116 );
not ( n348 , n323 );
or ( n349 , n347 , n348 );
and ( n350 , n328 , n111 );
not ( n351 , n114 );
not ( n352 , n231 );
or ( n353 , n351 , n352 );
nand ( n354 , n353 , n113 );
nor ( n355 , n350 , n354 );
nand ( n356 , n349 , n355 );
nor ( n357 , n93 , n121 );
nand ( n358 , n356 , n357 );
not ( n359 , n112 );
not ( n360 , n338 );
or ( n361 , n359 , n360 );
and ( n362 , n233 , n110 );
nand ( n363 , n328 , n107 );
nand ( n364 , n363 , n109 );
nor ( n365 , n362 , n364 );
nand ( n366 , n361 , n365 );
not ( n367 , n366 );
nor ( n368 , n358 , n367 );
and ( n369 , n233 , n106 );
not ( n370 , n103 );
not ( n371 , n328 );
or ( n372 , n370 , n371 );
nand ( n373 , n372 , n105 );
nor ( n374 , n369 , n373 );
not ( n375 , n374 );
nand ( n376 , n108 , n323 );
not ( n377 , n376 );
or ( n378 , n375 , n377 );
nand ( n379 , n104 , n338 );
and ( n380 , n233 , n102 );
not ( n381 , n99 );
not ( n382 , n328 );
or ( n383 , n381 , n382 );
nand ( n384 , n383 , n101 );
nor ( n385 , n380 , n384 );
nand ( n386 , n379 , n385 );
nand ( n387 , n378 , n386 );
not ( n388 , n387 );
and ( n389 , n346 , n368 , n388 );
and ( n390 , n324 , n92 );
and ( n391 , n233 , n90 );
nor ( n392 , n390 , n391 , n308 );
nor ( n393 , n389 , n392 );
buf ( n394 , n393 );
buf ( n395 , n394 );
nand ( n396 , n376 , n374 );
nand ( n397 , n344 , n396 );
not ( n398 , n397 );
nand ( n399 , n379 , n385 );
not ( n400 , n399 );
and ( n401 , n400 , n344 );
not ( n402 , n96 );
not ( n403 , n338 );
or ( n404 , n402 , n403 );
and ( n405 , n94 , n233 );
nor ( n406 , n405 , n258 );
nand ( n407 , n404 , n406 );
not ( n408 , n407 );
nor ( n409 , n401 , n408 );
nand ( n410 , n398 , n409 );
buf ( n411 , n410 );
buf ( n412 , n411 );
nand ( n413 , n367 , n399 );
or ( n414 , n397 , n413 );
not ( n415 , n387 );
not ( n416 , n356 );
and ( n417 , n415 , n416 );
nand ( n418 , n407 , n344 );
nor ( n419 , n417 , n418 );
nand ( n420 , n414 , n419 );
buf ( n421 , n420 );
buf ( n422 , n421 );
not ( n423 , n326 );
not ( n424 , n331 );
and ( n425 , n423 , n356 , n424 );
and ( n426 , n396 , n367 );
nor ( n427 , n425 , n426 );
or ( n428 , n427 , n345 );
nand ( n429 , n428 , n409 );
buf ( n430 , n429 );
buf ( n431 , n430 );
endmodule

