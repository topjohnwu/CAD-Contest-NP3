//
// Conformal-LEC Version 16.10-d005 ( 21-Apr-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 ;
output n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 ;

wire n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
     n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
     n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , 
     n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , 
     n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , 
     n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , 
     n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , 
     n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
     n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
     n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
     n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
     n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
     n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
     n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
     n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
     n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
     n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
     n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
     n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
     n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
     n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
     n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
     n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
     n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
     n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
     n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
     n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
     n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
     n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
     n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
     n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
     n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , 
     n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , 
     n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
     n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , 
     n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
     n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , 
     n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
     n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
     n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
     n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , 
     n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
     n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
     n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
     n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
     n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
     n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
     n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
     n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
     n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
     n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
     n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
     n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
     n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , 
     n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , 
     n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , 
     n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , 
     n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , 
     n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , 
     n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , 
     n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
     n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , 
     n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , 
     n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , 
     n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , 
     n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , 
     n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , 
     n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , 
     n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , 
     n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , 
     n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , 
     n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , 
     n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , 
     n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , 
     n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , 
     n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
     n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
     n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
     n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
     n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
     n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
     n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
     n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
     n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
     n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
     n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
     n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
     n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
     n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
     n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , 
     n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , 
     n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
     n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , 
     n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , 
     n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , 
     n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , 
     n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , 
     n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , 
     n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , 
     n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , 
     n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
     n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , 
     n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , 
     n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , 
     n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
     n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , 
     n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , 
     n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
     n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , 
     n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , 
     n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , 
     n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , 
     n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , 
     n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , 
     n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , 
     n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , 
     n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , 
     n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , 
     n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , 
     n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , 
     n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , 
     n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , 
     n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , 
     n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , 
     n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , 
     n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , 
     n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
     n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , 
     n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , 
     n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , 
     n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , 
     n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , 
     n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , 
     n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , 
     n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , 
     n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , 
     n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , 
     n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , 
     n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , 
     n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , 
     n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , 
     n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , 
     n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , 
     n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , 
     n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , 
     n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , 
     n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , 
     n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , 
     n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , 
     n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , 
     n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , 
     n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , 
     n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , 
     n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , 
     n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , 
     n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , 
     n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , 
     n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , 
     n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , 
     n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , 
     n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , 
     n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , 
     n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , 
     n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , 
     n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , 
     n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , 
     n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , 
     n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , 
     n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , 
     n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , 
     n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , 
     n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , 
     n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , 
     n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , 
     n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , 
     n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , 
     n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , 
     n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , 
     n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , 
     n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , 
     n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , 
     n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , 
     n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , 
     n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , 
     n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , 
     n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , 
     n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , 
     n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , 
     n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , 
     n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , 
     n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , 
     n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , 
     n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , 
     n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , 
     n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , 
     n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , 
     n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , 
     n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , 
     n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , 
     n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , 
     n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , 
     n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , 
     n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , 
     n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , 
     n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , 
     n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , 
     n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , 
     n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , 
     n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , 
     n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , 
     n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , 
     n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , 
     n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , 
     n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , 
     n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , 
     n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , 
     n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , 
     n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , 
     n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , 
     n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , 
     n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , 
     n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , 
     n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , 
     n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , 
     n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , 
     n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , 
     n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , 
     n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , 
     n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , 
     n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , 
     n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , 
     n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , 
     n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , 
     n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , 
     n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , 
     n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , 
     n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , 
     n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , 
     n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , 
     n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , 
     n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , 
     n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , 
     n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , 
     n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , 
     n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , 
     n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , 
     n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , 
     n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , 
     n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , 
     n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , 
     n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , 
     n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , 
     n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , 
     n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , 
     n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , 
     n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , 
     n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , 
     n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , 
     n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , 
     n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , 
     n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , 
     n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , 
     n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , 
     n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , 
     n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , 
     n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , 
     n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , 
     n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , 
     n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , 
     n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , 
     n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , 
     n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , 
     n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , 
     n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , 
     n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , 
     n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , 
     n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , 
     n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , 
     n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , 
     n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , 
     n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , 
     n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , 
     n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , 
     n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , 
     n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , 
     n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , 
     n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , 
     n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , 
     n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , 
     n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , 
     n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , 
     n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , 
     n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , 
     n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , 
     n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , 
     n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , 
     n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , 
     n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , 
     n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , 
     n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , 
     n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , 
     n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , 
     n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , 
     n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , 
     n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , 
     n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , 
     n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , 
     n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , 
     n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , 
     n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , 
     n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , 
     n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , 
     n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , 
     n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , 
     n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , 
     n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , 
     n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , 
     n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , 
     n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , 
     n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , 
     n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , 
     n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , 
     n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , 
     n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , 
     n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , 
     n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , 
     n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , 
     n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , 
     n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , 
     n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , 
     n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , 
     n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , 
     n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , 
     n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , 
     n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , 
     n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , 
     n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , 
     n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , 
     n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , 
     n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , 
     n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , 
     n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , 
     n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , 
     n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , 
     n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , 
     n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , 
     n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , 
     n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , 
     n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , 
     n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , 
     n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , 
     n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , 
     n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , 
     n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , 
     n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , 
     n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , 
     n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , 
     n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , 
     n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , 
     n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , 
     n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , 
     n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , 
     n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , 
     n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , 
     n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , 
     n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , 
     n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , 
     n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , 
     n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , 
     n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , 
     n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , 
     n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , 
     n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , 
     n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , 
     n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , 
     n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , 
     n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , 
     n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , 
     n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , 
     n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , 
     n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , 
     n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , 
     n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , 
     n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , 
     n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , 
     n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , 
     n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , 
     n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , 
     n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , 
     n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , 
     n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , 
     n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , 
     n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , 
     n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , 
     n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , 
     n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , 
     n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , 
     n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , 
     n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , 
     n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , 
     n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , 
     n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , 
     n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , 
     n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , 
     n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , 
     n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , 
     n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , 
     n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , 
     n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , 
     n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , 
     n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , 
     n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , 
     n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , 
     n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , 
     n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , 
     n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , 
     n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , 
     n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , 
     n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , 
     n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , 
     n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , 
     n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , 
     n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , 
     n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , 
     n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , 
     n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , 
     n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , 
     n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , 
     n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , 
     n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , 
     n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , 
     n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , 
     n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , 
     n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , 
     n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , 
     n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , 
     n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , 
     n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , 
     n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , 
     n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , 
     n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , 
     n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , 
     n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , 
     n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , 
     n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , 
     n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , 
     n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , 
     n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , 
     n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , 
     n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , 
     n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , 
     n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , 
     n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , 
     n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , 
     n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , 
     n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , 
     n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , 
     n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , 
     n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , 
     n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , 
     n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , 
     n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , 
     n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , 
     n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , 
     n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , 
     n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , 
     n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , 
     n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , 
     n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , 
     n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , 
     n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , 
     n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , 
     n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , 
     n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , 
     n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , 
     n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , 
     n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , 
     n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , 
     n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , 
     n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , 
     n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , 
     n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , 
     n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , 
     n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , 
     n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , 
     n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , 
     n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , 
     n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , 
     n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , 
     n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , 
     n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , 
     n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , 
     n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , 
     n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , 
     n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , 
     n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , 
     n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , 
     n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , 
     n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , 
     n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , 
     n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , 
     n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , 
     n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , 
     n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , 
     n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , 
     n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , 
     n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , 
     n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , 
     n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , 
     n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , 
     n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , 
     n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , 
     n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , 
     n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , 
     n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , 
     n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , 
     n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , 
     n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , 
     n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , 
     n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , 
     n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , 
     n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , 
     n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , 
     n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , 
     n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , 
     n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , 
     n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , 
     n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , 
     n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , 
     n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , 
     n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , 
     n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , 
     n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , 
     n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , 
     n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , 
     n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , 
     n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , 
     n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , 
     n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , 
     n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , 
     n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , 
     n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , 
     n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , 
     n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , 
     n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , 
     n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , 
     n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , 
     n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , 
     n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , 
     n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , 
     n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , 
     n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , 
     n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , 
     n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , 
     n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , 
     n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , 
     n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , 
     n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , 
     n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , 
     n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , 
     n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , 
     n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , 
     n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , 
     n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , 
     n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , 
     n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , 
     n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , 
     n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , 
     n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , 
     n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , 
     n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , 
     n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , 
     n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , 
     n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , 
     n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , 
     n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , 
     n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , 
     n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , 
     n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , 
     n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , 
     n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , 
     n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , 
     n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , 
     n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , 
     n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , 
     n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , 
     n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , 
     n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , 
     n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , 
     n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , 
     n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , 
     n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , 
     n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , 
     n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , 
     n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , 
     n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , 
     n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , 
     n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , 
     n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , 
     n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , 
     n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , 
     n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , 
     n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , 
     n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , 
     n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , 
     n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , 
     n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , 
     n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , 
     n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , 
     n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , 
     n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , 
     n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , 
     n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , 
     n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , 
     n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , 
     n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , 
     n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , 
     n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , 
     n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , 
     n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , 
     n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , 
     n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , 
     n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , 
     n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , 
     n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , 
     n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , 
     n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , 
     n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , 
     n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , 
     n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , 
     n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , 
     n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , 
     n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , 
     n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , 
     n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , 
     n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , 
     n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , 
     n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , 
     n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , 
     n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , 
     n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , 
     n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , 
     n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , 
     n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , 
     n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , 
     n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , 
     n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , 
     n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , 
     n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , 
     n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , 
     n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , 
     n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , 
     n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , 
     n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , 
     n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , 
     n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , 
     n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , 
     n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , 
     n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , 
     n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , 
     n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , 
     n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , 
     n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , 
     n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , 
     n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , 
     n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , 
     n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , 
     n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , 
     n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , 
     n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , 
     n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , 
     n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , 
     n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , 
     n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , 
     n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , 
     n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , 
     n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , 
     n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , 
     n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , 
     n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , 
     n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , 
     n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , 
     n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , 
     n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , 
     n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , 
     n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , 
     n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , 
     n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , 
     n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , 
     n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , 
     n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , 
     n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , 
     n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , 
     n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , 
     n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , 
     n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , 
     n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , 
     n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , 
     n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , 
     n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , 
     n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , 
     n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , 
     n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , 
     n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , 
     n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , 
     n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , 
     n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , 
     n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , 
     n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , 
     n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , 
     n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , 
     n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , 
     n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , 
     n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , 
     n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , 
     n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , 
     n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , 
     n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , 
     n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , 
     n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , 
     n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , 
     n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , 
     n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , 
     n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , 
     n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , 
     n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , 
     n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , 
     n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , 
     n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , 
     n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , 
     n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , 
     n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , 
     n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , 
     n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , 
     n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , 
     n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , 
     n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , 
     n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , 
     n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , 
     n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , 
     n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , 
     n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , 
     n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , 
     n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , 
     n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , 
     n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , 
     n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , 
     n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , 
     n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , 
     n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , 
     n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , 
     n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , 
     n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , 
     n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , 
     n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , 
     n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , 
     n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , 
     n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , 
     n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , 
     n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , 
     n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , 
     n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , 
     n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , 
     n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , 
     n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , 
     n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , 
     n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , 
     n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , 
     n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , 
     n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , 
     n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , 
     n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , 
     n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , 
     n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , 
     n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , 
     n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , 
     n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , 
     n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , 
     n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , 
     n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , 
     n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , 
     n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , 
     n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , 
     n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , 
     n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , 
     n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , 
     n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , 
     n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , 
     n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , 
     n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , 
     n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , 
     n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , 
     n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , 
     n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , 
     n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , 
     n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , 
     n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , 
     n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , 
     n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , 
     n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , 
     n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , 
     n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , 
     n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , 
     n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , 
     n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , 
     n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , 
     n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , 
     n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , 
     n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , 
     n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , 
     n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , 
     n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , 
     n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , 
     n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , 
     n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , 
     n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , 
     n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , 
     n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , 
     n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , 
     n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , 
     n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , 
     n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , 
     n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , 
     n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , 
     n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , 
     n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , 
     n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , 
     n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , 
     n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , 
     n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , 
     n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , 
     n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , 
     n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , 
     n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , 
     n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , 
     n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , 
     n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , 
     n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , 
     n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , 
     n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , 
     n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , 
     n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , 
     n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , 
     n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , 
     n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , 
     n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , 
     n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , 
     n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , 
     n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , 
     n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , 
     n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , 
     n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , 
     n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , 
     n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , 
     n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , 
     n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , 
     n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , 
     n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , 
     n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , 
     n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , 
     n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , 
     n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , 
     n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , 
     n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , 
     n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , 
     n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , 
     n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , 
     n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , 
     n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , 
     n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , 
     n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , 
     n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , 
     n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , 
     n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , 
     n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , 
     n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , 
     n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , 
     n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , 
     n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , 
     n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , 
     n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , 
     n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , 
     n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , 
     n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , 
     n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , 
     n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , 
     n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , 
     n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , 
     n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , 
     n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , 
     n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , 
     n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , 
     n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , 
     n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , 
     n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , 
     n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , 
     n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , 
     n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , 
     n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , 
     n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , 
     n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , 
     n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , 
     n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , 
     n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , 
     n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , 
     n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , 
     n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , 
     n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , 
     n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , 
     n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , 
     n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , 
     n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , 
     n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , 
     n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , 
     n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , 
     n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , 
     n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , 
     n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , 
     n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , 
     n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , 
     n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , 
     n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , 
     n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , 
     n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , 
     n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , 
     n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , 
     n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , 
     n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , 
     n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , 
     n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , 
     n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , 
     n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , 
     n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , 
     n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , 
     n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , 
     n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , 
     n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , 
     n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , 
     n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , 
     n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , 
     n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , 
     n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , 
     n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , 
     n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , 
     n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , 
     n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , 
     n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , 
     n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , 
     n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , 
     n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , 
     n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , 
     n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , 
     n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , 
     n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , 
     n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , 
     n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , 
     n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , 
     n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , 
     n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , 
     n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , 
     n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , 
     n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , 
     n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , 
     n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , 
     n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , 
     n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , 
     n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , 
     n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , 
     n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , 
     n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , 
     n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , 
     n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , 
     n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , 
     n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , 
     n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , 
     n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , 
     n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , 
     n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , 
     n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , 
     n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , 
     n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , 
     n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , 
     n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , 
     n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , 
     n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , 
     n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , 
     n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , 
     n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , 
     n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , 
     n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , 
     n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , 
     n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , 
     n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , 
     n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , 
     n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , 
     n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , 
     n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , 
     n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , 
     n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , 
     n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , 
     n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , 
     n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , 
     n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , 
     n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , 
     n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , 
     n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , 
     n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , 
     n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , 
     n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , 
     n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , 
     n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , 
     n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , 
     n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , 
     n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , 
     n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , 
     n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , 
     n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , 
     n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , 
     n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , 
     n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , 
     n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , 
     n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , 
     n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , 
     n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , 
     n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , 
     n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , 
     n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , 
     n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , 
     n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , 
     n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , 
     n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , 
     n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , 
     n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , 
     n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , 
     n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , 
     n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , 
     n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , 
     n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , 
     n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , 
     n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , 
     n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , 
     n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , 
     n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , 
     n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , 
     n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , 
     n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , 
     n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , 
     n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , 
     n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , 
     n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , 
     n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , 
     n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , 
     n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , 
     n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , 
     n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , 
     n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , 
     n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , 
     n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , 
     n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , 
     n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , 
     n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , 
     n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , 
     n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , 
     n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , 
     n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , 
     n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , 
     n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , 
     n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , 
     n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , 
     n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , 
     n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , 
     n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , 
     n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , 
     n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , 
     n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , 
     n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , 
     n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , 
     n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , 
     n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , 
     n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , 
     n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , 
     n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , 
     n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , 
     n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , 
     n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , 
     n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , 
     n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , 
     n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , 
     n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , 
     n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , 
     n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , 
     n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , 
     n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , 
     n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , 
     n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , 
     n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , 
     n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , 
     n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , 
     n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , 
     n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , 
     n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , 
     n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , 
     n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , 
     n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , 
     n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , 
     n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , 
     n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , 
     n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , 
     n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , 
     n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , 
     n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , 
     n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , 
     n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , 
     n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , 
     n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , 
     n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , 
     n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , 
     n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , 
     n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , 
     n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , 
     n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , 
     n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , 
     n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , 
     n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , 
     n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , 
     n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , 
     n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , 
     n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , 
     n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , 
     n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , 
     n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , 
     n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , 
     n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , 
     n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , 
     n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , 
     n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , 
     n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , 
     n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , 
     n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , 
     n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , 
     n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , 
     n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , 
     n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , 
     n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , 
     n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , 
     n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , 
     n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , 
     n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , 
     n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , 
     n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , 
     n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , 
     n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , 
     n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , 
     n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , 
     n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , 
     n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , 
     n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , 
     n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , 
     n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , 
     n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , 
     n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , 
     n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , 
     n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , 
     n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , 
     n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , 
     n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , 
     n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , 
     n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , 
     n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , 
     n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , 
     n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , 
     n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , 
     n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , 
     n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , 
     n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , 
     n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , 
     n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , 
     n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , 
     n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , 
     n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , 
     n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , 
     n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , 
     n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , 
     n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , 
     n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , 
     n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , 
     n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , 
     n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , 
     n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , 
     n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , 
     n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , 
     n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , 
     n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , 
     n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , 
     n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , 
     n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , 
     n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , 
     n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , 
     n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , 
     n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , 
     n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , 
     n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , 
     n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , 
     n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , 
     n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , 
     n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , 
     n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , 
     n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , 
     n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , 
     n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , 
     n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , 
     n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , 
     n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , 
     n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , 
     n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , 
     n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , 
     n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , 
     n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , 
     n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , 
     n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , 
     n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , 
     n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , 
     n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , 
     n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , 
     n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , 
     n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , 
     n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , 
     n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , 
     n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , 
     n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , 
     n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , 
     n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , 
     n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , 
     n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , 
     n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , 
     n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , 
     n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , 
     n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , 
     n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , 
     n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , 
     n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , 
     n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , 
     n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , 
     n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , 
     n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , 
     n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , 
     n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , 
     n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , 
     n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , 
     n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , 
     n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , 
     n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , 
     n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , 
     n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , 
     n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , 
     n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , 
     n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , 
     n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , 
     n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , 
     n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , 
     n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , 
     n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , 
     n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , 
     n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , 
     n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , 
     n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , 
     n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , 
     n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , 
     n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , 
     n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , 
     n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , 
     n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , 
     n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , 
     n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , 
     n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , 
     n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , 
     n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , 
     n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , 
     n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , 
     n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , 
     n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , 
     n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , 
     n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , 
     n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , 
     n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , 
     n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , 
     n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , 
     n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , 
     n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , 
     n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , 
     n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , 
     n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , 
     n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , 
     n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , 
     n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , 
     n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , 
     n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , 
     n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , 
     n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , 
     n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , 
     n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , 
     n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , 
     n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , 
     n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , 
     n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , 
     n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , 
     n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , 
     n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , 
     n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , 
     n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , 
     n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , 
     n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , 
     n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , 
     n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , 
     n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , 
     n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , 
     n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , 
     n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , 
     n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , 
     n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , 
     n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , 
     n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , 
     n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , 
     n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , 
     n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , 
     n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , 
     n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , 
     n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , 
     n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , 
     n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , 
     n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , 
     n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , 
     n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , 
     n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , 
     n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , 
     n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , 
     n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , 
     n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , 
     n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , 
     n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , 
     n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , 
     n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , 
     n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , 
     n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , 
     n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , 
     n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , 
     n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , 
     n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , 
     n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , 
     n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , 
     n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , 
     n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , 
     n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , 
     n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , 
     n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , 
     n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , 
     n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , 
     n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , 
     n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , 
     n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , 
     n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , 
     n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , 
     n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , 
     n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , 
     n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , 
     n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , 
     n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , 
     n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , 
     n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , 
     n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , 
     n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , 
     n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , 
     n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , 
     n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , 
     n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , 
     n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , 
     n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , 
     n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , 
     n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , 
     n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , 
     n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , 
     n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , 
     n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , 
     n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , 
     n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , 
     n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , 
     n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , 
     n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , 
     n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , 
     n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , 
     n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , 
     n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , 
     n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , 
     n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , 
     n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , 
     n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , 
     n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , 
     n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , 
     n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , 
     n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , 
     n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , 
     n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , 
     n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , 
     n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , 
     n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , 
     n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , 
     n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , 
     n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , 
     n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , 
     n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , 
     n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , 
     n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , 
     n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , 
     n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , 
     n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , 
     n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , 
     n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , 
     n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , 
     n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , 
     n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , 
     n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , 
     n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , 
     n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , 
     n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , 
     n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , 
     n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , 
     n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , 
     n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , 
     n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , 
     n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , 
     n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , 
     n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , 
     n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , 
     n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , 
     n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , 
     n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , 
     n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , 
     n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , 
     n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , 
     n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , 
     n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , 
     n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , 
     n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , 
     n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , 
     n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , 
     n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , 
     n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , 
     n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , 
     n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , 
     n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , 
     n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , 
     n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , 
     n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , 
     n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , 
     n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , 
     n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , 
     n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , 
     n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , 
     n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , 
     n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , 
     n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , 
     n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , 
     n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , 
     n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , 
     n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , 
     n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , 
     n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , 
     n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , 
     n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , 
     n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , 
     n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , 
     n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , 
     n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , 
     n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , 
     n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , 
     n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , 
     n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , 
     n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , 
     n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , 
     n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , 
     n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , 
     n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , 
     n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , 
     n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , 
     n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , 
     n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , 
     n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , 
     n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , 
     n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , 
     n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , 
     n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , 
     n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , 
     n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , 
     n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , 
     n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , 
     n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , 
     n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , 
     n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , 
     n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , 
     n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , 
     n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , 
     n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , 
     n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , 
     n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , 
     n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , 
     n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , 
     n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , 
     n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , 
     n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , 
     n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , 
     n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , 
     n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , 
     n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , 
     n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , 
     n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , 
     n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , 
     n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , 
     n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , 
     n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , 
     n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , 
     n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , 
     n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , 
     n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , 
     n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , 
     n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , 
     n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , 
     n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , 
     n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , 
     n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , 
     n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , 
     n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , 
     n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , 
     n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , 
     n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , 
     n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , 
     n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , 
     n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , 
     n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , 
     n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , 
     n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , 
     n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , 
     n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , 
     n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , 
     n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , 
     n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , 
     n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , 
     n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , 
     n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , 
     n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , 
     n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , 
     n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , 
     n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , 
     n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , 
     n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , 
     n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , 
     n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , 
     n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , 
     n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , 
     n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , 
     n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , 
     n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , 
     n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , 
     n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , 
     n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , 
     n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , 
     n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , 
     n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , 
     n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , 
     n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , 
     n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , 
     n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , 
     n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , 
     n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , 
     n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , 
     n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , 
     n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , 
     n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , 
     n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , 
     n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , 
     n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , 
     n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , 
     n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , 
     n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , 
     n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , 
     n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , 
     n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , 
     n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , 
     n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , 
     n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , 
     n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , 
     n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , 
     n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , 
     n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , 
     n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , 
     n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , 
     n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , 
     n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , 
     n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , 
     n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , 
     n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , 
     n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , 
     n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , 
     n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , 
     n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , 
     n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , 
     n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , 
     n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , 
     n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , 
     n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , 
     n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , 
     n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , 
     n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , 
     n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , 
     n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , 
     n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , 
     n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , 
     n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , 
     n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , 
     n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , 
     n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , 
     n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , 
     n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , 
     n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , 
     n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , 
     n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , 
     n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , 
     n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , 
     n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , 
     n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , 
     n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , 
     n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , 
     n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , 
     n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , 
     n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , 
     n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , 
     n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , 
     n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , 
     n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , 
     n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , 
     n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , 
     n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , 
     n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , 
     n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , 
     n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , 
     n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , 
     n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , 
     n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , 
     n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , 
     n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , 
     n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , 
     n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , 
     n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , 
     n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , 
     n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , 
     n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , 
     n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , 
     n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , 
     n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , 
     n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , 
     n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , 
     n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , 
     n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , 
     n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , 
     n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , 
     n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , 
     n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , 
     n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , 
     n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , 
     n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , 
     n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , 
     n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , 
     n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , 
     n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , 
     n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , 
     n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , 
     n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , 
     n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , 
     n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , 
     n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , 
     n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , 
     n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , 
     n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , 
     n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , 
     n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , 
     n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , 
     n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , 
     n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , 
     n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , 
     n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , 
     n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , 
     n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , 
     n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , 
     n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , 
     n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , 
     n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , 
     n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , 
     n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , 
     n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , 
     n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , 
     n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , 
     n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , 
     n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , 
     n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , 
     n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , 
     n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , 
     n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , 
     n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , 
     n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , 
     n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , 
     n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , 
     n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , 
     n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , 
     n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , 
     n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , 
     n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , 
     n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , 
     n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , 
     n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , 
     n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , 
     n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , 
     n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , 
     n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , 
     n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , 
     n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , 
     n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , 
     n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , 
     n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , 
     n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , 
     n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , 
     n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , 
     n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , 
     n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , 
     n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , 
     n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , 
     n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , 
     n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , 
     n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , 
     n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , 
     n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , 
     n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , 
     n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , 
     n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , 
     n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , 
     n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , 
     n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , 
     n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , 
     n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , 
     n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , 
     n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , 
     n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , 
     n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , 
     n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , 
     n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , 
     n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , 
     n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , 
     n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , 
     n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , 
     n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , 
     n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , 
     n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , 
     n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , 
     n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , 
     n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , 
     n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , 
     n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , 
     n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , 
     n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , 
     n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , 
     n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , 
     n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , 
     n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , 
     n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , 
     n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , 
     n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , 
     n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , 
     n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , 
     n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , 
     n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , 
     n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , 
     n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , 
     n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , 
     n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , 
     n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , 
     n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , 
     n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , 
     n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , 
     n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , 
     n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , 
     n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , 
     n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , 
     n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , 
     n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , 
     n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , 
     n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , 
     n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , 
     n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , 
     n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , 
     n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , 
     n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , 
     n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , 
     n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , 
     n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , 
     n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , 
     n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , 
     n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , 
     n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , 
     n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , 
     n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , 
     n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , 
     n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , 
     n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , 
     n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , 
     n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , 
     n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , 
     n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , 
     n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , 
     n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , 
     n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , 
     n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , 
     n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , 
     n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , 
     n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , 
     n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , 
     n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , 
     n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , 
     n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , 
     n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , 
     n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , 
     n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , 
     n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , 
     n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , 
     n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , 
     n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , 
     n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , 
     n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , 
     n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , 
     n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , 
     n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , 
     n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , 
     n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , 
     n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , 
     n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , 
     n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , 
     n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , 
     n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , 
     n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , 
     n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , 
     n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , 
     n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , 
     n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , 
     n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , 
     n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , 
     n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , 
     n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , 
     n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , 
     n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , 
     n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , 
     n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , 
     n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , 
     n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , 
     n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , 
     n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , 
     n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , 
     n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , 
     n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , 
     n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , 
     n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , 
     n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , 
     n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , 
     n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , 
     n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , 
     n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , 
     n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , 
     n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , 
     n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , 
     n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , 
     n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , 
     n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , 
     n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , 
     n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , 
     n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , 
     n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , 
     n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , 
     n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , 
     n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , 
     n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , 
     n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , 
     n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , 
     n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , 
     n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , 
     n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , 
     n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , 
     n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , 
     n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , 
     n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , 
     n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , 
     n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , 
     n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , 
     n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , 
     n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , 
     n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , 
     n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , 
     n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , 
     n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , 
     n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , 
     n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , 
     n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , 
     n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , 
     n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , 
     n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , 
     n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , 
     n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , 
     n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , 
     n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , 
     n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , 
     n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , 
     n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , 
     n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , 
     n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , 
     n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , 
     n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , 
     n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , 
     n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , 
     n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , 
     n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , 
     n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , 
     n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , 
     n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , 
     n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , 
     n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , 
     n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , 
     n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , 
     n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , 
     n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , 
     n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , 
     n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , 
     n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , 
     n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , 
     n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , 
     n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , 
     n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , 
     n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , 
     n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , 
     n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , 
     n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , 
     n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , 
     n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , 
     n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , 
     n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , 
     n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , 
     n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , 
     n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , 
     n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , 
     n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , 
     n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , 
     n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , 
     n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , 
     n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , 
     n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , 
     n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , 
     n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , 
     n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , 
     n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , 
     n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , 
     n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , 
     n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , 
     n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , 
     n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , 
     n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , 
     n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , 
     n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , 
     n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , 
     n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , 
     n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , 
     n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , 
     n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , 
     n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , 
     n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , 
     n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , 
     n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , 
     n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , 
     n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , 
     n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , 
     n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , 
     n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , 
     n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , 
     n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , 
     n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , 
     n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , 
     n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , 
     n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , 
     n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , 
     n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , 
     n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , 
     n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , 
     n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , 
     n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , 
     n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , 
     n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , 
     n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , 
     n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , 
     n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , 
     n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , 
     n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , 
     n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , 
     n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , 
     n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , 
     n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , 
     n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , 
     n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , 
     n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , 
     n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , 
     n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , 
     n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , 
     n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , 
     n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , 
     n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , 
     n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , 
     n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , 
     n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , 
     n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , 
     n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , 
     n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , 
     n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , 
     n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , 
     n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , 
     n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , 
     n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , 
     n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , 
     n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , 
     n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , 
     n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , 
     n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , 
     n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , 
     n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , 
     n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , 
     n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , 
     n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , 
     n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , 
     n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , 
     n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , 
     n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , 
     n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , 
     n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , 
     n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , 
     n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , 
     n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , 
     n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , 
     n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , 
     n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , 
     n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , 
     n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , 
     n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , 
     n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , 
     n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , 
     n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , 
     n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , 
     n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , 
     n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , 
     n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , 
     n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , 
     n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , 
     n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , 
     n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , 
     n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , 
     n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , 
     n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , 
     n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , 
     n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , 
     n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , 
     n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , 
     n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , 
     n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , 
     n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , 
     n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , 
     n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , 
     n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , 
     n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , 
     n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , 
     n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , 
     n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , 
     n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , 
     n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , 
     n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , 
     n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , 
     n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , 
     n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , 
     n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , 
     n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , 
     n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , 
     n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , 
     n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , 
     n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , 
     n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , 
     n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , 
     n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , 
     n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , 
     n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , 
     n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , 
     n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , 
     n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , 
     n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , 
     n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , 
     n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , 
     n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , 
     n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , 
     n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , 
     n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , 
     n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , 
     n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , 
     n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , 
     n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , 
     n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , 
     n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , 
     n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , 
     n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , 
     n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , 
     n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , 
     n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , 
     n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , 
     n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , 
     n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , 
     n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , 
     n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , 
     n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , 
     n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , 
     n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , 
     n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , 
     n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , 
     n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , 
     n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , 
     n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , 
     n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , 
     n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , 
     n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , 
     n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , 
     n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , 
     n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , 
     n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , 
     n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , 
     n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , 
     n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , 
     n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , 
     n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , 
     n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , 
     n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , 
     n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , 
     n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , 
     n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , 
     n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , 
     n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , 
     n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , 
     n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , 
     n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , 
     n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , 
     n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , 
     n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , 
     n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , 
     n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , 
     n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , 
     n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , 
     n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , 
     n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , 
     n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , 
     n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , 
     n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , 
     n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , 
     n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , 
     n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , 
     n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , 
     n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , 
     n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , 
     n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , 
     n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , 
     n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , 
     n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , 
     n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , 
     n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , 
     n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , 
     n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , 
     n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , 
     n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , 
     n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , 
     n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , 
     n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , 
     n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , 
     n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , 
     n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , 
     n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , 
     n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , 
     n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , 
     n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , 
     n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , 
     n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , 
     n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , 
     n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , 
     n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , 
     n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , 
     n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , 
     n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , 
     n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , 
     n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , 
     n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , 
     n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , 
     n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , 
     n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , 
     n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , 
     n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , 
     n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , 
     n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , 
     n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , 
     n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , 
     n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , 
     n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , 
     n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , 
     n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , 
     n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , 
     n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , 
     n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , 
     n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , 
     n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , 
     n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , 
     n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , 
     n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , 
     n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , 
     n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , 
     n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , 
     n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , 
     n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , 
     n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , 
     n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , 
     n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , 
     n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , 
     n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , 
     n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , 
     n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , 
     n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , 
     n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , 
     n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , 
     n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , 
     n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , 
     n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , 
     n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , 
     n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , 
     n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , 
     n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , 
     n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , 
     n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , 
     n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , 
     n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , 
     n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , 
     n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , 
     n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , 
     n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , 
     n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , 
     n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , 
     n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , 
     n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , 
     n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , 
     n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , 
     n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , 
     n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , 
     n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , 
     n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , 
     n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , 
     n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , 
     n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , 
     n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , 
     n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , 
     n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , 
     n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , 
     n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , 
     n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , 
     n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , 
     n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , 
     n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , 
     n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , 
     n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , 
     n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , 
     n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , 
     n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , 
     n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , 
     n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , 
     n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , 
     n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , 
     n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , 
     n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , 
     n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , 
     n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , 
     n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , 
     n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , 
     n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , 
     n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , 
     n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , 
     n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , 
     n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , 
     n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , 
     n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , 
     n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , 
     n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , 
     n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , 
     n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , 
     n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , 
     n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , 
     n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , 
     n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , 
     n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , 
     n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , 
     n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , 
     n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , 
     n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , 
     n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , 
     n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , 
     n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , 
     n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , 
     n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , 
     n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , 
     n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , 
     n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , 
     n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , 
     n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , 
     n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , 
     n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , 
     n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , 
     n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , 
     n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , 
     n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , 
     n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , 
     n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , 
     n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , 
     n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , 
     n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , 
     n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , 
     n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , 
     n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , 
     n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , 
     n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , 
     n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , 
     n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , 
     n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , 
     n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , 
     n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , 
     n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , 
     n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , 
     n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , 
     n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , 
     n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , 
     n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , 
     n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , 
     n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , 
     n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , 
     n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , 
     n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , 
     n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , 
     n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , 
     n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , 
     n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , 
     n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , 
     n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , 
     n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , 
     n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , 
     n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , 
     n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , 
     n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , 
     n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , 
     n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , 
     n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , 
     n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , 
     n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , 
     n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , 
     n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , 
     n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , 
     n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , 
     n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , 
     n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , 
     n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , 
     n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , 
     n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , 
     n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , 
     n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , 
     n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , 
     n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , 
     n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , 
     n28151 ;
buf ( n2160 , n13359 );
buf ( n2158 , n17817 );
buf ( n2152 , n20981 );
buf ( n2157 , n21742 );
buf ( n2156 , n23073 );
buf ( n2151 , n24731 );
buf ( n2153 , n25632 );
buf ( n2155 , n26703 );
buf ( n2154 , n27224 );
buf ( n2159 , n28151 );
buf ( n4324 , n387 );
buf ( n4325 , n1678 );
buf ( n4326 , n137 );
buf ( n4327 , n1077 );
buf ( n4328 , n52 );
buf ( n4329 , n426 );
buf ( n4330 , n2024 );
buf ( n4331 , n1146 );
buf ( n4332 , n1897 );
buf ( n4333 , n1333 );
buf ( n4334 , n280 );
buf ( n4335 , n848 );
buf ( n4336 , n824 );
buf ( n4337 , n1122 );
buf ( n4338 , n2028 );
buf ( n4339 , n735 );
buf ( n4340 , n1217 );
buf ( n4341 , n394 );
buf ( n4342 , n1043 );
buf ( n4343 , n1880 );
buf ( n4344 , n980 );
buf ( n4345 , n694 );
buf ( n4346 , n1679 );
buf ( n4347 , n350 );
buf ( n4348 , n294 );
buf ( n4349 , n1647 );
buf ( n4350 , n871 );
buf ( n4351 , n404 );
buf ( n4352 , n894 );
buf ( n4353 , n1789 );
buf ( n4354 , n890 );
buf ( n4355 , n149 );
buf ( n4356 , n6 );
buf ( n4357 , n1412 );
buf ( n4358 , n859 );
buf ( n4359 , n2016 );
buf ( n4360 , n1300 );
buf ( n4361 , n616 );
buf ( n4362 , n508 );
buf ( n4363 , n102 );
buf ( n4364 , n1596 );
buf ( n4365 , n567 );
buf ( n4366 , n1640 );
buf ( n4367 , n303 );
buf ( n4368 , n2 );
buf ( n4369 , n2083 );
buf ( n4370 , n1219 );
buf ( n4371 , n115 );
buf ( n4372 , n249 );
buf ( n4373 , n407 );
buf ( n4374 , n1616 );
buf ( n4375 , n572 );
buf ( n4376 , n17 );
buf ( n4377 , n1461 );
buf ( n4378 , n401 );
buf ( n4379 , n71 );
buf ( n4380 , n719 );
buf ( n4381 , n136 );
buf ( n4382 , n8 );
buf ( n4383 , n1029 );
buf ( n4384 , n1358 );
buf ( n4385 , n13 );
buf ( n4386 , n677 );
buf ( n4387 , n997 );
buf ( n4388 , n1262 );
buf ( n4389 , n448 );
buf ( n4390 , n857 );
buf ( n4391 , n465 );
buf ( n4392 , n1574 );
buf ( n4393 , n1697 );
buf ( n4394 , n1685 );
buf ( n4395 , n1735 );
buf ( n4396 , n1368 );
buf ( n4397 , n1176 );
buf ( n4398 , n340 );
buf ( n4399 , n364 );
buf ( n4400 , n1282 );
buf ( n4401 , n1500 );
buf ( n4402 , n543 );
buf ( n4403 , n100 );
buf ( n4404 , n403 );
buf ( n4405 , n81 );
buf ( n4406 , n774 );
buf ( n4407 , n98 );
buf ( n4408 , n510 );
buf ( n4409 , n829 );
buf ( n4410 , n1795 );
buf ( n4411 , n615 );
buf ( n4412 , n582 );
buf ( n4413 , n158 );
buf ( n4414 , n964 );
buf ( n4415 , n909 );
buf ( n4416 , n1786 );
buf ( n4417 , n91 );
buf ( n4418 , n1297 );
buf ( n4419 , n689 );
buf ( n4420 , n1359 );
buf ( n4421 , n2087 );
buf ( n4422 , n1086 );
buf ( n4423 , n1209 );
buf ( n4424 , n1452 );
buf ( n4425 , n1650 );
buf ( n4426 , n1486 );
buf ( n4427 , n936 );
buf ( n4428 , n736 );
buf ( n4429 , n1932 );
buf ( n4430 , n1603 );
buf ( n4431 , n1166 );
buf ( n4432 , n1095 );
buf ( n4433 , n1347 );
buf ( n4434 , n18 );
buf ( n4435 , n287 );
buf ( n4436 , n1249 );
buf ( n4437 , n880 );
buf ( n4438 , n29 );
buf ( n4439 , n1075 );
buf ( n4440 , n1831 );
buf ( n4441 , n1134 );
buf ( n4442 , n1482 );
buf ( n4443 , n682 );
buf ( n4444 , n1658 );
buf ( n4445 , n32 );
buf ( n4446 , n1076 );
buf ( n4447 , n211 );
buf ( n4448 , n2143 );
buf ( n4449 , n799 );
buf ( n4450 , n786 );
buf ( n4451 , n146 );
buf ( n4452 , n1722 );
buf ( n4453 , n488 );
buf ( n4454 , n1406 );
buf ( n4455 , n1799 );
buf ( n4456 , n2082 );
buf ( n4457 , n492 );
buf ( n4458 , n557 );
buf ( n4459 , n1885 );
buf ( n4460 , n2025 );
buf ( n4461 , n1607 );
buf ( n4462 , n1884 );
buf ( n4463 , n116 );
buf ( n4464 , n182 );
buf ( n4465 , n1054 );
buf ( n4466 , n670 );
buf ( n4467 , n297 );
buf ( n4468 , n120 );
buf ( n4469 , n1206 );
buf ( n4470 , n1531 );
buf ( n4471 , n2102 );
buf ( n4472 , n1959 );
buf ( n4473 , n49 );
buf ( n4474 , n1132 );
buf ( n4475 , n180 );
buf ( n4476 , n691 );
buf ( n4477 , n724 );
buf ( n4478 , n1576 );
buf ( n4479 , n1979 );
buf ( n4480 , n1097 );
buf ( n4481 , n150 );
buf ( n4482 , n326 );
buf ( n4483 , n1048 );
buf ( n4484 , n1775 );
buf ( n4485 , n633 );
buf ( n4486 , n377 );
buf ( n4487 , n529 );
buf ( n4488 , n1085 );
buf ( n4489 , n1674 );
buf ( n4490 , n1727 );
buf ( n4491 , n370 );
buf ( n4492 , n1879 );
buf ( n4493 , n701 );
buf ( n4494 , n1992 );
buf ( n4495 , n507 );
buf ( n4496 , n676 );
buf ( n4497 , n173 );
buf ( n4498 , n1568 );
buf ( n4499 , n1600 );
buf ( n4500 , n707 );
buf ( n4501 , n798 );
buf ( n4502 , n1150 );
buf ( n4503 , n470 );
buf ( n4504 , n2091 );
buf ( n4505 , n524 );
buf ( n4506 , n1394 );
buf ( n4507 , n1337 );
buf ( n4508 , n53 );
buf ( n4509 , n395 );
buf ( n4510 , n1652 );
buf ( n4511 , n477 );
buf ( n4512 , n1275 );
buf ( n4513 , n341 );
buf ( n4514 , n184 );
buf ( n4515 , n673 );
buf ( n4516 , n509 );
buf ( n4517 , n396 );
buf ( n4518 , n1100 );
buf ( n4519 , n1309 );
buf ( n4520 , n708 );
buf ( n4521 , n1222 );
buf ( n4522 , n1349 );
buf ( n4523 , n1039 );
buf ( n4524 , n70 );
buf ( n4525 , n261 );
buf ( n4526 , n1202 );
buf ( n4527 , n808 );
buf ( n4528 , n1157 );
buf ( n4529 , n84 );
buf ( n4530 , n769 );
buf ( n4531 , n776 );
buf ( n4532 , n90 );
buf ( n4533 , n992 );
buf ( n4534 , n1191 );
buf ( n4535 , n1400 );
buf ( n4536 , n1824 );
buf ( n4537 , n117 );
buf ( n4538 , n1464 );
buf ( n4539 , n929 );
buf ( n4540 , n1882 );
buf ( n4541 , n1378 );
buf ( n4542 , n1285 );
buf ( n4543 , n1105 );
buf ( n4544 , n1614 );
buf ( n4545 , n2075 );
buf ( n4546 , n667 );
buf ( n4547 , n960 );
buf ( n4548 , n578 );
buf ( n4549 , n1754 );
buf ( n4550 , n1881 );
buf ( n4551 , n245 );
buf ( n4552 , n1872 );
buf ( n4553 , n837 );
buf ( n4554 , n399 );
buf ( n4555 , n503 );
buf ( n4556 , n143 );
buf ( n4557 , n1205 );
buf ( n4558 , n1371 );
buf ( n4559 , n422 );
buf ( n4560 , n1721 );
buf ( n4561 , n398 );
buf ( n4562 , n331 );
buf ( n4563 , n830 );
buf ( n4564 , n1170 );
buf ( n4565 , n1855 );
buf ( n4566 , n1023 );
buf ( n4567 , n1380 );
buf ( n4568 , n1668 );
buf ( n4569 , n63 );
buf ( n4570 , n1033 );
buf ( n4571 , n2049 );
buf ( n4572 , n780 );
buf ( n4573 , n1955 );
buf ( n4574 , n74 );
buf ( n4575 , n218 );
buf ( n4576 , n1495 );
buf ( n4577 , n1283 );
buf ( n4578 , n660 );
buf ( n4579 , n322 );
buf ( n4580 , n449 );
buf ( n4581 , n35 );
buf ( n4582 , n271 );
buf ( n4583 , n2040 );
buf ( n4584 , n505 );
buf ( n4585 , n1562 );
buf ( n4586 , n906 );
buf ( n4587 , n1171 );
buf ( n4588 , n378 );
buf ( n4589 , n28 );
buf ( n4590 , n1370 );
buf ( n4591 , n659 );
buf ( n4592 , n983 );
buf ( n4593 , n1733 );
buf ( n4594 , n675 );
buf ( n4595 , n821 );
buf ( n4596 , n114 );
buf ( n4597 , n1526 );
buf ( n4598 , n1611 );
buf ( n4599 , n1505 );
buf ( n4600 , n496 );
buf ( n4601 , n2071 );
buf ( n4602 , n812 );
buf ( n4603 , n2029 );
buf ( n4604 , n307 );
buf ( n4605 , n931 );
buf ( n4606 , n1090 );
buf ( n4607 , n282 );
buf ( n4608 , n683 );
buf ( n4609 , n889 );
buf ( n4610 , n1318 );
buf ( n4611 , n316 );
buf ( n4612 , n1063 );
buf ( n4613 , n990 );
buf ( n4614 , n167 );
buf ( n4615 , n1962 );
buf ( n4616 , n33 );
buf ( n4617 , n2148 );
buf ( n4618 , n1492 );
buf ( n4619 , n1755 );
buf ( n4620 , n1409 );
buf ( n4621 , n487 );
buf ( n4622 , n699 );
buf ( n4623 , n1985 );
buf ( n4624 , n816 );
buf ( n4625 , n1136 );
buf ( n4626 , n686 );
buf ( n4627 , n1550 );
buf ( n4628 , n1145 );
buf ( n4629 , n1812 );
buf ( n4630 , n214 );
buf ( n4631 , n1952 );
buf ( n4632 , n954 );
buf ( n4633 , n1776 );
buf ( n4634 , n904 );
buf ( n4635 , n942 );
buf ( n4636 , n2013 );
buf ( n4637 , n1391 );
buf ( n4638 , n1625 );
buf ( n4639 , n782 );
buf ( n4640 , n1021 );
buf ( n4641 , n372 );
buf ( n4642 , n1228 );
buf ( n4643 , n730 );
buf ( n4644 , n762 );
buf ( n4645 , n1970 );
buf ( n4646 , n1488 );
buf ( n4647 , n225 );
buf ( n4648 , n1529 );
buf ( n4649 , n1620 );
buf ( n4650 , n1268 );
buf ( n4651 , n2109 );
buf ( n4652 , n371 );
buf ( n4653 , n1348 );
buf ( n4654 , n725 );
buf ( n4655 , n1737 );
buf ( n4656 , n1621 );
buf ( n4657 , n1714 );
buf ( n4658 , n832 );
buf ( n4659 , n662 );
buf ( n4660 , n775 );
buf ( n4661 , n1762 );
buf ( n4662 , n384 );
buf ( n4663 , n641 );
buf ( n4664 , n632 );
buf ( n4665 , n1973 );
buf ( n4666 , n1846 );
buf ( n4667 , n484 );
buf ( n4668 , n1656 );
buf ( n4669 , n1689 );
buf ( n4670 , n1525 );
buf ( n4671 , n882 );
buf ( n4672 , n986 );
buf ( n4673 , n688 );
buf ( n4674 , n1728 );
buf ( n4675 , n860 );
buf ( n4676 , n206 );
buf ( n4677 , n171 );
buf ( n4678 , n1458 );
buf ( n4679 , n362 );
buf ( n4680 , n1372 );
buf ( n4681 , n363 );
buf ( n4682 , n760 );
buf ( n4683 , n666 );
buf ( n4684 , n631 );
buf ( n4685 , n2095 );
buf ( n4686 , n1852 );
buf ( n4687 , n994 );
buf ( n4688 , n77 );
buf ( n4689 , n2100 );
buf ( n4690 , n1366 );
buf ( n4691 , n1017 );
buf ( n4692 , n335 );
buf ( n4693 , n1137 );
buf ( n4694 , n841 );
buf ( n4695 , n2026 );
buf ( n4696 , n984 );
buf ( n4697 , n2015 );
buf ( n4698 , n1314 );
buf ( n4699 , n365 );
buf ( n4700 , n648 );
buf ( n4701 , n553 );
buf ( n4702 , n1854 );
buf ( n4703 , n134 );
buf ( n4704 , n1538 );
buf ( n4705 , n1585 );
buf ( n4706 , n2123 );
buf ( n4707 , n1207 );
buf ( n4708 , n926 );
buf ( n4709 , n621 );
buf ( n4710 , n976 );
buf ( n4711 , n958 );
buf ( n4712 , n518 );
buf ( n4713 , n1379 );
buf ( n4714 , n288 );
buf ( n4715 , n1565 );
buf ( n4716 , n1436 );
buf ( n4717 , n636 );
buf ( n4718 , n1045 );
buf ( n4719 , n2022 );
buf ( n4720 , n1618 );
buf ( n4721 , n2090 );
buf ( n4722 , n456 );
buf ( n4723 , n629 );
buf ( n4724 , n1290 );
buf ( n4725 , n2031 );
buf ( n4726 , n558 );
buf ( n4727 , n560 );
buf ( n4728 , n1947 );
buf ( n4729 , n1287 );
buf ( n4730 , n1354 );
buf ( n4731 , n169 );
buf ( n4732 , n1582 );
buf ( n4733 , n2072 );
buf ( n4734 , n907 );
buf ( n4735 , n1558 );
buf ( n4736 , n272 );
buf ( n4737 , n1951 );
buf ( n4738 , n247 );
buf ( n4739 , n1001 );
buf ( n4740 , n1158 );
buf ( n4741 , n2020 );
buf ( n4742 , n205 );
buf ( n4743 , n207 );
buf ( n4744 , n908 );
buf ( n4745 , n1459 );
buf ( n4746 , n468 );
buf ( n4747 , n1633 );
buf ( n4748 , n577 );
buf ( n4749 , n191 );
buf ( n4750 , n1922 );
buf ( n4751 , n59 );
buf ( n4752 , n1113 );
buf ( n4753 , n1426 );
buf ( n4754 , n687 );
buf ( n4755 , n1351 );
buf ( n4756 , n1109 );
buf ( n4757 , n924 );
buf ( n4758 , n379 );
buf ( n4759 , n765 );
buf ( n4760 , n1042 );
buf ( n4761 , n2027 );
buf ( n4762 , n1225 );
buf ( n4763 , n68 );
buf ( n4764 , n915 );
buf ( n4765 , n2036 );
buf ( n4766 , n1820 );
buf ( n4767 , n1629 );
buf ( n4768 , n1630 );
buf ( n4769 , n1752 );
buf ( n4770 , n181 );
buf ( n4771 , n437 );
buf ( n4772 , n1323 );
buf ( n4773 , n834 );
buf ( n4774 , n1553 );
buf ( n4775 , n1156 );
buf ( n4776 , n820 );
buf ( n4777 , n2117 );
buf ( n4778 , n1455 );
buf ( n4779 , n825 );
buf ( n4780 , n1385 );
buf ( n4781 , n2058 );
buf ( n4782 , n1057 );
buf ( n4783 , n1875 );
buf ( n4784 , n1481 );
buf ( n4785 , n1356 );
buf ( n4786 , n727 );
buf ( n4787 , n1164 );
buf ( n4788 , n1663 );
buf ( n4789 , n988 );
buf ( n4790 , n1334 );
buf ( n4791 , n232 );
buf ( n4792 , n1696 );
buf ( n4793 , n127 );
buf ( n4794 , n1512 );
buf ( n4795 , n746 );
buf ( n4796 , n1773 );
buf ( n4797 , n1528 );
buf ( n4798 , n1294 );
buf ( n4799 , n594 );
buf ( n4800 , n903 );
buf ( n4801 , n1948 );
buf ( n4802 , n1027 );
buf ( n4803 , n298 );
buf ( n4804 , n2066 );
buf ( n4805 , n131 );
buf ( n4806 , n1676 );
buf ( n4807 , n1816 );
buf ( n4808 , n1592 );
buf ( n4809 , n886 );
buf ( n4810 , n1507 );
buf ( n4811 , n2077 );
buf ( n4812 , n1401 );
buf ( n4813 , n1871 );
buf ( n4814 , n1231 );
buf ( n4815 , n1088 );
buf ( n4816 , n1240 );
buf ( n4817 , n1811 );
buf ( n4818 , n1431 );
buf ( n4819 , n917 );
buf ( n4820 , n1587 );
buf ( n4821 , n1913 );
buf ( n4822 , n1230 );
buf ( n4823 , n1093 );
buf ( n4824 , n34 );
buf ( n4825 , n772 );
buf ( n4826 , n2039 );
buf ( n4827 , n1950 );
buf ( n4828 , n1965 );
buf ( n4829 , n1129 );
buf ( n4830 , n1670 );
buf ( n4831 , n1648 );
buf ( n4832 , n1916 );
buf ( n4833 , n1660 );
buf ( n4834 , n1067 );
buf ( n4835 , n749 );
buf ( n4836 , n1544 );
buf ( n4837 , n1794 );
buf ( n4838 , n1848 );
buf ( n4839 , n1987 );
buf ( n4840 , n19 );
buf ( n4841 , n1866 );
buf ( n4842 , n2068 );
buf ( n4843 , n2018 );
buf ( n4844 , n2103 );
buf ( n4845 , n1243 );
buf ( n4846 , n1098 );
buf ( n4847 , n412 );
buf ( n4848 , n172 );
buf ( n4849 , n121 );
buf ( n4850 , n1766 );
buf ( n4851 , n87 );
buf ( n4852 , n2063 );
buf ( n4853 , n728 );
buf ( n4854 , n1244 );
buf ( n4855 , n563 );
buf ( n4856 , n1059 );
buf ( n4857 , n76 );
buf ( n4858 , n1694 );
buf ( n4859 , n1998 );
buf ( n4860 , n1167 );
buf ( n4861 , n123 );
buf ( n4862 , n101 );
buf ( n4863 , n1609 );
buf ( n4864 , n584 );
buf ( n4865 , n1849 );
buf ( n4866 , n354 );
buf ( n4867 , n777 );
buf ( n4868 , n406 );
buf ( n4869 , n2107 );
buf ( n4870 , n2142 );
buf ( n4871 , n822 );
buf ( n4872 , n490 );
buf ( n4873 , n2053 );
buf ( n4874 , n2076 );
buf ( n4875 , n846 );
buf ( n4876 , n1019 );
buf ( n4877 , n1858 );
buf ( n4878 , n1099 );
buf ( n4879 , n1800 );
buf ( n4880 , n1430 );
buf ( n4881 , n2114 );
buf ( n4882 , n1277 );
buf ( n4883 , n1997 );
buf ( n4884 , n1447 );
buf ( n4885 , n1454 );
buf ( n4886 , n1612 );
buf ( n4887 , n1691 );
buf ( n4888 , n302 );
buf ( n4889 , n2124 );
buf ( n4890 , n733 );
buf ( n4891 , n2074 );
buf ( n4892 , n571 );
buf ( n4893 , n1438 );
buf ( n4894 , n818 );
buf ( n4895 , n548 );
buf ( n4896 , n498 );
buf ( n4897 , n2005 );
buf ( n4898 , n62 );
buf ( n4899 , n201 );
buf ( n4900 , n1506 );
buf ( n4901 , n732 );
buf ( n4902 , n528 );
buf ( n4903 , n933 );
buf ( n4904 , n586 );
buf ( n4905 , n1966 );
buf ( n4906 , n1295 );
buf ( n4907 , n588 );
buf ( n4908 , n2136 );
buf ( n4909 , n262 );
buf ( n4910 , n2135 );
buf ( n4911 , n423 );
buf ( n4912 , n1725 );
buf ( n4913 , n539 );
buf ( n4914 , n1623 );
buf ( n4915 , n1497 );
buf ( n4916 , n1140 );
buf ( n4917 , n944 );
buf ( n4918 , n1608 );
buf ( n4919 , n140 );
buf ( n4920 , n221 );
buf ( n4921 , n1102 );
buf ( n4922 , n1271 );
buf ( n4923 , n312 );
buf ( n4924 , n635 );
buf ( n4925 , n853 );
buf ( n4926 , n1357 );
buf ( n4927 , n1269 );
buf ( n4928 , n1024 );
buf ( n4929 , n30 );
buf ( n4930 , n828 );
buf ( n4931 , n1473 );
buf ( n4932 , n705 );
buf ( n4933 , n436 );
buf ( n4934 , n2011 );
buf ( n4935 , n1716 );
buf ( n4936 , n946 );
buf ( n4937 , n1200 );
buf ( n4938 , n1825 );
buf ( n4939 , n1583 );
buf ( n4940 , n1873 );
buf ( n4941 , n601 );
buf ( n4942 , n1851 );
buf ( n4943 , n1169 );
buf ( n4944 , n1980 );
buf ( n4945 , n23 );
buf ( n4946 , n328 );
buf ( n4947 , n618 );
buf ( n4948 , n483 );
buf ( n4949 , n1655 );
buf ( n4950 , n1330 );
buf ( n4951 , n1031 );
buf ( n4952 , n836 );
buf ( n4953 , n431 );
buf ( n4954 , n1511 );
buf ( n4955 , n1631 );
buf ( n4956 , n471 );
buf ( n4957 , n869 );
buf ( n4958 , n428 );
buf ( n4959 , n1386 );
buf ( n4960 , n1301 );
buf ( n4961 , n650 );
buf ( n4962 , n810 );
buf ( n4963 , n1296 );
buf ( n4964 , n369 );
buf ( n4965 , n1777 );
buf ( n4966 , n1489 );
buf ( n4967 , n458 );
buf ( n4968 , n575 );
buf ( n4969 , n1343 );
buf ( n4970 , n132 );
buf ( n4971 , n1332 );
buf ( n4972 , n969 );
buf ( n4973 , n1261 );
buf ( n4974 , n1131 );
buf ( n4975 , n255 );
buf ( n4976 , n1772 );
buf ( n4977 , n1325 );
buf ( n4978 , n382 );
buf ( n4979 , n1888 );
buf ( n4980 , n1224 );
buf ( n4981 , n1702 );
buf ( n4982 , n1597 );
buf ( n4983 , n858 );
buf ( n4984 , n88 );
buf ( n4985 , n1874 );
buf ( n4986 , n743 );
buf ( n4987 , n568 );
buf ( n4988 , n1047 );
buf ( n4989 , n891 );
buf ( n4990 , n1779 );
buf ( n4991 , n301 );
buf ( n4992 , n1478 );
buf ( n4993 , n522 );
buf ( n4994 , n1013 );
buf ( n4995 , n1477 );
buf ( n4996 , n1404 );
buf ( n4997 , n610 );
buf ( n4998 , n1111 );
buf ( n4999 , n1518 );
buf ( n5000 , n1149 );
buf ( n5001 , n1808 );
buf ( n5002 , n1700 );
buf ( n5003 , n763 );
buf ( n5004 , n462 );
buf ( n5005 , n1078 );
buf ( n5006 , n709 );
buf ( n5007 , n700 );
buf ( n5008 , n852 );
buf ( n5009 , n658 );
buf ( n5010 , n961 );
buf ( n5011 , n461 );
buf ( n5012 , n850 );
buf ( n5013 , n1120 );
buf ( n5014 , n1619 );
buf ( n5015 , n721 );
buf ( n5016 , n576 );
buf ( n5017 , n800 );
buf ( n5018 , n1485 );
buf ( n5019 , n1941 );
buf ( n5020 , n695 );
buf ( n5021 , n292 );
buf ( n5022 , n923 );
buf ( n5023 , n1432 );
buf ( n5024 , n717 );
buf ( n5025 , n1767 );
buf ( n5026 , n1598 );
buf ( n5027 , n566 );
buf ( n5028 , n176 );
buf ( n5029 , n2131 );
buf ( n5030 , n383 );
buf ( n5031 , n1499 );
buf ( n5032 , n83 );
buf ( n5033 , n1590 );
buf ( n5034 , n1672 );
buf ( n5035 , n1192 );
buf ( n5036 , n1073 );
buf ( n5037 , n663 );
buf ( n5038 , n442 );
buf ( n5039 , n1508 );
buf ( n5040 , n1116 );
buf ( n5041 , n1765 );
buf ( n5042 , n293 );
buf ( n5043 , n856 );
buf ( n5044 , n645 );
buf ( n5045 , n2120 );
buf ( n5046 , n1594 );
buf ( n5047 , n640 );
buf ( n5048 , n713 );
buf ( n5049 , n113 );
buf ( n5050 , n242 );
buf ( n5051 , n96 );
buf ( n5052 , n1460 );
buf ( n5053 , n344 );
buf ( n5054 , n779 );
buf ( n5055 , n5 );
buf ( n5056 , n1778 );
buf ( n5057 , n217 );
buf ( n5058 , n165 );
buf ( n5059 , n1135 );
buf ( n5060 , n1863 );
buf ( n5061 , n530 );
buf ( n5062 , n469 );
buf ( n5063 , n1204 );
buf ( n5064 , n1144 );
buf ( n5065 , n1822 );
buf ( n5066 , n1154 );
buf ( n5067 , n863 );
buf ( n5068 , n1845 );
buf ( n5069 , n99 );
buf ( n5070 , n1197 );
buf ( n5071 , n414 );
buf ( n5072 , n108 );
buf ( n5073 , n823 );
buf ( n5074 , n706 );
buf ( n5075 , n951 );
buf ( n5076 , n368 );
buf ( n5077 , n606 );
buf ( n5078 , n93 );
buf ( n5079 , n684 );
buf ( n5080 , n2134 );
buf ( n5081 , n1839 );
buf ( n5082 , n1410 );
buf ( n5083 , n646 );
buf ( n5084 , n1387 );
buf ( n5085 , n2045 );
buf ( n5086 , n435 );
buf ( n5087 , n905 );
buf ( n5088 , n1901 );
buf ( n5089 , n296 );
buf ( n5090 , n410 );
buf ( n5091 , n896 );
buf ( n5092 , n1520 );
buf ( n5093 , n987 );
buf ( n5094 , n2064 );
buf ( n5095 , n213 );
buf ( n5096 , n1742 );
buf ( n5097 , n2054 );
buf ( n5098 , n1444 );
buf ( n5099 , n1456 );
buf ( n5100 , n1286 );
buf ( n5101 , n42 );
buf ( n5102 , n643 );
buf ( n5103 , n1793 );
buf ( n5104 , n1889 );
buf ( n5105 , n1450 );
buf ( n5106 , n1316 );
buf ( n5107 , n956 );
buf ( n5108 , n1654 );
buf ( n5109 , n1914 );
buf ( n5110 , n41 );
buf ( n5111 , n2048 );
buf ( n5112 , n1101 );
buf ( n5113 , n1764 );
buf ( n5114 , n202 );
buf ( n5115 , n996 );
buf ( n5116 , n1007 );
buf ( n5117 , n612 );
buf ( n5118 , n1740 );
buf ( n5119 , n559 );
buf ( n5120 , n323 );
buf ( n5121 , n152 );
buf ( n5122 , n875 );
buf ( n5123 , n358 );
buf ( n5124 , n1353 );
buf ( n5125 , n1524 );
buf ( n5126 , n460 );
buf ( n5127 , n1699 );
buf ( n5128 , n1252 );
buf ( n5129 , n353 );
buf ( n5130 , n948 );
buf ( n5131 , n1428 );
buf ( n5132 , n827 );
buf ( n5133 , n642 );
buf ( n5134 , n231 );
buf ( n5135 , n40 );
buf ( n5136 , n199 );
buf ( n5137 , n1308 );
buf ( n5138 , n1943 );
buf ( n5139 , n1003 );
buf ( n5140 , n644 );
buf ( n5141 , n1589 );
buf ( n5142 , n2097 );
buf ( n5143 , n319 );
buf ( n5144 , n425 );
buf ( n5145 , n2008 );
buf ( n5146 , n1449 );
buf ( n5147 , n1960 );
buf ( n5148 , n1055 );
buf ( n5149 , n409 );
buf ( n5150 , n1472 );
buf ( n5151 , n2037 );
buf ( n5152 , n718 );
buf ( n5153 , n107 );
buf ( n5154 , n2116 );
buf ( n5155 , n268 );
buf ( n5156 , n1709 );
buf ( n5157 , n228 );
buf ( n5158 , n1352 );
buf ( n5159 , n922 );
buf ( n5160 , n1850 );
buf ( n5161 , n1004 );
buf ( n5162 , n1815 );
buf ( n5163 , n844 );
buf ( n5164 , n1165 );
buf ( n5165 , n2144 );
buf ( n5166 , n1719 );
buf ( n5167 , n486 );
buf ( n5168 , n1586 );
buf ( n5169 , n1983 );
buf ( n5170 , n1257 );
buf ( n5171 , n796 );
buf ( n5172 , n967 );
buf ( n5173 , n1841 );
buf ( n5174 , n2141 );
buf ( n5175 , n391 );
buf ( n5176 , n500 );
buf ( n5177 , n1637 );
buf ( n5178 , n881 );
buf ( n5179 , n864 );
buf ( n5180 , n1977 );
buf ( n5181 , n1094 );
buf ( n5182 , n866 );
buf ( n5183 , n453 );
buf ( n5184 , n161 );
buf ( n5185 , n595 );
buf ( n5186 , n1974 );
buf ( n5187 , n248 );
buf ( n5188 , n971 );
buf ( n5189 , n1706 );
buf ( n5190 , n1963 );
buf ( n5191 , n540 );
buf ( n5192 , n758 );
buf ( n5193 , n1251 );
buf ( n5194 , n1218 );
buf ( n5195 , n1324 );
buf ( n5196 , n1265 );
buf ( n5197 , n959 );
buf ( n5198 , n1091 );
buf ( n5199 , n1784 );
buf ( n5200 , n1703 );
buf ( n5201 , n1730 );
buf ( n5202 , n1530 );
buf ( n5203 , n1 );
buf ( n5204 , n1311 );
buf ( n5205 , n450 );
buf ( n5206 , n22 );
buf ( n5207 , n1266 );
buf ( n5208 , n122 );
buf ( n5209 , n1080 );
buf ( n5210 , n1972 );
buf ( n5211 , n2033 );
buf ( n5212 , n1179 );
buf ( n5213 , n943 );
buf ( n5214 , n1000 );
buf ( n5215 , n1726 );
buf ( n5216 , n1369 );
buf ( n5217 , n2052 );
buf ( n5218 , n981 );
buf ( n5219 , n1491 );
buf ( n5220 , n2092 );
buf ( n5221 , n1201 );
buf ( n5222 , n259 );
buf ( n5223 , n160 );
buf ( n5224 , n290 );
buf ( n5225 , n603 );
buf ( n5226 , n597 );
buf ( n5227 , n2065 );
buf ( n5228 , n1537 );
buf ( n5229 , n1912 );
buf ( n5230 , n545 );
buf ( n5231 , n1175 );
buf ( n5232 , n147 );
buf ( n5233 , n72 );
buf ( n5234 , n1919 );
buf ( n5235 , n2043 );
buf ( n5236 , n1493 );
buf ( n5237 , n698 );
buf ( n5238 , n916 );
buf ( n5239 , n1212 );
buf ( n5240 , n1365 );
buf ( n5241 , n338 );
buf ( n5242 , n653 );
buf ( n5243 , n1264 );
buf ( n5244 , n1515 );
buf ( n5245 , n957 );
buf ( n5246 , n989 );
buf ( n5247 , n1425 );
buf ( n5248 , n494 );
buf ( n5249 , n550 );
buf ( n5250 , n1396 );
buf ( n5251 , n1364 );
buf ( n5252 , n457 );
buf ( n5253 , n1025 );
buf ( n5254 , n1305 );
buf ( n5255 , n286 );
buf ( n5256 , n2118 );
buf ( n5257 , n1281 );
buf ( n5258 , n1758 );
buf ( n5259 , n1546 );
buf ( n5260 , n443 );
buf ( n5261 , n797 );
buf ( n5262 , n1688 );
buf ( n5263 , n1548 );
buf ( n5264 , n119 );
buf ( n5265 , n671 );
buf ( n5266 , n1326 );
buf ( n5267 , n2034 );
buf ( n5268 , n1946 );
buf ( n5269 , n1479 );
buf ( n5270 , n277 );
buf ( n5271 , n356 );
buf ( n5272 , n1475 );
buf ( n5273 , n1104 );
buf ( n5274 , n3 );
buf ( n5275 , n1613 );
buf ( n5276 , n1053 );
buf ( n5277 , n1862 );
buf ( n5278 , n79 );
buf ( n5279 , n940 );
buf ( n5280 , n2149 );
buf ( n5281 , n139 );
buf ( n5282 , n1575 );
buf ( n5283 , n1556 );
buf ( n5284 , n219 );
buf ( n5285 , n223 );
buf ( n5286 , n227 );
buf ( n5287 , n1214 );
buf ( n5288 , n783 );
buf ( n5289 , n472 );
buf ( n5290 , n1707 );
buf ( n5291 , n1738 );
buf ( n5292 , n142 );
buf ( n5293 , n1837 );
buf ( n5294 , n1990 );
buf ( n5295 , n1198 );
buf ( n5296 , n1016 );
buf ( n5297 , n1355 );
buf ( n5298 , n1012 );
buf ( n5299 , n1126 );
buf ( n5300 , n352 );
buf ( n5301 , n1687 );
buf ( n5302 , n1020 );
buf ( n5303 , n887 );
buf ( n5304 , n979 );
buf ( n5305 , n962 );
buf ( n5306 , n0 );
buf ( n5307 , n895 );
buf ( n5308 , n10 );
buf ( n5309 , n1756 );
buf ( n5310 , n950 );
buf ( n5311 , n2108 );
buf ( n5312 , n1227 );
buf ( n5313 , n1805 );
buf ( n5314 , n991 );
buf ( n5315 , n741 );
buf ( n5316 , n570 );
buf ( n5317 , n795 );
buf ( n5318 , n941 );
buf ( n5319 , n623 );
buf ( n5320 , n385 );
buf ( n5321 , n210 );
buf ( n5322 , n1921 );
buf ( n5323 , n865 );
buf ( n5324 , n75 );
buf ( n5325 , n757 );
buf ( n5326 , n963 );
buf ( n5327 , n678 );
buf ( n5328 , n1645 );
buf ( n5329 , n813 );
buf ( n5330 , n526 );
buf ( n5331 , n2096 );
buf ( n5332 , n46 );
buf ( n5333 , n2147 );
buf ( n5334 , n1178 );
buf ( n5335 , n26 );
buf ( n5336 , n148 );
buf ( n5337 , n1968 );
buf ( n5338 , n1632 );
buf ( n5339 , n253 );
buf ( n5340 , n427 );
buf ( n5341 , n1256 );
buf ( n5342 , n497 );
buf ( n5343 , n1761 );
buf ( n5344 , n1405 );
buf ( n5345 , n1810 );
buf ( n5346 , n65 );
buf ( n5347 , n476 );
buf ( n5348 , n1836 );
buf ( n5349 , n1903 );
buf ( n5350 , n2007 );
buf ( n5351 , n411 );
buf ( n5352 , n478 );
buf ( n5353 , n1028 );
buf ( n5354 , n1939 );
buf ( n5355 , n1490 );
buf ( n5356 , n1501 );
buf ( n5357 , n1014 );
buf ( n5358 , n1342 );
buf ( n5359 , n151 );
buf ( n5360 , n1434 );
buf ( n5361 , n651 );
buf ( n5362 , n804 );
buf ( n5363 , n1739 );
buf ( n5364 , n599 );
buf ( n5365 , n1693 );
buf ( n5366 , n1686 );
buf ( n5367 , n1573 );
buf ( n5368 , n1991 );
buf ( n5369 , n734 );
buf ( n5370 , n284 );
buf ( n5371 , n1747 );
buf ( n5372 , n1052 );
buf ( n5373 , n420 );
buf ( n5374 , n80 );
buf ( n5375 , n1533 );
buf ( n5376 , n649 );
buf ( n5377 , n1636 );
buf ( n5378 , n1894 );
buf ( n5379 , n118 );
buf ( n5380 , n473 );
buf ( n5381 , n314 );
buf ( n5382 , n878 );
buf ( n5383 , n1956 );
buf ( n5384 , n1302 );
buf ( n5385 , n516 );
buf ( n5386 , n1298 );
buf ( n5387 , n788 );
buf ( n5388 , n1878 );
buf ( n5389 , n1790 );
buf ( n5390 , n1341 );
buf ( n5391 , n1671 );
buf ( n5392 , n868 );
buf ( n5393 , n2057 );
buf ( n5394 , n1232 );
buf ( n5395 , n1712 );
buf ( n5396 , n1010 );
buf ( n5397 , n1542 );
buf ( n5398 , n1383 );
buf ( n5399 , n1788 );
buf ( n5400 , n840 );
buf ( n5401 , n585 );
buf ( n5402 , n1065 );
buf ( n5403 , n1695 );
buf ( n5404 , n1433 );
buf ( n5405 , n283 );
buf ( n5406 , n1994 );
buf ( n5407 , n1856 );
buf ( n5408 , n898 );
buf ( n5409 , n1651 );
buf ( n5410 , n1139 );
buf ( n5411 , n58 );
buf ( n5412 , n637 );
buf ( n5413 , n562 );
buf ( n5414 , n600 );
buf ( n5415 , n1108 );
buf ( n5416 , n1509 );
buf ( n5417 , n622 );
buf ( n5418 , n92 );
buf ( n5419 , n681 );
buf ( n5420 , n921 );
buf ( n5421 , n2089 );
buf ( n5422 , n2094 );
buf ( n5423 , n541 );
buf ( n5424 , n418 );
buf ( n5425 , n405 );
buf ( n5426 , n939 );
buf ( n5427 , n1599 );
buf ( n5428 , n726 );
buf ( n5429 , n1666 );
buf ( n5430 , n421 );
buf ( n5431 , n1254 );
buf ( n5432 , n1248 );
buf ( n5433 , n514 );
buf ( n5434 , n416 );
buf ( n5435 , n1928 );
buf ( n5436 , n579 );
buf ( n5437 , n129 );
buf ( n5438 , n1060 );
buf ( n5439 , n1187 );
buf ( n5440 , n4 );
buf ( n5441 , n475 );
buf ( n5442 , n1715 );
buf ( n5443 , n1969 );
buf ( n5444 , n2046 );
buf ( n5445 , n2080 );
buf ( n5446 , n531 );
buf ( n5447 , n2150 );
buf ( n5448 , n1566 );
buf ( n5449 , n285 );
buf ( n5450 , n1675 );
buf ( n5451 , n366 );
buf ( n5452 , n793 );
buf ( n5453 , n1422 );
buf ( n5454 , n1121 );
buf ( n5455 , n664 );
buf ( n5456 , n792 );
buf ( n5457 , n222 );
buf ( n5458 , n771 );
buf ( n5459 , n1338 );
buf ( n5460 , n835 );
buf ( n5461 , n1074 );
buf ( n5462 , n1321 );
buf ( n5463 , n78 );
buf ( n5464 , n246 );
buf ( n5465 , n710 );
buf ( n5466 , n690 );
buf ( n5467 , n109 );
buf ( n5468 , n1933 );
buf ( n5469 , n1237 );
buf ( n5470 , n587 );
buf ( n5471 , n1905 );
buf ( n5472 , n417 );
buf ( n5473 , n1906 );
buf ( n5474 , n254 );
buf ( n5475 , n1834 );
buf ( n5476 , n1617 );
buf ( n5477 , n1103 );
buf ( n5478 , n1964 );
buf ( n5479 , n1306 );
buf ( n5480 , n408 );
buf ( n5481 , n1981 );
buf ( n5482 , n1909 );
buf ( n5483 , n1284 );
buf ( n5484 , n1569 );
buf ( n5485 , n534 );
buf ( n5486 , n1993 );
buf ( n5487 , n1760 );
buf ( n5488 , n974 );
buf ( n5489 , n305 );
buf ( n5490 , n549 );
buf ( n5491 , n1669 );
buf ( n5492 , n351 );
buf ( n5493 , n1032 );
buf ( n5494 , n1046 );
buf ( n5495 , n1622 );
buf ( n5496 , n945 );
buf ( n5497 , n376 );
buf ( n5498 , n1830 );
buf ( n5499 , n50 );
buf ( n5500 , n1940 );
buf ( n5501 , n680 );
buf ( n5502 , n1051 );
buf ( n5503 , n1868 );
buf ( n5504 , n1945 );
buf ( n5505 , n1665 );
buf ( n5506 , n778 );
buf ( n5507 , n1593 );
buf ( n5508 , n1624 );
buf ( n5509 , n714 );
buf ( n5510 , n723 );
buf ( n5511 , n1220 );
buf ( n5512 , n224 );
buf ( n5513 , n754 );
buf ( n5514 , n1279 );
buf ( n5515 , n234 );
buf ( n5516 , n1177 );
buf ( n5517 , n794 );
buf ( n5518 , n15 );
buf ( n5519 , n69 );
buf ( n5520 , n874 );
buf ( n5521 , n1234 );
buf ( n5522 , n748 );
buf ( n5523 , n1944 );
buf ( n5524 , n1659 );
buf ( n5525 , n1570 );
buf ( n5526 , n1195 );
buf ( n5527 , n273 );
buf ( n5528 , n432 );
buf ( n5529 , n343 );
buf ( n5530 , n346 );
buf ( n5531 , n2021 );
buf ( n5532 , n2138 );
buf ( n5533 , n1870 );
buf ( n5534 , n1746 );
buf ( n5535 , n455 );
buf ( n5536 , n1514 );
buf ( n5537 , n1929 );
buf ( n5538 , n2121 );
buf ( n5539 , n459 );
buf ( n5540 , n2101 );
buf ( n5541 , n1162 );
buf ( n5542 , n674 );
buf ( n5543 , n838 );
buf ( n5544 , n870 );
buf ( n5545 , n2006 );
buf ( n5546 , n192 );
buf ( n5547 , n2051 );
buf ( n5548 , n1774 );
buf ( n5549 , n1527 );
buf ( n5550 , n499 );
buf ( n5551 , n2023 );
buf ( n5552 , n1610 );
buf ( n5553 , n16 );
buf ( n5554 , n502 );
buf ( n5555 , n1189 );
buf ( n5556 , n2070 );
buf ( n5557 , n607 );
buf ( n5558 , n1690 );
buf ( n5559 , n2001 );
buf ( n5560 , n281 );
buf ( n5561 , n153 );
buf ( n5562 , n998 );
buf ( n5563 , n270 );
buf ( n5564 , n64 );
buf ( n5565 , n1821 );
buf ( n5566 , n1040 );
buf ( n5567 , n37 );
buf ( n5568 , n2038 );
buf ( n5569 , n215 );
buf ( n5570 , n1345 );
buf ( n5571 , n57 );
buf ( n5572 , n1470 );
buf ( n5573 , n715 );
buf ( n5574 , n1147 );
buf ( n5575 , n2113 );
buf ( n5576 , n2104 );
buf ( n5577 , n1081 );
buf ( n5578 , n1415 );
buf ( n5579 , n441 );
buf ( n5580 , n1299 );
buf ( n5581 , n1554 );
buf ( n5582 , n1516 );
buf ( n5583 , n1559 );
buf ( n5584 , n1936 );
buf ( n5585 , n9 );
buf ( n5586 , n814 );
buf ( n5587 , n2129 );
buf ( n5588 , n581 );
buf ( n5589 , n94 );
buf ( n5590 , n1893 );
buf ( n5591 , n1861 );
buf ( n5592 , n1168 );
buf ( n5593 , n1842 );
buf ( n5594 , n790 );
buf ( n5595 , n590 );
buf ( n5596 , n1392 );
buf ( n5597 , n233 );
buf ( n5598 , n1796 );
buf ( n5599 , n564 );
buf ( n5600 , n2030 );
buf ( n5601 , n1887 );
buf ( n5602 , n1484 );
buf ( n5603 , n1591 );
buf ( n5604 , n791 );
buf ( n5605 , n1211 );
buf ( n5606 , n1417 );
buf ( n5607 , n1729 );
buf ( n5608 , n1448 );
buf ( n5609 , n444 );
buf ( n5610 , n1931 );
buf ( n5611 , n1375 );
buf ( n5612 , n1440 );
buf ( n5613 , n168 );
buf ( n5614 , n1843 );
buf ( n5615 , n1971 );
buf ( n5616 , n1233 );
buf ( n5617 , n1106 );
buf ( n5618 , n1163 );
buf ( n5619 , n574 );
buf ( n5620 , n1190 );
buf ( n5621 , n1639 );
buf ( n5622 , n1838 );
buf ( n5623 , n1902 );
buf ( n5624 , n1421 );
buf ( n5625 , n1124 );
buf ( n5626 , n2099 );
buf ( n5627 , n815 );
buf ( n5628 , n1934 );
buf ( n5629 , n620 );
buf ( n5630 , n1635 );
buf ( n5631 , n313 );
buf ( n5632 , n704 );
buf ( n5633 , n781 );
buf ( n5634 , n1847 );
buf ( n5635 , n1161 );
buf ( n5636 , n982 );
buf ( n5637 , n968 );
buf ( n5638 , n1734 );
buf ( n5639 , n1978 );
buf ( n5640 , n2059 );
buf ( n5641 , n243 );
buf ( n5642 , n1278 );
buf ( n5643 , n624 );
buf ( n5644 , n614 );
buf ( n5645 , n1817 );
buf ( n5646 , n1270 );
buf ( n5647 , n806 );
buf ( n5648 , n1335 );
buf ( n5649 , n2061 );
buf ( n5650 , n1865 );
buf ( n5651 , n1304 );
buf ( n5652 , n608 );
buf ( n5653 , n613 );
buf ( n5654 , n1967 );
buf ( n5655 , n1503 );
buf ( n5656 , n970 );
buf ( n5657 , n589 );
buf ( n5658 , n1521 );
buf ( n5659 , n2139 );
buf ( n5660 , n2047 );
buf ( n5661 , n913 );
buf ( n5662 , n1402 );
buf ( n5663 , n985 );
buf ( n5664 , n357 );
buf ( n5665 , n1539 );
buf ( n5666 , n126 );
buf ( n5667 , n1938 );
buf ( n5668 , n1008 );
buf ( n5669 , n1022 );
buf ( n5670 , n1153 );
buf ( n5671 , n1818 );
buf ( n5672 , n56 );
buf ( n5673 , n299 );
buf ( n5674 , n155 );
buf ( n5675 , n1953 );
buf ( n5676 , n1215 );
buf ( n5677 , n1711 );
buf ( n5678 , n1183 );
buf ( n5679 , n203 );
buf ( n5680 , n1976 );
buf ( n5681 , n1487 );
buf ( n5682 , n520 );
buf ( n5683 , n47 );
buf ( n5684 , n1626 );
buf ( n5685 , n212 );
buf ( n5686 , n291 );
buf ( n5687 , n1915 );
buf ( n5688 , n1474 );
buf ( n5689 , n1567 );
buf ( n5690 , n573 );
buf ( n5691 , n849 );
buf ( n5692 , n1857 );
buf ( n5693 , n355 );
buf ( n5694 , n1900 );
buf ( n5695 , n1649 );
buf ( n5696 , n867 );
buf ( n5697 , n230 );
buf ( n5698 , n1246 );
buf ( n5699 , n1112 );
buf ( n5700 , n729 );
buf ( n5701 , n2078 );
buf ( n5702 , n452 );
buf ( n5703 , n742 );
buf ( n5704 , n1549 );
buf ( n5705 , n761 );
buf ( n5706 , n1641 );
buf ( n5707 , n1638 );
buf ( n5708 , n517 );
buf ( n5709 , n1339 );
buf ( n5710 , n1937 );
buf ( n5711 , n447 );
buf ( n5712 , n1272 );
buf ( n5713 , n750 );
buf ( n5714 , n1155 );
buf ( n5715 , n85 );
buf ( n5716 , n317 );
buf ( n5717 , n1259 );
buf ( n5718 , n1859 );
buf ( n5719 , n267 );
buf ( n5720 , n1280 );
buf ( n5721 , n532 );
buf ( n5722 , n278 );
buf ( n5723 , n1453 );
buf ( n5724 , n593 );
buf ( n5725 , n739 );
buf ( n5726 , n1543 );
buf ( n5727 , n373 );
buf ( n5728 , n1717 );
buf ( n5729 , n1340 );
buf ( n5730 , n554 );
buf ( n5731 , n993 );
buf ( n5732 , n1536 );
buf ( n5733 , n388 );
buf ( n5734 , n638 );
buf ( n5735 , n1185 );
buf ( n5736 , n485 );
buf ( n5737 , n1288 );
buf ( n5738 , n133 );
buf ( n5739 , n27 );
buf ( n5740 , n669 );
buf ( n5741 , n1041 );
buf ( n5742 , n1718 );
buf ( n5743 , n185 );
buf ( n5744 , n1193 );
buf ( n5745 , n135 );
buf ( n5746 , n1011 );
buf ( n5747 , n901 );
buf ( n5748 , n306 );
buf ( n5749 , n1267 );
buf ( n5750 , n347 );
buf ( n5751 , n1628 );
buf ( n5752 , n999 );
buf ( n5753 , n1780 );
buf ( n5754 , n1864 );
buf ( n5755 , n1083 );
buf ( n5756 , n1035 );
buf ( n5757 , n767 );
buf ( n5758 , n479 );
buf ( n5759 , n1026 );
buf ( n5760 , n803 );
buf ( n5761 , n1034 );
buf ( n5762 , n2086 );
buf ( n5763 , n995 );
buf ( n5764 , n138 );
buf ( n5765 , n1236 );
buf ( n5766 , n513 );
buf ( n5767 , n1677 );
buf ( n5768 , n110 );
buf ( n5769 , n200 );
buf ( n5770 , n257 );
buf ( n5771 , n235 );
buf ( n5772 , n1445 );
buf ( n5773 , n877 );
buf ( n5774 , n1443 );
buf ( n5775 , n229 );
buf ( n5776 , n2126 );
buf ( n5777 , n104 );
buf ( n5778 , n753 );
buf ( n5779 , n851 );
buf ( n5780 , n1984 );
buf ( n5781 , n111 );
buf ( n5782 , n911 );
buf ( n5783 , n157 );
buf ( n5784 , n899 );
buf ( n5785 , n237 );
buf ( n5786 , n1062 );
buf ( n5787 , n738 );
buf ( n5788 , n702 );
buf ( n5789 , n1627 );
buf ( n5790 , n1595 );
buf ( n5791 , n1089 );
buf ( n5792 , n740 );
buf ( n5793 , n1958 );
buf ( n5794 , n1749 );
buf ( n5795 , n1429 );
buf ( n5796 , n2137 );
buf ( n5797 , n523 );
buf ( n5798 , n266 );
buf ( n5799 , n308 );
buf ( n5800 , n252 );
buf ( n5801 , n264 );
buf ( n5802 , n2133 );
buf ( n5803 , n1125 );
buf ( n5804 , n1925 );
buf ( n5805 , n324 );
buf ( n5806 , n2140 );
buf ( n5807 , n937 );
buf ( n5808 , n1291 );
buf ( n5809 , n745 );
buf ( n5810 , n1117 );
buf ( n5811 , n1564 );
buf ( n5812 , n2004 );
buf ( n5813 , n1315 );
buf ( n5814 , n1079 );
buf ( n5815 , n1064 );
buf ( n5816 , n1273 );
buf ( n5817 , n360 );
buf ( n5818 , n1322 );
buf ( n5819 , n1327 );
buf ( n5820 , n1247 );
buf ( n5821 , n756 );
buf ( n5822 , n617 );
buf ( n5823 , n1390 );
buf ( n5824 , n807 );
buf ( n5825 , n48 );
buf ( n5826 , n920 );
buf ( n5827 , n1751 );
buf ( n5828 , n1466 );
buf ( n5829 , n504 );
buf ( n5830 , n1683 );
buf ( n5831 , n1009 );
buf ( n5832 , n1920 );
buf ( n5833 , n1471 );
buf ( n5834 , n491 );
buf ( n5835 , n392 );
buf ( n5836 , n495 );
buf ( n5837 , n1911 );
buf ( n5838 , n2000 );
buf ( n5839 , n2085 );
buf ( n5840 , n1181 );
buf ( n5841 , n1701 );
buf ( n5842 , n105 );
buf ( n5843 , n433 );
buf ( n5844 , n1182 );
buf ( n5845 , n438 );
buf ( n5846 , n661 );
buf ( n5847 , n24 );
buf ( n5848 , n1744 );
buf ( n5849 , n1704 );
buf ( n5850 , n21 );
buf ( n5851 , n972 );
buf ( n5852 , n1732 );
buf ( n5853 , n1107 );
buf ( n5854 , n402 );
buf ( n5855 , n1827 );
buf ( n5856 , n1092 );
buf ( n5857 , n240 );
buf ( n5858 , n1561 );
buf ( n5859 , n1005 );
buf ( n5860 , n716 );
buf ( n5861 , n565 );
buf ( n5862 , n289 );
buf ( n5863 , n1239 );
buf ( n5864 , n1420 );
buf ( n5865 , n1133 );
buf ( n5866 , n2105 );
buf ( n5867 , n311 );
buf ( n5868 , n805 );
buf ( n5869 , n45 );
buf ( n5870 , n1657 );
buf ( n5871 , n177 );
buf ( n5872 , n679 );
buf ( n5873 , n556 );
buf ( n5874 , n236 );
buf ( n5875 , n1319 );
buf ( n5876 , n333 );
buf ( n5877 , n61 );
buf ( n5878 , n1844 );
buf ( n5879 , n332 );
buf ( n5880 , n209 );
buf ( n5881 , n279 );
buf ( n5882 , n327 );
buf ( n5883 , n1741 );
buf ( n5884 , n555 );
buf ( n5885 , n1226 );
buf ( n5886 , n1572 );
buf ( n5887 , n250 );
buf ( n5888 , n389 );
buf ( n5889 , n873 );
buf ( n5890 , n1253 );
buf ( n5891 , n1961 );
buf ( n5892 , n1289 );
buf ( n5893 , n1552 );
buf ( n5894 , n14 );
buf ( n5895 , n1713 );
buf ( n5896 , n619 );
buf ( n5897 , n888 );
buf ( n5898 , n2084 );
buf ( n5899 , n1118 );
buf ( n5900 , n897 );
buf ( n5901 , n1876 );
buf ( n5902 , n1310 );
buf ( n5903 , n592 );
buf ( n5904 , n668 );
buf ( n5905 , n1250 );
buf ( n5906 , n1439 );
buf ( n5907 , n336 );
buf ( n5908 , n1463 );
buf ( n5909 , n1293 );
buf ( n5910 , n2056 );
buf ( n5911 , n1441 );
buf ( n5912 , n755 );
buf ( n5913 , n397 );
buf ( n5914 , n770 );
buf ( n5915 , n1049 );
buf ( n5916 , n1407 );
buf ( n5917 , n269 );
buf ( n5918 , n1890 );
buf ( n5919 , n1255 );
buf ( n5920 , n2145 );
buf ( n5921 , n1877 );
buf ( n5922 , n1899 );
buf ( n5923 , n872 );
buf ( n5924 , n274 );
buf ( n5925 , n1606 );
buf ( n5926 , n439 );
buf ( n5927 , n1037 );
buf ( n5928 , n552 );
buf ( n5929 , n481 );
buf ( n5930 , n537 );
buf ( n5931 , n381 );
buf ( n5932 , n1807 );
buf ( n5933 , n159 );
buf ( n5934 , n652 );
buf ( n5935 , n339 );
buf ( n5936 , n722 );
buf ( n5937 , n1221 );
buf ( n5938 , n1361 );
buf ( n5939 , n2062 );
buf ( n5940 , n130 );
buf ( n5941 , n1989 );
buf ( n5942 , n1924 );
buf ( n5943 , n885 );
buf ( n5944 , n125 );
buf ( n5945 , n1413 );
buf ( n5946 , n2009 );
buf ( n5947 , n605 );
buf ( n5948 , n1208 );
buf ( n5949 , n546 );
buf ( n5950 , n36 );
buf ( n5951 , n2012 );
buf ( n5952 , n720 );
buf ( n5953 , n415 );
buf ( n5954 , n752 );
buf ( n5955 , n2146 );
buf ( n5956 , n1886 );
buf ( n5957 , n359 );
buf ( n5958 , n1498 );
buf ( n5959 , n1513 );
buf ( n5960 , n1832 );
buf ( n5961 , n1954 );
buf ( n5962 , n1360 );
buf ( n5963 , n1551 );
buf ( n5964 , n2079 );
buf ( n5965 , n1720 );
buf ( n5966 , n1891 );
buf ( n5967 , n1374 );
buf ( n5968 , n1759 );
buf ( n5969 , n1127 );
buf ( n5970 , n54 );
buf ( n5971 , n551 );
buf ( n5972 , n2127 );
buf ( n5973 , n1557 );
buf ( n5974 , n1532 );
buf ( n5975 , n361 );
buf ( n5976 , n1804 );
buf ( n5977 , n1895 );
buf ( n5978 , n1303 );
buf ( n5979 , n1982 );
buf ( n5980 , n919 );
buf ( n5981 , n2032 );
buf ( n5982 , n876 );
buf ( n5983 , n197 );
buf ( n5984 , n1229 );
buf ( n5985 , n2110 );
buf ( n5986 , n1317 );
buf ( n5987 , n1130 );
buf ( n5988 , n1186 );
buf ( n5989 , n2119 );
buf ( n5990 , n1350 );
buf ( n5991 , n819 );
buf ( n5992 , n190 );
buf ( n5993 , n429 );
buf ( n5994 , n367 );
buf ( n5995 , n1398 );
buf ( n5996 , n12 );
buf ( n5997 , n1602 );
buf ( n5998 , n1753 );
buf ( n5999 , n295 );
buf ( n6000 , n1242 );
buf ( n6001 , n1465 );
buf ( n6002 , n665 );
buf ( n6003 , n1577 );
buf ( n6004 , n591 );
buf ( n6005 , n731 );
buf ( n6006 , n413 );
buf ( n6007 , n1781 );
buf ( n6008 , n966 );
buf ( n6009 , n226 );
buf ( n6010 , n86 );
buf ( n6011 , n1194 );
buf ( n6012 , n655 );
buf ( n6013 , n1263 );
buf ( n6014 , n466 );
buf ( n6015 , n464 );
buf ( n6016 , n1056 );
buf ( n6017 , n39 );
buf ( n6018 , n1072 );
buf ( n6019 , n2002 );
buf ( n6020 , n2019 );
buf ( n6021 , n501 );
buf ( n6022 , n737 );
buf ( n6023 , n318 );
buf ( n6024 , n1692 );
buf ( n6025 , n598 );
buf ( n6026 , n626 );
buf ( n6027 , n611 );
buf ( n6028 , n1745 );
buf ( n6029 , n1036 );
buf ( n6030 , n1667 );
buf ( n6031 , n925 );
buf ( n6032 , n1312 );
buf ( n6033 , n162 );
buf ( n6034 , n1584 );
buf ( n6035 , n1828 );
buf ( n6036 , n744 );
buf ( n6037 , n166 );
buf ( n6038 , n826 );
buf ( n6039 , n1540 );
buf ( n6040 , n580 );
buf ( n6041 , n1115 );
buf ( n6042 , n1986 );
buf ( n6043 , n1803 );
buf ( n6044 , n845 );
buf ( n6045 , n930 );
buf ( n6046 , n186 );
buf ( n6047 , n1860 );
buf ( n6048 , n1030 );
buf ( n6049 , n847 );
buf ( n6050 , n1414 );
buf ( n6051 , n839 );
buf ( n6052 , n325 );
buf ( n6053 , n525 );
buf ( n6054 , n569 );
buf ( n6055 , n189 );
buf ( n6056 , n1643 );
buf ( n6057 , n2106 );
buf ( n6058 , n1705 );
buf ( n6059 , n375 );
buf ( n6060 , n1069 );
buf ( n6061 , n978 );
buf ( n6062 , n893 );
buf ( n6063 , n1579 );
buf ( n6064 , n1523 );
buf ( n6065 , n440 );
buf ( n6066 , n1792 );
buf ( n6067 , n1908 );
buf ( n6068 , n198 );
buf ( n6069 , n1393 );
buf ( n6070 , n861 );
buf ( n6071 , n97 );
buf ( n6072 , n1235 );
buf ( n6073 , n1384 );
buf ( n6074 , n1469 );
buf ( n6075 , n1927 );
buf ( n6076 , n766 );
buf ( n6077 , n602 );
buf ( n6078 , n2112 );
buf ( n6079 , n1119 );
buf ( n6080 , n1174 );
buf ( n6081 , n1006 );
buf ( n6082 , n604 );
buf ( n6083 , n337 );
buf ( n6084 , n634 );
buf ( n6085 , n784 );
buf ( n6086 , n1898 );
buf ( n6087 , n1363 );
buf ( n6088 , n2132 );
buf ( n6089 , n1673 );
buf ( n6090 , n1457 );
buf ( n6091 , n1159 );
buf ( n6092 , n195 );
buf ( n6093 , n103 );
buf ( n6094 , n124 );
buf ( n6095 , n260 );
buf ( n6096 , n1806 );
buf ( n6097 , n1942 );
buf ( n6098 , n1435 );
buf ( n6099 , n1138 );
buf ( n6100 , n1160 );
buf ( n6101 , n515 );
buf ( n6102 , n1547 );
buf ( n6103 , n1173 );
buf ( n6104 , n511 );
buf ( n6105 , n654 );
buf ( n6106 , n692 );
buf ( n6107 , n1110 );
buf ( n6108 , n334 );
buf ( n6109 , n1223 );
buf ( n6110 , n463 );
buf ( n6111 , n1084 );
buf ( n6112 , n512 );
buf ( n6113 , n1833 );
buf ( n6114 , n1814 );
buf ( n6115 , n842 );
buf ( n6116 , n789 );
buf ( n6117 , n1867 );
buf ( n6118 , n1680 );
buf ( n6119 , n1835 );
buf ( n6120 , n106 );
buf ( n6121 , n1797 );
buf ( n6122 , n1058 );
buf ( n6123 , n163 );
buf ( n6124 , n128 );
buf ( n6125 , n2122 );
buf ( n6126 , n480 );
buf ( n6127 , n430 );
buf ( n6128 , n902 );
buf ( n6129 , n258 );
buf ( n6130 , n349 );
buf ( n6131 , n178 );
buf ( n6132 , n544 );
buf ( n6133 , n1388 );
buf ( n6134 , n1292 );
buf ( n6135 , n241 );
buf ( n6136 , n1813 );
buf ( n6137 , n275 );
buf ( n6138 , n263 );
buf ( n6139 , n451 );
buf ( n6140 , n910 );
buf ( n6141 , n697 );
buf ( n6142 , n374 );
buf ( n6143 , n1681 );
buf ( n6144 , n424 );
buf ( n6145 , n657 );
buf ( n6146 , n276 );
buf ( n6147 , n811 );
buf ( n6148 , n1819 );
buf ( n6149 , n89 );
buf ( n6150 , n1397 );
buf ( n6151 , n1995 );
buf ( n6152 , n329 );
buf ( n6153 , n1826 );
buf ( n6154 , n1274 );
buf ( n6155 , n802 );
buf ( n6156 , n1245 );
buf ( n6157 , n647 );
buf ( n6158 , n1999 );
buf ( n6159 , n1152 );
buf ( n6160 , n949 );
buf ( n6161 , n2014 );
buf ( n6162 , n208 );
buf ( n6163 , n2088 );
buf ( n6164 , n1061 );
buf ( n6165 , n1180 );
buf ( n6166 , n521 );
buf ( n6167 , n1601 );
buf ( n6168 , n630 );
buf ( n6169 , n1869 );
buf ( n6170 , n639 );
buf ( n6171 , n914 );
buf ( n6172 , n251 );
buf ( n6173 , n751 );
buf ( n6174 , n95 );
buf ( n6175 , n747 );
buf ( n6176 , n179 );
buf ( n6177 , n1580 );
buf ( n6178 , n1467 );
buf ( n6179 , n1768 );
buf ( n6180 , n82 );
buf ( n6181 , n1555 );
buf ( n6182 , n1723 );
buf ( n6183 , n141 );
buf ( n6184 , n953 );
buf ( n6185 , n38 );
buf ( n6186 , n1682 );
buf ( n6187 , n2098 );
buf ( n6188 , n938 );
buf ( n6189 , n239 );
buf ( n6190 , n583 );
buf ( n6191 , n1757 );
buf ( n6192 , n55 );
buf ( n6193 , n1634 );
buf ( n6194 , n66 );
buf ( n6195 , n467 );
buf ( n6196 , n1534 );
buf ( n6197 , n60 );
buf ( n6198 , n1328 );
buf ( n6199 , n1403 );
buf ( n6200 , n2035 );
buf ( n6201 , n884 );
buf ( n6202 , n918 );
buf ( n6203 , n51 );
buf ( n6204 , n928 );
buf ( n6205 , n1763 );
buf ( n6206 , n1427 );
buf ( n6207 , n1241 );
buf ( n6208 , n345 );
buf ( n6209 , n1408 );
buf ( n6210 , n315 );
buf ( n6211 , n1172 );
buf ( n6212 , n1071 );
buf ( n6213 , n1829 );
buf ( n6214 , n1783 );
buf ( n6215 , n1923 );
buf ( n6216 , n535 );
buf ( n6217 , n183 );
buf ( n6218 , n965 );
buf ( n6219 , n1213 );
buf ( n6220 , n20 );
buf ( n6221 , n1782 );
buf ( n6222 , n1646 );
buf ( n6223 , n609 );
buf ( n6224 , n975 );
buf ( n6225 , n1798 );
buf ( n6226 , n174 );
buf ( n6227 , n1038 );
buf ( n6228 , n1416 );
buf ( n6229 , n1423 );
buf ( n6230 , n204 );
buf ( n6231 , n1918 );
buf ( n6232 , n1748 );
buf ( n6233 , n596 );
buf ( n6234 , n1949 );
buf ( n6235 , n400 );
buf ( n6236 , n768 );
buf ( n6237 , n1128 );
buf ( n6238 , n310 );
buf ( n6239 , n386 );
buf ( n6240 , n1771 );
buf ( n6241 , n1522 );
buf ( n6242 , n1770 );
buf ( n6243 , n703 );
buf ( n6244 , n1320 );
buf ( n6245 , n533 );
buf ( n6246 , n2069 );
buf ( n6247 , n2081 );
buf ( n6248 , n1785 );
buf ( n6249 , n2044 );
buf ( n6250 , n1399 );
buf ( n6251 , n955 );
buf ( n6252 , n773 );
buf ( n6253 , n1446 );
buf ( n6254 , n1480 );
buf ( n6255 , n1605 );
buf ( n6256 , n434 );
buf ( n6257 , n1362 );
buf ( n6258 , n1381 );
buf ( n6259 , n1910 );
buf ( n6260 , n1769 );
buf ( n6261 , n1853 );
buf ( n6262 , n1710 );
buf ( n6263 , n947 );
buf ( n6264 , n672 );
buf ( n6265 , n1437 );
buf ( n6266 , n112 );
buf ( n6267 , n380 );
buf ( n6268 , n1451 );
buf ( n6269 , n321 );
buf ( n6270 , n1494 );
buf ( n6271 , n1996 );
buf ( n6272 , n1258 );
buf ( n6273 , n2060 );
buf ( n6274 , n1802 );
buf ( n6275 , n1517 );
buf ( n6276 , n2010 );
buf ( n6277 , n1068 );
buf ( n6278 , n393 );
buf ( n6279 , n759 );
buf ( n6280 , n1216 );
buf ( n6281 , n764 );
buf ( n6282 , n1367 );
buf ( n6283 , n519 );
buf ( n6284 , n1615 );
buf ( n6285 , n304 );
buf ( n6286 , n348 );
buf ( n6287 , n506 );
buf ( n6288 , n1644 );
buf ( n6289 , n300 );
buf ( n6290 , n320 );
buf ( n6291 , n1892 );
buf ( n6292 , n831 );
buf ( n6293 , n1329 );
buf ( n6294 , n1066 );
buf ( n6295 , n1684 );
buf ( n6296 , n482 );
buf ( n6297 , n1199 );
buf ( n6298 , n194 );
buf ( n6299 , n1588 );
buf ( n6300 , n1896 );
buf ( n6301 , n833 );
buf ( n6302 , n1346 );
buf ( n6303 , n547 );
buf ( n6304 , n536 );
buf ( n6305 , n935 );
buf ( n6306 , n1307 );
buf ( n6307 , n862 );
buf ( n6308 , n1188 );
buf ( n6309 , n892 );
buf ( n6310 , n1519 );
buf ( n6311 , n170 );
buf ( n6312 , n474 );
buf ( n6313 , n1698 );
buf ( n6314 , n696 );
buf ( n6315 , n1662 );
buf ( n6316 , n855 );
buf ( n6317 , n1395 );
buf ( n6318 , n1087 );
buf ( n6319 , n446 );
buf ( n6320 , n1750 );
buf ( n6321 , n1571 );
buf ( n6322 , n144 );
buf ( n6323 , n1373 );
buf ( n6324 , n628 );
buf ( n6325 , n1468 );
buf ( n6326 , n977 );
buf ( n6327 , n1988 );
buf ( n6328 , n1823 );
buf ( n6329 , n1260 );
buf ( n6330 , n1142 );
buf ( n6331 , n1904 );
buf ( n6332 , n1545 );
buf ( n6333 , n787 );
buf ( n6334 , n2073 );
buf ( n6335 , n1809 );
buf ( n6336 , n1563 );
buf ( n6337 , n164 );
buf ( n6338 , n1975 );
buf ( n6339 , n238 );
buf ( n6340 , n1411 );
buf ( n6341 , n390 );
buf ( n6342 , n1070 );
buf ( n6343 , n2111 );
buf ( n6344 , n627 );
buf ( n6345 , n1483 );
buf ( n6346 , n256 );
buf ( n6347 , n1418 );
buf ( n6348 , n1560 );
buf ( n6349 , n1642 );
buf ( n6350 , n1114 );
buf ( n6351 , n1917 );
buf ( n6352 , n952 );
buf ( n6353 , n1203 );
buf ( n6354 , n1184 );
buf ( n6355 , n2125 );
buf ( n6356 , n2041 );
buf ( n6357 , n1883 );
buf ( n6358 , n817 );
buf ( n6359 , n1044 );
buf ( n6360 , n711 );
buf ( n6361 , n1376 );
buf ( n6362 , n1504 );
buf ( n6363 , n1664 );
buf ( n6364 , n1442 );
buf ( n6365 , n1424 );
buf ( n6366 , n809 );
buf ( n6367 , n934 );
buf ( n6368 , n1148 );
buf ( n6369 , n342 );
buf ( n6370 , n1743 );
buf ( n6371 , n2128 );
buf ( n6372 , n1736 );
buf ( n6373 , n973 );
buf ( n6374 , n1907 );
buf ( n6375 , n2003 );
buf ( n6376 , n1018 );
buf ( n6377 , n2115 );
buf ( n6378 , n1653 );
buf ( n6379 , n1389 );
buf ( n6380 , n216 );
buf ( n6381 , n1336 );
buf ( n6382 , n7 );
buf ( n6383 , n1930 );
buf ( n6384 , n220 );
buf ( n6385 , n1276 );
buf ( n6386 , n693 );
buf ( n6387 , n1141 );
buf ( n6388 , n1210 );
buf ( n6389 , n883 );
buf ( n6390 , n1419 );
buf ( n6391 , n656 );
buf ( n6392 , n1123 );
buf ( n6393 , n561 );
buf ( n6394 , n1015 );
buf ( n6395 , n1377 );
buf ( n6396 , n309 );
buf ( n6397 , n1096 );
buf ( n6398 , n2050 );
buf ( n6399 , n1926 );
buf ( n6400 , n801 );
buf ( n6401 , n2067 );
buf ( n6402 , n1724 );
buf ( n6403 , n900 );
buf ( n6404 , n1801 );
buf ( n6405 , n1143 );
buf ( n6406 , n1331 );
buf ( n6407 , n1731 );
buf ( n6408 , n1535 );
buf ( n6409 , n1151 );
buf ( n6410 , n1604 );
buf ( n6411 , n932 );
buf ( n6412 , n196 );
buf ( n6413 , n419 );
buf ( n6414 , n1957 );
buf ( n6415 , n1002 );
buf ( n6416 , n43 );
buf ( n6417 , n244 );
buf ( n6418 , n1840 );
buf ( n6419 , n175 );
buf ( n6420 , n2017 );
buf ( n6421 , n542 );
buf ( n6422 , n927 );
buf ( n6423 , n67 );
buf ( n6424 , n685 );
buf ( n6425 , n1661 );
buf ( n6426 , n1502 );
buf ( n6427 , n1382 );
buf ( n6428 , n156 );
buf ( n6429 , n188 );
buf ( n6430 , n538 );
buf ( n6431 , n1082 );
buf ( n6432 , n1462 );
buf ( n6433 , n11 );
buf ( n6434 , n2055 );
buf ( n6435 , n2042 );
buf ( n6436 , n2130 );
buf ( n6437 , n1791 );
buf ( n6438 , n785 );
buf ( n6439 , n445 );
buf ( n6440 , n879 );
buf ( n6441 , n493 );
buf ( n6442 , n1476 );
buf ( n6443 , n489 );
buf ( n6444 , n527 );
buf ( n6445 , n843 );
buf ( n6446 , n145 );
buf ( n6447 , n1313 );
buf ( n6448 , n1541 );
buf ( n6449 , n193 );
buf ( n6450 , n31 );
buf ( n6451 , n1787 );
buf ( n6452 , n1196 );
buf ( n6453 , n44 );
buf ( n6454 , n187 );
buf ( n6455 , n154 );
buf ( n6456 , n1578 );
buf ( n6457 , n712 );
buf ( n6458 , n854 );
buf ( n6459 , n1581 );
buf ( n6460 , n1496 );
buf ( n6461 , n330 );
buf ( n6462 , n1050 );
buf ( n6463 , n1344 );
buf ( n6464 , n912 );
buf ( n6465 , n625 );
buf ( n6466 , n1935 );
buf ( n6467 , n25 );
buf ( n6468 , n454 );
buf ( n6469 , n2093 );
buf ( n6470 , n73 );
buf ( n6471 , n265 );
buf ( n6472 , n1238 );
buf ( n6473 , n1510 );
buf ( n6474 , n1708 );
buf ( n6475 , n4324 );
not ( n6476 , n6475 );
not ( n6477 , n6476 );
buf ( n6478 , n4325 );
buf ( n6479 , n6478 );
not ( n6480 , n6479 );
buf ( n6481 , n4326 );
not ( n6482 , n6481 );
not ( n6483 , n6482 );
or ( n6484 , n6480 , n6483 );
not ( n6485 , n6478 );
buf ( n6486 , n6481 );
nand ( n6487 , n6485 , n6486 );
nand ( n6488 , n6484 , n6487 );
buf ( n6489 , n4327 );
buf ( n6490 , n6489 );
and ( n6491 , n6488 , n6490 );
not ( n6492 , n6488 );
not ( n6493 , n6489 );
and ( n6494 , n6492 , n6493 );
nor ( n6495 , n6491 , n6494 );
buf ( n6496 , n4328 );
not ( n6497 , n6496 );
buf ( n6498 , n4329 );
nand ( n6499 , n6497 , n6498 );
not ( n6500 , n6499 );
buf ( n6501 , n6500 );
buf ( n6502 , n6501 );
buf ( n6503 , n4330 );
nand ( n6504 , n6502 , n6503 );
buf ( n6505 , n4331 );
buf ( n6506 , n6505 );
and ( n6507 , n6504 , n6506 );
not ( n6508 , n6504 );
not ( n6509 , n6505 );
and ( n6510 , n6508 , n6509 );
nor ( n6511 , n6507 , n6510 );
xor ( n6512 , n6495 , n6511 );
buf ( n6513 , n6500 );
buf ( n6514 , n6513 );
buf ( n6515 , n6514 );
buf ( n6516 , n4332 );
nand ( n6517 , n6515 , n6516 );
buf ( n6518 , n4333 );
buf ( n6519 , n6518 );
and ( n6520 , n6517 , n6519 );
not ( n6521 , n6517 );
not ( n6522 , n6518 );
and ( n6523 , n6521 , n6522 );
nor ( n6524 , n6520 , n6523 );
xnor ( n6525 , n6512 , n6524 );
not ( n6526 , n6525 );
not ( n6527 , n6526 );
or ( n6528 , n6477 , n6527 );
not ( n6529 , n6476 );
nand ( n6530 , n6529 , n6525 );
nand ( n6531 , n6528 , n6530 );
buf ( n6532 , n4334 );
buf ( n6533 , n6532 );
not ( n6534 , n6533 );
buf ( n6535 , n4335 );
not ( n6536 , n6535 );
not ( n6537 , n6536 );
or ( n6538 , n6534 , n6537 );
not ( n6539 , n6532 );
buf ( n6540 , n6535 );
nand ( n6541 , n6539 , n6540 );
nand ( n6542 , n6538 , n6541 );
buf ( n6543 , n4336 );
buf ( n6544 , n6543 );
and ( n6545 , n6542 , n6544 );
not ( n6546 , n6542 );
not ( n6547 , n6543 );
and ( n6548 , n6546 , n6547 );
nor ( n6549 , n6545 , n6548 );
buf ( n6550 , n4337 );
nand ( n6551 , n6502 , n6550 );
buf ( n6552 , n4338 );
xor ( n6553 , n6551 , n6552 );
xor ( n6554 , n6549 , n6553 );
buf ( n6555 , n6500 );
buf ( n6556 , n6555 );
buf ( n6557 , n6556 );
buf ( n6558 , n6557 );
buf ( n6559 , n4339 );
nand ( n6560 , n6558 , n6559 );
buf ( n6561 , n4340 );
buf ( n6562 , n6561 );
and ( n6563 , n6560 , n6562 );
not ( n6564 , n6560 );
not ( n6565 , n6561 );
and ( n6566 , n6564 , n6565 );
nor ( n6567 , n6563 , n6566 );
xnor ( n6568 , n6554 , n6567 );
not ( n6569 , n6568 );
and ( n6570 , n6531 , n6569 );
not ( n6571 , n6531 );
buf ( n6572 , n6568 );
and ( n6573 , n6571 , n6572 );
nor ( n6574 , n6570 , n6573 );
not ( n6575 , n6574 );
buf ( n6576 , n6555 );
buf ( n6577 , n6576 );
buf ( n6578 , n4341 );
nand ( n6579 , n6577 , n6578 );
buf ( n6580 , n4342 );
buf ( n6581 , n6580 );
and ( n6582 , n6579 , n6581 );
not ( n6583 , n6579 );
not ( n6584 , n6580 );
and ( n6585 , n6583 , n6584 );
nor ( n6586 , n6582 , n6585 );
buf ( n6587 , n6586 );
not ( n6588 , n6587 );
buf ( n6589 , n4343 );
buf ( n6590 , n4344 );
not ( n6591 , n6590 );
buf ( n6592 , n4345 );
buf ( n6593 , n6592 );
and ( n6594 , n6591 , n6593 );
not ( n6595 , n6591 );
not ( n6596 , n6592 );
and ( n6597 , n6595 , n6596 );
nor ( n6598 , n6594 , n6597 );
not ( n6599 , n6598 );
xor ( n6600 , n6589 , n6599 );
buf ( n6601 , n4346 );
buf ( n6602 , n4347 );
xor ( n6603 , n6601 , n6602 );
buf ( n6604 , n6556 );
buf ( n6605 , n6604 );
buf ( n6606 , n4348 );
nand ( n6607 , n6605 , n6606 );
xnor ( n6608 , n6603 , n6607 );
xnor ( n6609 , n6600 , n6608 );
not ( n6610 , n6609 );
not ( n6611 , n6610 );
or ( n6612 , n6588 , n6611 );
or ( n6613 , n6610 , n6587 );
nand ( n6614 , n6612 , n6613 );
buf ( n6615 , n4349 );
buf ( n6616 , n6615 );
not ( n6617 , n6616 );
buf ( n6618 , n4350 );
not ( n6619 , n6618 );
not ( n6620 , n6619 );
or ( n6621 , n6617 , n6620 );
not ( n6622 , n6615 );
buf ( n6623 , n6618 );
nand ( n6624 , n6622 , n6623 );
nand ( n6625 , n6621 , n6624 );
buf ( n6626 , n4351 );
not ( n6627 , n6626 );
and ( n6628 , n6625 , n6627 );
not ( n6629 , n6625 );
buf ( n6630 , n6626 );
and ( n6631 , n6629 , n6630 );
nor ( n6632 , n6628 , n6631 );
buf ( n6633 , n6513 );
buf ( n6634 , n6633 );
buf ( n6635 , n4352 );
nand ( n6636 , n6634 , n6635 );
buf ( n6637 , n4353 );
buf ( n6638 , n6637 );
and ( n6639 , n6636 , n6638 );
not ( n6640 , n6636 );
not ( n6641 , n6637 );
and ( n6642 , n6640 , n6641 );
nor ( n6643 , n6639 , n6642 );
xor ( n6644 , n6632 , n6643 );
buf ( n6645 , n6500 );
buf ( n6646 , n6645 );
buf ( n6647 , n6646 );
buf ( n6648 , n4354 );
nand ( n6649 , n6647 , n6648 );
buf ( n6650 , n4355 );
buf ( n6651 , n6650 );
and ( n6652 , n6649 , n6651 );
not ( n6653 , n6649 );
not ( n6654 , n6650 );
and ( n6655 , n6653 , n6654 );
nor ( n6656 , n6652 , n6655 );
not ( n6657 , n6656 );
xnor ( n6658 , n6644 , n6657 );
buf ( n6659 , n6658 );
and ( n6660 , n6614 , n6659 );
not ( n6661 , n6614 );
not ( n6662 , n6659 );
and ( n6663 , n6661 , n6662 );
nor ( n6664 , n6660 , n6663 );
not ( n6665 , n6664 );
nand ( n6666 , n6575 , n6665 );
not ( n6667 , n6666 );
buf ( n6668 , n4356 );
buf ( n6669 , n4357 );
not ( n6670 , n6669 );
buf ( n6671 , n4358 );
buf ( n6672 , n6671 );
nand ( n6673 , n6670 , n6672 );
not ( n6674 , n6671 );
buf ( n6675 , n6669 );
nand ( n6676 , n6674 , n6675 );
and ( n6677 , n6673 , n6676 );
xor ( n6678 , n6668 , n6677 );
buf ( n6679 , n4359 );
buf ( n6680 , n4360 );
xor ( n6681 , n6679 , n6680 );
buf ( n6682 , n4361 );
nand ( n6683 , n6605 , n6682 );
xnor ( n6684 , n6681 , n6683 );
xnor ( n6685 , n6678 , n6684 );
not ( n6686 , n6685 );
buf ( n6687 , n4362 );
buf ( n6688 , n6687 );
not ( n6689 , n6688 );
buf ( n6690 , n4363 );
buf ( n6691 , n6690 );
not ( n6692 , n6691 );
buf ( n6693 , n4364 );
not ( n6694 , n6693 );
not ( n6695 , n6694 );
or ( n6696 , n6692 , n6695 );
not ( n6697 , n6690 );
buf ( n6698 , n6693 );
nand ( n6699 , n6697 , n6698 );
nand ( n6700 , n6696 , n6699 );
buf ( n6701 , n4365 );
not ( n6702 , n6701 );
and ( n6703 , n6700 , n6702 );
not ( n6704 , n6700 );
buf ( n6705 , n6701 );
and ( n6706 , n6704 , n6705 );
nor ( n6707 , n6703 , n6706 );
buf ( n6708 , n4366 );
nand ( n6709 , n6502 , n6708 );
buf ( n6710 , n4367 );
buf ( n6711 , n6710 );
and ( n6712 , n6709 , n6711 );
not ( n6713 , n6709 );
not ( n6714 , n6710 );
and ( n6715 , n6713 , n6714 );
nor ( n6716 , n6712 , n6715 );
xor ( n6717 , n6707 , n6716 );
buf ( n6718 , n6513 );
buf ( n6719 , n6718 );
buf ( n6720 , n4368 );
nand ( n6721 , n6719 , n6720 );
buf ( n6722 , n4369 );
buf ( n6723 , n6722 );
and ( n6724 , n6721 , n6723 );
not ( n6725 , n6721 );
not ( n6726 , n6722 );
and ( n6727 , n6725 , n6726 );
nor ( n6728 , n6724 , n6727 );
xor ( n6729 , n6717 , n6728 );
not ( n6730 , n6729 );
not ( n6731 , n6730 );
not ( n6732 , n6731 );
or ( n6733 , n6689 , n6732 );
not ( n6734 , n6729 );
not ( n6735 , n6687 );
nand ( n6736 , n6734 , n6735 );
nand ( n6737 , n6733 , n6736 );
not ( n6738 , n6737 );
not ( n6739 , n6738 );
or ( n6740 , n6686 , n6739 );
not ( n6741 , n6685 );
nand ( n6742 , n6741 , n6737 );
nand ( n6743 , n6740 , n6742 );
not ( n6744 , n6743 );
and ( n6745 , n6667 , n6744 );
not ( n6746 , n6574 );
nand ( n6747 , n6746 , n6665 );
and ( n6748 , n6747 , n6743 );
nor ( n6749 , n6745 , n6748 );
not ( n6750 , n6749 );
not ( n6751 , n6750 );
buf ( n6752 , n4370 );
buf ( n6753 , n6752 );
not ( n6754 , n6753 );
buf ( n6755 , n4371 );
not ( n6756 , n6755 );
not ( n6757 , n6756 );
or ( n6758 , n6754 , n6757 );
not ( n6759 , n6752 );
buf ( n6760 , n6755 );
nand ( n6761 , n6759 , n6760 );
nand ( n6762 , n6758 , n6761 );
buf ( n6763 , n4372 );
not ( n6764 , n6763 );
and ( n6765 , n6762 , n6764 );
not ( n6766 , n6762 );
buf ( n6767 , n6763 );
and ( n6768 , n6766 , n6767 );
nor ( n6769 , n6765 , n6768 );
buf ( n6770 , n6501 );
buf ( n6771 , n4373 );
nand ( n6772 , n6770 , n6771 );
buf ( n6773 , n4374 );
buf ( n6774 , n6773 );
and ( n6775 , n6772 , n6774 );
not ( n6776 , n6772 );
not ( n6777 , n6773 );
and ( n6778 , n6776 , n6777 );
nor ( n6779 , n6775 , n6778 );
xor ( n6780 , n6769 , n6779 );
buf ( n6781 , n4375 );
nand ( n6782 , n6557 , n6781 );
buf ( n6783 , n4376 );
buf ( n6784 , n6783 );
and ( n6785 , n6782 , n6784 );
not ( n6786 , n6782 );
not ( n6787 , n6783 );
and ( n6788 , n6786 , n6787 );
nor ( n6789 , n6785 , n6788 );
not ( n6790 , n6789 );
xnor ( n6791 , n6780 , n6790 );
buf ( n6792 , n6791 );
not ( n6793 , n6792 );
buf ( n6794 , n4377 );
buf ( n6795 , n6794 );
not ( n6796 , n6795 );
buf ( n6797 , n4378 );
buf ( n6798 , n6797 );
not ( n6799 , n6798 );
buf ( n6800 , n4379 );
not ( n6801 , n6800 );
not ( n6802 , n6801 );
or ( n6803 , n6799 , n6802 );
not ( n6804 , n6797 );
buf ( n6805 , n6800 );
nand ( n6806 , n6804 , n6805 );
nand ( n6807 , n6803 , n6806 );
buf ( n6808 , n4380 );
not ( n6809 , n6808 );
and ( n6810 , n6807 , n6809 );
not ( n6811 , n6807 );
buf ( n6812 , n6808 );
and ( n6813 , n6811 , n6812 );
nor ( n6814 , n6810 , n6813 );
buf ( n6815 , n6645 );
buf ( n6816 , n6815 );
buf ( n6817 , n4381 );
nand ( n6818 , n6816 , n6817 );
buf ( n6819 , n4382 );
buf ( n6820 , n6819 );
and ( n6821 , n6818 , n6820 );
not ( n6822 , n6818 );
not ( n6823 , n6819 );
and ( n6824 , n6822 , n6823 );
nor ( n6825 , n6821 , n6824 );
xor ( n6826 , n6814 , n6825 );
buf ( n6827 , n6555 );
buf ( n6828 , n6827 );
buf ( n6829 , n4383 );
nand ( n6830 , n6828 , n6829 );
buf ( n6831 , n4384 );
buf ( n6832 , n6831 );
and ( n6833 , n6830 , n6832 );
not ( n6834 , n6830 );
not ( n6835 , n6831 );
and ( n6836 , n6834 , n6835 );
nor ( n6837 , n6833 , n6836 );
not ( n6838 , n6837 );
xnor ( n6839 , n6826 , n6838 );
not ( n6840 , n6839 );
or ( n6841 , n6796 , n6840 );
xor ( n6842 , n6814 , n6837 );
buf ( n6843 , n6825 );
xnor ( n6844 , n6842 , n6843 );
not ( n6845 , n6794 );
nand ( n6846 , n6844 , n6845 );
nand ( n6847 , n6841 , n6846 );
not ( n6848 , n6847 );
or ( n6849 , n6793 , n6848 );
or ( n6850 , n6847 , n6791 );
nand ( n6851 , n6849 , n6850 );
not ( n6852 , n6851 );
buf ( n6853 , n4385 );
buf ( n6854 , n6853 );
not ( n6855 , n6854 );
buf ( n6856 , n4386 );
not ( n6857 , n6856 );
not ( n6858 , n6857 );
or ( n6859 , n6855 , n6858 );
not ( n6860 , n6853 );
buf ( n6861 , n6856 );
nand ( n6862 , n6860 , n6861 );
nand ( n6863 , n6859 , n6862 );
buf ( n6864 , n4387 );
not ( n6865 , n6864 );
and ( n6866 , n6863 , n6865 );
not ( n6867 , n6863 );
buf ( n6868 , n6864 );
and ( n6869 , n6867 , n6868 );
nor ( n6870 , n6866 , n6869 );
buf ( n6871 , n6827 );
buf ( n6872 , n4388 );
nand ( n6873 , n6871 , n6872 );
buf ( n6874 , n4389 );
buf ( n6875 , n6874 );
and ( n6876 , n6873 , n6875 );
not ( n6877 , n6873 );
not ( n6878 , n6874 );
and ( n6879 , n6877 , n6878 );
nor ( n6880 , n6876 , n6879 );
xor ( n6881 , n6870 , n6880 );
buf ( n6882 , n4390 );
nand ( n6883 , n6647 , n6882 );
buf ( n6884 , n4391 );
not ( n6885 , n6884 );
and ( n6886 , n6883 , n6885 );
not ( n6887 , n6883 );
buf ( n6888 , n6884 );
and ( n6889 , n6887 , n6888 );
nor ( n6890 , n6886 , n6889 );
xnor ( n6891 , n6881 , n6890 );
not ( n6892 , n6891 );
not ( n6893 , n6892 );
not ( n6894 , n6893 );
buf ( n6895 , n4392 );
buf ( n6896 , n6895 );
not ( n6897 , n6896 );
buf ( n6898 , n4393 );
buf ( n6899 , n6898 );
not ( n6900 , n6899 );
buf ( n6901 , n4394 );
not ( n6902 , n6901 );
not ( n6903 , n6902 );
or ( n6904 , n6900 , n6903 );
not ( n6905 , n6898 );
buf ( n6906 , n6901 );
nand ( n6907 , n6905 , n6906 );
nand ( n6908 , n6904 , n6907 );
buf ( n6909 , n4395 );
buf ( n6910 , n6909 );
and ( n6911 , n6908 , n6910 );
not ( n6912 , n6908 );
not ( n6913 , n6909 );
and ( n6914 , n6912 , n6913 );
nor ( n6915 , n6911 , n6914 );
buf ( n6916 , n6827 );
buf ( n6917 , n4396 );
nand ( n6918 , n6916 , n6917 );
buf ( n6919 , n4397 );
buf ( n6920 , n6919 );
and ( n6921 , n6918 , n6920 );
not ( n6922 , n6918 );
not ( n6923 , n6919 );
and ( n6924 , n6922 , n6923 );
nor ( n6925 , n6921 , n6924 );
xor ( n6926 , n6915 , n6925 );
buf ( n6927 , n6645 );
buf ( n6928 , n4398 );
nand ( n6929 , n6927 , n6928 );
buf ( n6930 , n4399 );
buf ( n6931 , n6930 );
and ( n6932 , n6929 , n6931 );
not ( n6933 , n6929 );
not ( n6934 , n6930 );
and ( n6935 , n6933 , n6934 );
nor ( n6936 , n6932 , n6935 );
xnor ( n6937 , n6926 , n6936 );
not ( n6938 , n6937 );
or ( n6939 , n6897 , n6938 );
xor ( n6940 , n6915 , n6936 );
not ( n6941 , n6925 );
xnor ( n6942 , n6940 , n6941 );
not ( n6943 , n6895 );
nand ( n6944 , n6942 , n6943 );
nand ( n6945 , n6939 , n6944 );
not ( n6946 , n6945 );
or ( n6947 , n6894 , n6946 );
buf ( n6948 , n6891 );
buf ( n6949 , n6948 );
or ( n6950 , n6945 , n6949 );
nand ( n6951 , n6947 , n6950 );
nand ( n6952 , n6852 , n6951 );
buf ( n6953 , n4400 );
not ( n6954 , n6953 );
not ( n6955 , n6954 );
buf ( n6956 , n4401 );
buf ( n6957 , n4402 );
buf ( n6958 , n6957 );
not ( n6959 , n6958 );
buf ( n6960 , n4403 );
not ( n6961 , n6960 );
not ( n6962 , n6961 );
or ( n6963 , n6959 , n6962 );
not ( n6964 , n6957 );
buf ( n6965 , n6960 );
nand ( n6966 , n6964 , n6965 );
nand ( n6967 , n6963 , n6966 );
not ( n6968 , n6967 );
xor ( n6969 , n6956 , n6968 );
buf ( n6970 , n4404 );
buf ( n6971 , n4405 );
xor ( n6972 , n6970 , n6971 );
buf ( n6973 , n6916 );
buf ( n6974 , n4406 );
nand ( n6975 , n6973 , n6974 );
xnor ( n6976 , n6972 , n6975 );
xnor ( n6977 , n6969 , n6976 );
not ( n6978 , n6977 );
or ( n6979 , n6955 , n6978 );
not ( n6980 , n6954 );
xor ( n6981 , n6956 , n6967 );
xnor ( n6982 , n6981 , n6976 );
nand ( n6983 , n6980 , n6982 );
nand ( n6984 , n6979 , n6983 );
buf ( n6985 , n4407 );
buf ( n6986 , n6985 );
not ( n6987 , n6986 );
buf ( n6988 , n4408 );
not ( n6989 , n6988 );
not ( n6990 , n6989 );
or ( n6991 , n6987 , n6990 );
not ( n6992 , n6985 );
buf ( n6993 , n6988 );
nand ( n6994 , n6992 , n6993 );
nand ( n6995 , n6991 , n6994 );
buf ( n6996 , n4409 );
buf ( n6997 , n6996 );
and ( n6998 , n6995 , n6997 );
not ( n6999 , n6995 );
not ( n7000 , n6996 );
and ( n7001 , n6999 , n7000 );
nor ( n7002 , n6998 , n7001 );
buf ( n7003 , n4410 );
nand ( n7004 , n6514 , n7003 );
buf ( n7005 , n4411 );
buf ( n7006 , n7005 );
and ( n7007 , n7004 , n7006 );
not ( n7008 , n7004 );
not ( n7009 , n7005 );
and ( n7010 , n7008 , n7009 );
nor ( n7011 , n7007 , n7010 );
xor ( n7012 , n7002 , n7011 );
buf ( n7013 , n6513 );
buf ( n7014 , n7013 );
buf ( n7015 , n4412 );
nand ( n7016 , n7014 , n7015 );
buf ( n7017 , n4413 );
not ( n7018 , n7017 );
and ( n7019 , n7016 , n7018 );
not ( n7020 , n7016 );
buf ( n7021 , n7017 );
and ( n7022 , n7020 , n7021 );
nor ( n7023 , n7019 , n7022 );
xnor ( n7024 , n7012 , n7023 );
buf ( n7025 , n7024 );
not ( n7026 , n7025 );
and ( n7027 , n6984 , n7026 );
not ( n7028 , n6984 );
not ( n7029 , n7024 );
not ( n7030 , n7029 );
and ( n7031 , n7028 , n7030 );
nor ( n7032 , n7027 , n7031 );
and ( n7033 , n6952 , n7032 );
not ( n7034 , n6952 );
not ( n7035 , n7032 );
and ( n7036 , n7034 , n7035 );
nor ( n7037 , n7033 , n7036 );
not ( n7038 , n7037 );
not ( n7039 , n7038 );
not ( n7040 , n6743 );
nand ( n7041 , n7040 , n6574 );
not ( n7042 , n7041 );
buf ( n7043 , n4414 );
buf ( n7044 , n7043 );
not ( n7045 , n7044 );
buf ( n7046 , n4415 );
not ( n7047 , n7046 );
not ( n7048 , n7047 );
or ( n7049 , n7045 , n7048 );
not ( n7050 , n7043 );
buf ( n7051 , n7046 );
nand ( n7052 , n7050 , n7051 );
nand ( n7053 , n7049 , n7052 );
not ( n7054 , n7053 );
buf ( n7055 , n4416 );
not ( n7056 , n7055 );
buf ( n7057 , n4417 );
nand ( n7058 , n6577 , n7057 );
buf ( n7059 , n4418 );
buf ( n7060 , n7059 );
and ( n7061 , n7058 , n7060 );
not ( n7062 , n7058 );
not ( n7063 , n7059 );
and ( n7064 , n7062 , n7063 );
nor ( n7065 , n7061 , n7064 );
xor ( n7066 , n7056 , n7065 );
buf ( n7067 , n6770 );
buf ( n7068 , n4419 );
nand ( n7069 , n7067 , n7068 );
buf ( n7070 , n4420 );
not ( n7071 , n7070 );
and ( n7072 , n7069 , n7071 );
not ( n7073 , n7069 );
buf ( n7074 , n7070 );
and ( n7075 , n7073 , n7074 );
nor ( n7076 , n7072 , n7075 );
xnor ( n7077 , n7066 , n7076 );
not ( n7078 , n7077 );
or ( n7079 , n7054 , n7078 );
not ( n7080 , n7077 );
not ( n7081 , n7053 );
nand ( n7082 , n7080 , n7081 );
nand ( n7083 , n7079 , n7082 );
not ( n7084 , n7083 );
not ( n7085 , n7084 );
buf ( n7086 , n4421 );
buf ( n7087 , n7086 );
not ( n7088 , n7087 );
buf ( n7089 , n4422 );
buf ( n7090 , n7089 );
not ( n7091 , n7090 );
buf ( n7092 , n4423 );
not ( n7093 , n7092 );
not ( n7094 , n7093 );
or ( n7095 , n7091 , n7094 );
not ( n7096 , n7089 );
buf ( n7097 , n7092 );
nand ( n7098 , n7096 , n7097 );
nand ( n7099 , n7095 , n7098 );
buf ( n7100 , n4424 );
not ( n7101 , n7100 );
and ( n7102 , n7099 , n7101 );
not ( n7103 , n7099 );
buf ( n7104 , n7100 );
and ( n7105 , n7103 , n7104 );
nor ( n7106 , n7102 , n7105 );
buf ( n7107 , n6718 );
buf ( n7108 , n4425 );
nand ( n7109 , n7107 , n7108 );
buf ( n7110 , n4426 );
buf ( n7111 , n7110 );
and ( n7112 , n7109 , n7111 );
not ( n7113 , n7109 );
not ( n7114 , n7110 );
and ( n7115 , n7113 , n7114 );
nor ( n7116 , n7112 , n7115 );
xor ( n7117 , n7106 , n7116 );
buf ( n7118 , n4427 );
nand ( n7119 , n7067 , n7118 );
buf ( n7120 , n4428 );
buf ( n7121 , n7120 );
and ( n7122 , n7119 , n7121 );
not ( n7123 , n7119 );
not ( n7124 , n7120 );
and ( n7125 , n7123 , n7124 );
nor ( n7126 , n7122 , n7125 );
xnor ( n7127 , n7117 , n7126 );
buf ( n7128 , n7127 );
not ( n7129 , n7128 );
not ( n7130 , n7129 );
or ( n7131 , n7088 , n7130 );
or ( n7132 , n7129 , n7087 );
nand ( n7133 , n7131 , n7132 );
not ( n7134 , n7133 );
and ( n7135 , n7085 , n7134 );
not ( n7136 , n7083 );
and ( n7137 , n7136 , n7133 );
nor ( n7138 , n7135 , n7137 );
not ( n7139 , n7138 );
not ( n7140 , n7139 );
and ( n7141 , n7042 , n7140 );
and ( n7142 , n7041 , n7139 );
nor ( n7143 , n7141 , n7142 );
not ( n7144 , n7143 );
not ( n7145 , n7144 );
or ( n7146 , n7039 , n7145 );
nand ( n7147 , n7143 , n7037 );
nand ( n7148 , n7146 , n7147 );
buf ( n7149 , n4429 );
buf ( n7150 , n7149 );
buf ( n7151 , n4430 );
buf ( n7152 , n7151 );
not ( n7153 , n7152 );
buf ( n7154 , n4431 );
not ( n7155 , n7154 );
not ( n7156 , n7155 );
or ( n7157 , n7153 , n7156 );
not ( n7158 , n7151 );
buf ( n7159 , n7154 );
nand ( n7160 , n7158 , n7159 );
nand ( n7161 , n7157 , n7160 );
buf ( n7162 , n4432 );
buf ( n7163 , n7162 );
and ( n7164 , n7161 , n7163 );
not ( n7165 , n7161 );
not ( n7166 , n7162 );
and ( n7167 , n7165 , n7166 );
nor ( n7168 , n7164 , n7167 );
buf ( n7169 , n4433 );
nand ( n7170 , n6604 , n7169 );
buf ( n7171 , n4434 );
buf ( n7172 , n7171 );
and ( n7173 , n7170 , n7172 );
not ( n7174 , n7170 );
not ( n7175 , n7171 );
and ( n7176 , n7174 , n7175 );
nor ( n7177 , n7173 , n7176 );
xor ( n7178 , n7168 , n7177 );
buf ( n7179 , n4435 );
nand ( n7180 , n6816 , n7179 );
buf ( n7181 , n4436 );
not ( n7182 , n7181 );
and ( n7183 , n7180 , n7182 );
not ( n7184 , n7180 );
buf ( n7185 , n7181 );
and ( n7186 , n7184 , n7185 );
nor ( n7187 , n7183 , n7186 );
xnor ( n7188 , n7178 , n7187 );
buf ( n7189 , n7188 );
xor ( n7190 , n7150 , n7189 );
buf ( n7191 , n4437 );
buf ( n7192 , n4438 );
not ( n7193 , n7192 );
xor ( n7194 , n7191 , n7193 );
buf ( n7195 , n4439 );
not ( n7196 , n7195 );
buf ( n7197 , n6827 );
buf ( n7198 , n4440 );
nand ( n7199 , n7197 , n7198 );
not ( n7200 , n7199 );
or ( n7201 , n7196 , n7200 );
buf ( n7202 , n6576 );
nand ( n7203 , n7202 , n7198 );
or ( n7204 , n7203 , n7195 );
nand ( n7205 , n7201 , n7204 );
xnor ( n7206 , n7194 , n7205 );
not ( n7207 , n7206 );
not ( n7208 , n7207 );
buf ( n7209 , n4441 );
buf ( n7210 , n7209 );
not ( n7211 , n7210 );
buf ( n7212 , n4442 );
not ( n7213 , n7212 );
not ( n7214 , n7213 );
or ( n7215 , n7211 , n7214 );
not ( n7216 , n7209 );
buf ( n7217 , n7212 );
nand ( n7218 , n7216 , n7217 );
nand ( n7219 , n7215 , n7218 );
not ( n7220 , n7219 );
and ( n7221 , n7208 , n7220 );
and ( n7222 , n7207 , n7219 );
nor ( n7223 , n7221 , n7222 );
buf ( n7224 , n7223 );
xnor ( n7225 , n7190 , n7224 );
not ( n7226 , n7225 );
buf ( n7227 , n4443 );
not ( n7228 , n7227 );
buf ( n7229 , n4444 );
buf ( n7230 , n7229 );
not ( n7231 , n7230 );
buf ( n7232 , n4445 );
not ( n7233 , n7232 );
not ( n7234 , n7233 );
or ( n7235 , n7231 , n7234 );
not ( n7236 , n7229 );
buf ( n7237 , n7232 );
nand ( n7238 , n7236 , n7237 );
nand ( n7239 , n7235 , n7238 );
buf ( n7240 , n4446 );
not ( n7241 , n7240 );
and ( n7242 , n7239 , n7241 );
not ( n7243 , n7239 );
buf ( n7244 , n7240 );
and ( n7245 , n7243 , n7244 );
nor ( n7246 , n7242 , n7245 );
buf ( n7247 , n6514 );
buf ( n7248 , n4447 );
nand ( n7249 , n7247 , n7248 );
buf ( n7250 , n4448 );
buf ( n7251 , n7250 );
and ( n7252 , n7249 , n7251 );
not ( n7253 , n7249 );
not ( n7254 , n7250 );
and ( n7255 , n7253 , n7254 );
nor ( n7256 , n7252 , n7255 );
xor ( n7257 , n7246 , n7256 );
buf ( n7258 , n6514 );
buf ( n7259 , n7258 );
buf ( n7260 , n4449 );
nand ( n7261 , n7259 , n7260 );
buf ( n7262 , n4450 );
not ( n7263 , n7262 );
and ( n7264 , n7261 , n7263 );
not ( n7265 , n7261 );
buf ( n7266 , n7262 );
and ( n7267 , n7265 , n7266 );
nor ( n7268 , n7264 , n7267 );
xnor ( n7269 , n7257 , n7268 );
buf ( n7270 , n7269 );
not ( n7271 , n7270 );
or ( n7272 , n7228 , n7271 );
or ( n7273 , n7270 , n7227 );
nand ( n7274 , n7272 , n7273 );
buf ( n7275 , n4451 );
buf ( n7276 , n7275 );
not ( n7277 , n7276 );
buf ( n7278 , n4452 );
not ( n7279 , n7278 );
not ( n7280 , n7279 );
or ( n7281 , n7277 , n7280 );
not ( n7282 , n7275 );
buf ( n7283 , n7278 );
nand ( n7284 , n7282 , n7283 );
nand ( n7285 , n7281 , n7284 );
buf ( n7286 , n4453 );
not ( n7287 , n7286 );
and ( n7288 , n7285 , n7287 );
not ( n7289 , n7285 );
buf ( n7290 , n7286 );
and ( n7291 , n7289 , n7290 );
nor ( n7292 , n7288 , n7291 );
buf ( n7293 , n6576 );
buf ( n7294 , n4454 );
nand ( n7295 , n7293 , n7294 );
buf ( n7296 , n4455 );
buf ( n7297 , n7296 );
and ( n7298 , n7295 , n7297 );
not ( n7299 , n7295 );
not ( n7300 , n7296 );
and ( n7301 , n7299 , n7300 );
nor ( n7302 , n7298 , n7301 );
xor ( n7303 , n7292 , n7302 );
buf ( n7304 , n4456 );
nand ( n7305 , n7247 , n7304 );
buf ( n7306 , n4457 );
not ( n7307 , n7306 );
and ( n7308 , n7305 , n7307 );
not ( n7309 , n7305 );
buf ( n7310 , n7306 );
and ( n7311 , n7309 , n7310 );
nor ( n7312 , n7308 , n7311 );
xnor ( n7313 , n7303 , n7312 );
buf ( n7314 , n7313 );
buf ( n7315 , n7314 );
and ( n7316 , n7274 , n7315 );
not ( n7317 , n7274 );
not ( n7318 , n7314 );
and ( n7319 , n7317 , n7318 );
nor ( n7320 , n7316 , n7319 );
not ( n7321 , n7320 );
nand ( n7322 , n7226 , n7321 );
buf ( n7323 , n4458 );
buf ( n7324 , n7323 );
not ( n7325 , n7324 );
buf ( n7326 , n4459 );
buf ( n7327 , n7326 );
not ( n7328 , n7327 );
buf ( n7329 , n4460 );
not ( n7330 , n7329 );
not ( n7331 , n7330 );
or ( n7332 , n7328 , n7331 );
not ( n7333 , n7326 );
buf ( n7334 , n7329 );
nand ( n7335 , n7333 , n7334 );
nand ( n7336 , n7332 , n7335 );
buf ( n7337 , n4461 );
buf ( n7338 , n7337 );
and ( n7339 , n7336 , n7338 );
not ( n7340 , n7336 );
not ( n7341 , n7337 );
and ( n7342 , n7340 , n7341 );
nor ( n7343 , n7339 , n7342 );
buf ( n7344 , n6576 );
buf ( n7345 , n4462 );
nand ( n7346 , n7344 , n7345 );
buf ( n7347 , n4463 );
buf ( n7348 , n7347 );
and ( n7349 , n7346 , n7348 );
not ( n7350 , n7346 );
not ( n7351 , n7347 );
and ( n7352 , n7350 , n7351 );
nor ( n7353 , n7349 , n7352 );
xor ( n7354 , n7343 , n7353 );
buf ( n7355 , n6718 );
buf ( n7356 , n4464 );
nand ( n7357 , n7355 , n7356 );
buf ( n7358 , n4465 );
buf ( n7359 , n7358 );
and ( n7360 , n7357 , n7359 );
not ( n7361 , n7357 );
not ( n7362 , n7358 );
and ( n7363 , n7361 , n7362 );
nor ( n7364 , n7360 , n7363 );
not ( n7365 , n7364 );
xnor ( n7366 , n7354 , n7365 );
not ( n7367 , n7366 );
not ( n7368 , n7367 );
or ( n7369 , n7325 , n7368 );
not ( n7370 , n7366 );
or ( n7371 , n7370 , n7324 );
nand ( n7372 , n7369 , n7371 );
buf ( n7373 , n4466 );
buf ( n7374 , n7373 );
not ( n7375 , n7374 );
buf ( n7376 , n4467 );
not ( n7377 , n7376 );
not ( n7378 , n7377 );
or ( n7379 , n7375 , n7378 );
not ( n7380 , n7373 );
buf ( n7381 , n7376 );
nand ( n7382 , n7380 , n7381 );
nand ( n7383 , n7379 , n7382 );
buf ( n7384 , n4468 );
not ( n7385 , n7384 );
and ( n7386 , n7383 , n7385 );
not ( n7387 , n7383 );
buf ( n7388 , n7384 );
and ( n7389 , n7387 , n7388 );
nor ( n7390 , n7386 , n7389 );
buf ( n7391 , n4469 );
nand ( n7392 , n6815 , n7391 );
buf ( n7393 , n4470 );
not ( n7394 , n7393 );
and ( n7395 , n7392 , n7394 );
not ( n7396 , n7392 );
buf ( n7397 , n7393 );
and ( n7398 , n7396 , n7397 );
nor ( n7399 , n7395 , n7398 );
xor ( n7400 , n7390 , n7399 );
buf ( n7401 , n4471 );
nand ( n7402 , n6634 , n7401 );
buf ( n7403 , n4472 );
not ( n7404 , n7403 );
and ( n7405 , n7402 , n7404 );
not ( n7406 , n7402 );
buf ( n7407 , n7403 );
and ( n7408 , n7406 , n7407 );
nor ( n7409 , n7405 , n7408 );
xnor ( n7410 , n7400 , n7409 );
not ( n7411 , n7410 );
buf ( n7412 , n7411 );
and ( n7413 , n7372 , n7412 );
not ( n7414 , n7372 );
and ( n7415 , n7414 , n7410 );
nor ( n7416 , n7413 , n7415 );
buf ( n7417 , n7416 );
xnor ( n7418 , n7322 , n7417 );
not ( n7419 , n7418 );
and ( n7420 , n7148 , n7419 );
not ( n7421 , n7148 );
and ( n7422 , n7421 , n7418 );
nor ( n7423 , n7420 , n7422 );
not ( n7424 , n7423 );
not ( n7425 , n7424 );
buf ( n7426 , n4473 );
buf ( n7427 , n7426 );
not ( n7428 , n7427 );
buf ( n7429 , n4474 );
buf ( n7430 , n4475 );
buf ( n7431 , n7430 );
not ( n7432 , n7431 );
buf ( n7433 , n4476 );
not ( n7434 , n7433 );
not ( n7435 , n7434 );
or ( n7436 , n7432 , n7435 );
not ( n7437 , n7430 );
buf ( n7438 , n7433 );
nand ( n7439 , n7437 , n7438 );
nand ( n7440 , n7436 , n7439 );
xor ( n7441 , n7429 , n7440 );
buf ( n7442 , n4477 );
buf ( n7443 , n4478 );
not ( n7444 , n7443 );
xor ( n7445 , n7442 , n7444 );
buf ( n7446 , n4479 );
nand ( n7447 , n7067 , n7446 );
xnor ( n7448 , n7445 , n7447 );
xnor ( n7449 , n7441 , n7448 );
not ( n7450 , n7449 );
not ( n7451 , n7450 );
or ( n7452 , n7428 , n7451 );
not ( n7453 , n7449 );
or ( n7454 , n7453 , n7427 );
nand ( n7455 , n7452 , n7454 );
buf ( n7456 , n4480 );
not ( n7457 , n7456 );
buf ( n7458 , n4481 );
nand ( n7459 , n6514 , n7458 );
buf ( n7460 , n4482 );
buf ( n7461 , n7460 );
and ( n7462 , n7459 , n7461 );
not ( n7463 , n7459 );
not ( n7464 , n7460 );
and ( n7465 , n7463 , n7464 );
nor ( n7466 , n7462 , n7465 );
xor ( n7467 , n7457 , n7466 );
buf ( n7468 , n4483 );
nand ( n7469 , n6828 , n7468 );
buf ( n7470 , n4484 );
buf ( n7471 , n7470 );
and ( n7472 , n7469 , n7471 );
not ( n7473 , n7469 );
not ( n7474 , n7470 );
and ( n7475 , n7473 , n7474 );
nor ( n7476 , n7472 , n7475 );
xnor ( n7477 , n7467 , n7476 );
not ( n7478 , n7477 );
buf ( n7479 , n4485 );
buf ( n7480 , n7479 );
not ( n7481 , n7480 );
buf ( n7482 , n4486 );
not ( n7483 , n7482 );
not ( n7484 , n7483 );
or ( n7485 , n7481 , n7484 );
not ( n7486 , n7479 );
buf ( n7487 , n7482 );
nand ( n7488 , n7486 , n7487 );
nand ( n7489 , n7485 , n7488 );
not ( n7490 , n7489 );
not ( n7491 , n7490 );
and ( n7492 , n7478 , n7491 );
and ( n7493 , n7477 , n7490 );
nor ( n7494 , n7492 , n7493 );
buf ( n7495 , n7494 );
xor ( n7496 , n7455 , n7495 );
not ( n7497 , n7496 );
buf ( n7498 , n4487 );
buf ( n7499 , n7498 );
not ( n7500 , n7499 );
buf ( n7501 , n4488 );
buf ( n7502 , n7501 );
not ( n7503 , n7502 );
buf ( n7504 , n4489 );
not ( n7505 , n7504 );
not ( n7506 , n7505 );
or ( n7507 , n7503 , n7506 );
not ( n7508 , n7501 );
buf ( n7509 , n7504 );
nand ( n7510 , n7508 , n7509 );
nand ( n7511 , n7507 , n7510 );
buf ( n7512 , n4490 );
buf ( n7513 , n7512 );
and ( n7514 , n7511 , n7513 );
not ( n7515 , n7511 );
not ( n7516 , n7512 );
and ( n7517 , n7515 , n7516 );
nor ( n7518 , n7514 , n7517 );
buf ( n7519 , n4491 );
nand ( n7520 , n6634 , n7519 );
buf ( n7521 , n4492 );
buf ( n7522 , n7521 );
and ( n7523 , n7520 , n7522 );
not ( n7524 , n7520 );
not ( n7525 , n7521 );
and ( n7526 , n7524 , n7525 );
nor ( n7527 , n7523 , n7526 );
xor ( n7528 , n7518 , n7527 );
buf ( n7529 , n4493 );
nand ( n7530 , n6515 , n7529 );
buf ( n7531 , n4494 );
buf ( n7532 , n7531 );
and ( n7533 , n7530 , n7532 );
not ( n7534 , n7530 );
not ( n7535 , n7531 );
and ( n7536 , n7534 , n7535 );
nor ( n7537 , n7533 , n7536 );
buf ( n7538 , n7537 );
xnor ( n7539 , n7528 , n7538 );
buf ( n7540 , n7539 );
not ( n7541 , n7540 );
or ( n7542 , n7500 , n7541 );
or ( n7543 , n7540 , n7499 );
nand ( n7544 , n7542 , n7543 );
buf ( n7545 , n4495 );
buf ( n7546 , n7545 );
not ( n7547 , n7546 );
buf ( n7548 , n4496 );
not ( n7549 , n7548 );
not ( n7550 , n7549 );
or ( n7551 , n7547 , n7550 );
not ( n7552 , n7545 );
buf ( n7553 , n7548 );
nand ( n7554 , n7552 , n7553 );
nand ( n7555 , n7551 , n7554 );
buf ( n7556 , n4497 );
buf ( n7557 , n7556 );
and ( n7558 , n7555 , n7557 );
not ( n7559 , n7555 );
not ( n7560 , n7556 );
and ( n7561 , n7559 , n7560 );
nor ( n7562 , n7558 , n7561 );
buf ( n7563 , n6556 );
buf ( n7564 , n4498 );
nand ( n7565 , n7563 , n7564 );
buf ( n7566 , n4499 );
xor ( n7567 , n7565 , n7566 );
xor ( n7568 , n7562 , n7567 );
buf ( n7569 , n6502 );
buf ( n7570 , n4500 );
nand ( n7571 , n7569 , n7570 );
buf ( n7572 , n4501 );
buf ( n7573 , n7572 );
and ( n7574 , n7571 , n7573 );
not ( n7575 , n7571 );
not ( n7576 , n7572 );
and ( n7577 , n7575 , n7576 );
nor ( n7578 , n7574 , n7577 );
xnor ( n7579 , n7568 , n7578 );
buf ( n7580 , n7579 );
and ( n7581 , n7544 , n7580 );
not ( n7582 , n7544 );
not ( n7583 , n7580 );
and ( n7584 , n7582 , n7583 );
nor ( n7585 , n7581 , n7584 );
nand ( n7586 , n7497 , n7585 );
not ( n7587 , n7586 );
buf ( n7588 , n4502 );
buf ( n7589 , n7588 );
not ( n7590 , n7589 );
buf ( n7591 , n4503 );
not ( n7592 , n7591 );
not ( n7593 , n7592 );
or ( n7594 , n7590 , n7593 );
not ( n7595 , n7588 );
buf ( n7596 , n7591 );
nand ( n7597 , n7595 , n7596 );
nand ( n7598 , n7594 , n7597 );
buf ( n7599 , n4504 );
buf ( n7600 , n7599 );
and ( n7601 , n7598 , n7600 );
not ( n7602 , n7598 );
not ( n7603 , n7599 );
and ( n7604 , n7602 , n7603 );
nor ( n7605 , n7601 , n7604 );
buf ( n7606 , n6556 );
buf ( n7607 , n4505 );
nand ( n7608 , n7606 , n7607 );
buf ( n7609 , n4506 );
buf ( n7610 , n7609 );
and ( n7611 , n7608 , n7610 );
not ( n7612 , n7608 );
not ( n7613 , n7609 );
and ( n7614 , n7612 , n7613 );
nor ( n7615 , n7611 , n7614 );
xor ( n7616 , n7605 , n7615 );
buf ( n7617 , n4507 );
nand ( n7618 , n7606 , n7617 );
buf ( n7619 , n4508 );
buf ( n7620 , n7619 );
and ( n7621 , n7618 , n7620 );
not ( n7622 , n7618 );
not ( n7623 , n7619 );
and ( n7624 , n7622 , n7623 );
nor ( n7625 , n7621 , n7624 );
not ( n7626 , n7625 );
xor ( n7627 , n7616 , n7626 );
buf ( n7628 , n4509 );
buf ( n7629 , n7628 );
nand ( n7630 , n7627 , n7629 );
not ( n7631 , n7630 );
nor ( n7632 , n7627 , n7629 );
nor ( n7633 , n7631 , n7632 );
not ( n7634 , n7633 );
buf ( n7635 , n4510 );
buf ( n7636 , n7635 );
not ( n7637 , n7636 );
buf ( n7638 , n4511 );
not ( n7639 , n7638 );
not ( n7640 , n7639 );
or ( n7641 , n7637 , n7640 );
not ( n7642 , n7635 );
buf ( n7643 , n7638 );
nand ( n7644 , n7642 , n7643 );
nand ( n7645 , n7641 , n7644 );
not ( n7646 , n7645 );
not ( n7647 , n7646 );
buf ( n7648 , n4512 );
buf ( n7649 , n4513 );
not ( n7650 , n7649 );
xor ( n7651 , n7648 , n7650 );
buf ( n7652 , n4514 );
nand ( n7653 , n7247 , n7652 );
buf ( n7654 , n4515 );
not ( n7655 , n7654 );
and ( n7656 , n7653 , n7655 );
not ( n7657 , n7653 );
buf ( n7658 , n7654 );
and ( n7659 , n7657 , n7658 );
nor ( n7660 , n7656 , n7659 );
xnor ( n7661 , n7651 , n7660 );
not ( n7662 , n7661 );
or ( n7663 , n7647 , n7662 );
or ( n7664 , n7661 , n7646 );
nand ( n7665 , n7663 , n7664 );
buf ( n7666 , n7665 );
not ( n7667 , n7666 );
or ( n7668 , n7634 , n7667 );
or ( n7669 , n7666 , n7633 );
nand ( n7670 , n7668 , n7669 );
buf ( n7671 , n7670 );
not ( n7672 , n7671 );
and ( n7673 , n7587 , n7672 );
and ( n7674 , n7586 , n7671 );
nor ( n7675 , n7673 , n7674 );
not ( n7676 , n7675 );
not ( n7677 , n7676 );
buf ( n7678 , n4516 );
buf ( n7679 , n7678 );
buf ( n7680 , n4517 );
buf ( n7681 , n7680 );
not ( n7682 , n7681 );
buf ( n7683 , n4518 );
not ( n7684 , n7683 );
not ( n7685 , n7684 );
or ( n7686 , n7682 , n7685 );
not ( n7687 , n7680 );
buf ( n7688 , n7683 );
nand ( n7689 , n7687 , n7688 );
nand ( n7690 , n7686 , n7689 );
buf ( n7691 , n4519 );
buf ( n7692 , n7691 );
and ( n7693 , n7690 , n7692 );
not ( n7694 , n7690 );
not ( n7695 , n7691 );
and ( n7696 , n7694 , n7695 );
nor ( n7697 , n7693 , n7696 );
buf ( n7698 , n6513 );
buf ( n7699 , n4520 );
nand ( n7700 , n7698 , n7699 );
buf ( n7701 , n4521 );
buf ( n7702 , n7701 );
and ( n7703 , n7700 , n7702 );
not ( n7704 , n7700 );
not ( n7705 , n7701 );
and ( n7706 , n7704 , n7705 );
nor ( n7707 , n7703 , n7706 );
xor ( n7708 , n7697 , n7707 );
buf ( n7709 , n7197 );
buf ( n7710 , n4522 );
nand ( n7711 , n7709 , n7710 );
buf ( n7712 , n4523 );
not ( n7713 , n7712 );
and ( n7714 , n7711 , n7713 );
not ( n7715 , n7711 );
buf ( n7716 , n7712 );
and ( n7717 , n7715 , n7716 );
nor ( n7718 , n7714 , n7717 );
xnor ( n7719 , n7708 , n7718 );
buf ( n7720 , n7719 );
xor ( n7721 , n7679 , n7720 );
buf ( n7722 , n4524 );
buf ( n7723 , n4525 );
nand ( n7724 , n6927 , n7723 );
buf ( n7725 , n4526 );
buf ( n7726 , n7725 );
and ( n7727 , n7724 , n7726 );
not ( n7728 , n7724 );
not ( n7729 , n7725 );
and ( n7730 , n7728 , n7729 );
nor ( n7731 , n7727 , n7730 );
xor ( n7732 , n7722 , n7731 );
buf ( n7733 , n4527 );
nand ( n7734 , n7067 , n7733 );
buf ( n7735 , n4528 );
not ( n7736 , n7735 );
and ( n7737 , n7734 , n7736 );
not ( n7738 , n7734 );
buf ( n7739 , n7735 );
and ( n7740 , n7738 , n7739 );
nor ( n7741 , n7737 , n7740 );
xnor ( n7742 , n7732 , n7741 );
not ( n7743 , n7742 );
buf ( n7744 , n4529 );
not ( n7745 , n7744 );
buf ( n7746 , n4530 );
buf ( n7747 , n7746 );
and ( n7748 , n7745 , n7747 );
not ( n7749 , n7745 );
not ( n7750 , n7746 );
and ( n7751 , n7749 , n7750 );
nor ( n7752 , n7748 , n7751 );
not ( n7753 , n7752 );
and ( n7754 , n7743 , n7753 );
and ( n7755 , n7742 , n7752 );
nor ( n7756 , n7754 , n7755 );
xnor ( n7757 , n7721 , n7756 );
not ( n7758 , n7757 );
buf ( n7759 , n4531 );
buf ( n7760 , n7759 );
not ( n7761 , n7760 );
buf ( n7762 , n4532 );
not ( n7763 , n7762 );
buf ( n7764 , n4533 );
buf ( n7765 , n7764 );
not ( n7766 , n7765 );
buf ( n7767 , n4534 );
not ( n7768 , n7767 );
not ( n7769 , n7768 );
or ( n7770 , n7766 , n7769 );
not ( n7771 , n7764 );
buf ( n7772 , n7767 );
nand ( n7773 , n7771 , n7772 );
nand ( n7774 , n7770 , n7773 );
not ( n7775 , n7774 );
xor ( n7776 , n7763 , n7775 );
buf ( n7777 , n4535 );
nand ( n7778 , n7698 , n7777 );
buf ( n7779 , n4536 );
buf ( n7780 , n7779 );
and ( n7781 , n7778 , n7780 );
not ( n7782 , n7778 );
not ( n7783 , n7779 );
and ( n7784 , n7782 , n7783 );
nor ( n7785 , n7781 , n7784 );
not ( n7786 , n7785 );
buf ( n7787 , n6576 );
buf ( n7788 , n4537 );
nand ( n7789 , n7787 , n7788 );
buf ( n7790 , n4538 );
not ( n7791 , n7790 );
and ( n7792 , n7789 , n7791 );
not ( n7793 , n7789 );
buf ( n7794 , n7790 );
and ( n7795 , n7793 , n7794 );
nor ( n7796 , n7792 , n7795 );
not ( n7797 , n7796 );
or ( n7798 , n7786 , n7797 );
or ( n7799 , n7785 , n7796 );
nand ( n7800 , n7798 , n7799 );
xnor ( n7801 , n7776 , n7800 );
not ( n7802 , n7801 );
not ( n7803 , n7802 );
not ( n7804 , n7803 );
or ( n7805 , n7761 , n7804 );
or ( n7806 , n7803 , n7760 );
nand ( n7807 , n7805 , n7806 );
buf ( n7808 , n4539 );
buf ( n7809 , n7808 );
buf ( n7810 , n4540 );
buf ( n7811 , n7810 );
not ( n7812 , n7811 );
buf ( n7813 , n4541 );
not ( n7814 , n7813 );
not ( n7815 , n7814 );
or ( n7816 , n7812 , n7815 );
not ( n7817 , n7810 );
buf ( n7818 , n7813 );
nand ( n7819 , n7817 , n7818 );
nand ( n7820 , n7816 , n7819 );
xor ( n7821 , n7809 , n7820 );
buf ( n7822 , n4542 );
buf ( n7823 , n4543 );
xor ( n7824 , n7822 , n7823 );
buf ( n7825 , n4544 );
nand ( n7826 , n7067 , n7825 );
xnor ( n7827 , n7824 , n7826 );
xnor ( n7828 , n7821 , n7827 );
not ( n7829 , n7828 );
not ( n7830 , n7829 );
and ( n7831 , n7807 , n7830 );
not ( n7832 , n7807 );
buf ( n7833 , n7828 );
not ( n7834 , n7833 );
and ( n7835 , n7832 , n7834 );
nor ( n7836 , n7831 , n7835 );
not ( n7837 , n7836 );
nand ( n7838 , n7758 , n7837 );
not ( n7839 , n7838 );
buf ( n7840 , n4545 );
buf ( n7841 , n7840 );
not ( n7842 , n7841 );
buf ( n7843 , n4546 );
not ( n7844 , n7843 );
not ( n7845 , n7844 );
or ( n7846 , n7842 , n7845 );
not ( n7847 , n7840 );
buf ( n7848 , n7843 );
nand ( n7849 , n7847 , n7848 );
nand ( n7850 , n7846 , n7849 );
buf ( n7851 , n4547 );
buf ( n7852 , n7851 );
and ( n7853 , n7850 , n7852 );
not ( n7854 , n7850 );
not ( n7855 , n7851 );
and ( n7856 , n7854 , n7855 );
nor ( n7857 , n7853 , n7856 );
buf ( n7858 , n4548 );
nand ( n7859 , n6633 , n7858 );
buf ( n7860 , n4549 );
not ( n7861 , n7860 );
and ( n7862 , n7859 , n7861 );
not ( n7863 , n7859 );
buf ( n7864 , n7860 );
and ( n7865 , n7863 , n7864 );
nor ( n7866 , n7862 , n7865 );
xor ( n7867 , n7857 , n7866 );
buf ( n7868 , n6827 );
buf ( n7869 , n4550 );
nand ( n7870 , n7868 , n7869 );
buf ( n7871 , n4551 );
not ( n7872 , n7871 );
and ( n7873 , n7870 , n7872 );
not ( n7874 , n7870 );
buf ( n7875 , n7871 );
and ( n7876 , n7874 , n7875 );
nor ( n7877 , n7873 , n7876 );
xnor ( n7878 , n7867 , n7877 );
buf ( n7879 , n7878 );
not ( n7880 , n7879 );
buf ( n7881 , n4552 );
buf ( n7882 , n7881 );
not ( n7883 , n7882 );
buf ( n7884 , n4553 );
buf ( n7885 , n7884 );
not ( n7886 , n7885 );
buf ( n7887 , n4554 );
not ( n7888 , n7887 );
not ( n7889 , n7888 );
or ( n7890 , n7886 , n7889 );
not ( n7891 , n7884 );
buf ( n7892 , n7887 );
nand ( n7893 , n7891 , n7892 );
nand ( n7894 , n7890 , n7893 );
buf ( n7895 , n4555 );
not ( n7896 , n7895 );
and ( n7897 , n7894 , n7896 );
not ( n7898 , n7894 );
buf ( n7899 , n7895 );
and ( n7900 , n7898 , n7899 );
nor ( n7901 , n7897 , n7900 );
buf ( n7902 , n4556 );
nand ( n7903 , n6828 , n7902 );
buf ( n7904 , n4557 );
not ( n7905 , n7904 );
and ( n7906 , n7903 , n7905 );
not ( n7907 , n7903 );
buf ( n7908 , n7904 );
and ( n7909 , n7907 , n7908 );
nor ( n7910 , n7906 , n7909 );
xor ( n7911 , n7901 , n7910 );
buf ( n7912 , n6645 );
buf ( n7913 , n4558 );
nand ( n7914 , n7912 , n7913 );
buf ( n7915 , n4559 );
not ( n7916 , n7915 );
and ( n7917 , n7914 , n7916 );
not ( n7918 , n7914 );
buf ( n7919 , n7915 );
and ( n7920 , n7918 , n7919 );
nor ( n7921 , n7917 , n7920 );
xnor ( n7922 , n7911 , n7921 );
not ( n7923 , n7922 );
not ( n7924 , n7923 );
or ( n7925 , n7883 , n7924 );
buf ( n7926 , n7922 );
not ( n7927 , n7926 );
or ( n7928 , n7927 , n7882 );
nand ( n7929 , n7925 , n7928 );
not ( n7930 , n7929 );
or ( n7931 , n7880 , n7930 );
or ( n7932 , n7929 , n7879 );
nand ( n7933 , n7931 , n7932 );
not ( n7934 , n7933 );
not ( n7935 , n7934 );
not ( n7936 , n7935 );
and ( n7937 , n7839 , n7936 );
and ( n7938 , n7838 , n7935 );
nor ( n7939 , n7937 , n7938 );
not ( n7940 , n7939 );
or ( n7941 , n7677 , n7940 );
not ( n7942 , n7939 );
nand ( n7943 , n7942 , n7675 );
nand ( n7944 , n7941 , n7943 );
not ( n7945 , n7944 );
and ( n7946 , n7425 , n7945 );
and ( n7947 , n7424 , n7944 );
nor ( n7948 , n7946 , n7947 );
not ( n7949 , n7948 );
or ( n7950 , n6751 , n7949 );
not ( n7951 , n6750 );
not ( n7952 , n7423 );
not ( n7953 , n7944 );
not ( n7954 , n7953 );
or ( n7955 , n7952 , n7954 );
nand ( n7956 , n7424 , n7944 );
nand ( n7957 , n7955 , n7956 );
nand ( n7958 , n7951 , n7957 );
nand ( n7959 , n7950 , n7958 );
buf ( n7960 , n4560 );
not ( n7961 , n7960 );
buf ( n7962 , n4561 );
buf ( n7963 , n7962 );
not ( n7964 , n7963 );
buf ( n7965 , n4562 );
not ( n7966 , n7965 );
not ( n7967 , n7966 );
or ( n7968 , n7964 , n7967 );
not ( n7969 , n7962 );
buf ( n7970 , n7965 );
nand ( n7971 , n7969 , n7970 );
nand ( n7972 , n7968 , n7971 );
xor ( n7973 , n7961 , n7972 );
buf ( n7974 , n4563 );
not ( n7975 , n7974 );
not ( n7976 , n7975 );
buf ( n7977 , n6576 );
buf ( n7978 , n4564 );
nand ( n7979 , n7977 , n7978 );
buf ( n7980 , n4565 );
not ( n7981 , n7980 );
and ( n7982 , n7979 , n7981 );
not ( n7983 , n7979 );
buf ( n7984 , n7980 );
and ( n7985 , n7983 , n7984 );
nor ( n7986 , n7982 , n7985 );
not ( n7987 , n7986 );
or ( n7988 , n7976 , n7987 );
or ( n7989 , n7986 , n7975 );
nand ( n7990 , n7988 , n7989 );
xnor ( n7991 , n7973 , n7990 );
buf ( n7992 , n7991 );
not ( n7993 , n7992 );
buf ( n7994 , n4566 );
nand ( n7995 , n6558 , n7994 );
buf ( n7996 , n4567 );
buf ( n7997 , n7996 );
and ( n7998 , n7995 , n7997 );
not ( n7999 , n7995 );
not ( n8000 , n7996 );
and ( n8001 , n7999 , n8000 );
nor ( n8002 , n7998 , n8001 );
buf ( n8003 , n8002 );
buf ( n8004 , n4568 );
buf ( n8005 , n8004 );
not ( n8006 , n8005 );
buf ( n8007 , n4569 );
not ( n8008 , n8007 );
not ( n8009 , n8008 );
or ( n8010 , n8006 , n8009 );
not ( n8011 , n8004 );
buf ( n8012 , n8007 );
nand ( n8013 , n8011 , n8012 );
nand ( n8014 , n8010 , n8013 );
buf ( n8015 , n4570 );
not ( n8016 , n8015 );
and ( n8017 , n8014 , n8016 );
not ( n8018 , n8014 );
buf ( n8019 , n8015 );
and ( n8020 , n8018 , n8019 );
nor ( n8021 , n8017 , n8020 );
buf ( n8022 , n4571 );
nand ( n8023 , n7698 , n8022 );
buf ( n8024 , n4572 );
buf ( n8025 , n8024 );
and ( n8026 , n8023 , n8025 );
not ( n8027 , n8023 );
not ( n8028 , n8024 );
and ( n8029 , n8027 , n8028 );
nor ( n8030 , n8026 , n8029 );
xor ( n8031 , n8021 , n8030 );
buf ( n8032 , n7698 );
buf ( n8033 , n4573 );
nand ( n8034 , n8032 , n8033 );
buf ( n8035 , n4574 );
not ( n8036 , n8035 );
and ( n8037 , n8034 , n8036 );
not ( n8038 , n8034 );
buf ( n8039 , n8035 );
and ( n8040 , n8038 , n8039 );
nor ( n8041 , n8037 , n8040 );
xnor ( n8042 , n8031 , n8041 );
and ( n8043 , n8003 , n8042 );
not ( n8044 , n8003 );
xor ( n8045 , n8021 , n8030 );
xnor ( n8046 , n8045 , n8041 );
not ( n8047 , n8046 );
and ( n8048 , n8044 , n8047 );
nor ( n8049 , n8043 , n8048 );
xor ( n8050 , n7993 , n8049 );
buf ( n8051 , n4575 );
not ( n8052 , n8051 );
not ( n8053 , n6688 );
buf ( n8054 , n4576 );
not ( n8055 , n8054 );
not ( n8056 , n8055 );
or ( n8057 , n8053 , n8056 );
buf ( n8058 , n8054 );
nand ( n8059 , n6735 , n8058 );
nand ( n8060 , n8057 , n8059 );
buf ( n8061 , n4577 );
not ( n8062 , n8061 );
and ( n8063 , n8060 , n8062 );
not ( n8064 , n8060 );
buf ( n8065 , n8061 );
and ( n8066 , n8064 , n8065 );
nor ( n8067 , n8063 , n8066 );
buf ( n8068 , n6500 );
buf ( n8069 , n8068 );
buf ( n8070 , n8069 );
buf ( n8071 , n4578 );
nand ( n8072 , n8070 , n8071 );
buf ( n8073 , n4579 );
buf ( n8074 , n8073 );
and ( n8075 , n8072 , n8074 );
not ( n8076 , n8072 );
not ( n8077 , n8073 );
and ( n8078 , n8076 , n8077 );
nor ( n8079 , n8075 , n8078 );
xor ( n8080 , n8067 , n8079 );
buf ( n8081 , n4580 );
nand ( n8082 , n7107 , n8081 );
buf ( n8083 , n4581 );
buf ( n8084 , n8083 );
and ( n8085 , n8082 , n8084 );
not ( n8086 , n8082 );
not ( n8087 , n8083 );
and ( n8088 , n8086 , n8087 );
nor ( n8089 , n8085 , n8088 );
not ( n8090 , n8089 );
xnor ( n8091 , n8080 , n8090 );
not ( n8092 , n8091 );
or ( n8093 , n8052 , n8092 );
or ( n8094 , n8091 , n8051 );
nand ( n8095 , n8093 , n8094 );
buf ( n8096 , n4582 );
buf ( n8097 , n8096 );
not ( n8098 , n8097 );
buf ( n8099 , n4583 );
not ( n8100 , n8099 );
not ( n8101 , n8100 );
or ( n8102 , n8098 , n8101 );
not ( n8103 , n8096 );
buf ( n8104 , n8099 );
nand ( n8105 , n8103 , n8104 );
nand ( n8106 , n8102 , n8105 );
buf ( n8107 , n4584 );
buf ( n8108 , n8107 );
and ( n8109 , n8106 , n8108 );
not ( n8110 , n8106 );
not ( n8111 , n8107 );
and ( n8112 , n8110 , n8111 );
nor ( n8113 , n8109 , n8112 );
buf ( n8114 , n4585 );
nand ( n8115 , n6577 , n8114 );
buf ( n8116 , n4586 );
buf ( n8117 , n8116 );
and ( n8118 , n8115 , n8117 );
not ( n8119 , n8115 );
not ( n8120 , n8116 );
and ( n8121 , n8119 , n8120 );
nor ( n8122 , n8118 , n8121 );
xor ( n8123 , n8113 , n8122 );
buf ( n8124 , n6645 );
buf ( n8125 , n8124 );
buf ( n8126 , n4587 );
nand ( n8127 , n8125 , n8126 );
buf ( n8128 , n4588 );
buf ( n8129 , n8128 );
and ( n8130 , n8127 , n8129 );
not ( n8131 , n8127 );
not ( n8132 , n8128 );
and ( n8133 , n8131 , n8132 );
nor ( n8134 , n8130 , n8133 );
xnor ( n8135 , n8123 , n8134 );
not ( n8136 , n8135 );
and ( n8137 , n8095 , n8136 );
not ( n8138 , n8095 );
not ( n8139 , n8135 );
not ( n8140 , n8139 );
and ( n8141 , n8138 , n8140 );
nor ( n8142 , n8137 , n8141 );
nand ( n8143 , n8050 , n8142 );
not ( n8144 , n8143 );
buf ( n8145 , n4589 );
buf ( n8146 , n8145 );
not ( n8147 , n8146 );
buf ( n8148 , n4590 );
buf ( n8149 , n8148 );
not ( n8150 , n8149 );
buf ( n8151 , n4591 );
not ( n8152 , n8151 );
not ( n8153 , n8152 );
or ( n8154 , n8150 , n8153 );
not ( n8155 , n8148 );
buf ( n8156 , n8151 );
nand ( n8157 , n8155 , n8156 );
nand ( n8158 , n8154 , n8157 );
buf ( n8159 , n4592 );
buf ( n8160 , n8159 );
and ( n8161 , n8158 , n8160 );
not ( n8162 , n8158 );
not ( n8163 , n8159 );
and ( n8164 , n8162 , n8163 );
nor ( n8165 , n8161 , n8164 );
buf ( n8166 , n4593 );
nand ( n8167 , n6828 , n8166 );
buf ( n8168 , n4594 );
buf ( n8169 , n8168 );
and ( n8170 , n8167 , n8169 );
not ( n8171 , n8167 );
not ( n8172 , n8168 );
and ( n8173 , n8171 , n8172 );
nor ( n8174 , n8170 , n8173 );
xor ( n8175 , n8165 , n8174 );
buf ( n8176 , n6827 );
buf ( n8177 , n4595 );
nand ( n8178 , n8176 , n8177 );
buf ( n8179 , n4596 );
buf ( n8180 , n8179 );
and ( n8181 , n8178 , n8180 );
not ( n8182 , n8178 );
not ( n8183 , n8179 );
and ( n8184 , n8182 , n8183 );
nor ( n8185 , n8181 , n8184 );
xnor ( n8186 , n8175 , n8185 );
not ( n8187 , n8186 );
or ( n8188 , n8147 , n8187 );
not ( n8189 , n8146 );
xor ( n8190 , n8165 , n8185 );
not ( n8191 , n8174 );
xnor ( n8192 , n8190 , n8191 );
nand ( n8193 , n8189 , n8192 );
nand ( n8194 , n8188 , n8193 );
buf ( n8195 , n4597 );
buf ( n8196 , n8195 );
not ( n8197 , n8196 );
buf ( n8198 , n4598 );
not ( n8199 , n8198 );
not ( n8200 , n8199 );
or ( n8201 , n8197 , n8200 );
not ( n8202 , n8195 );
buf ( n8203 , n8198 );
nand ( n8204 , n8202 , n8203 );
nand ( n8205 , n8201 , n8204 );
buf ( n8206 , n4599 );
not ( n8207 , n8206 );
and ( n8208 , n8205 , n8207 );
not ( n8209 , n8205 );
buf ( n8210 , n8206 );
and ( n8211 , n8209 , n8210 );
nor ( n8212 , n8208 , n8211 );
buf ( n8213 , n4600 );
nand ( n8214 , n7247 , n8213 );
buf ( n8215 , n4601 );
buf ( n8216 , n8215 );
and ( n8217 , n8214 , n8216 );
not ( n8218 , n8214 );
not ( n8219 , n8215 );
and ( n8220 , n8218 , n8219 );
nor ( n8221 , n8217 , n8220 );
xor ( n8222 , n8212 , n8221 );
buf ( n8223 , n7698 );
buf ( n8224 , n4602 );
nand ( n8225 , n8223 , n8224 );
buf ( n8226 , n4603 );
buf ( n8227 , n8226 );
and ( n8228 , n8225 , n8227 );
not ( n8229 , n8225 );
not ( n8230 , n8226 );
and ( n8231 , n8229 , n8230 );
nor ( n8232 , n8228 , n8231 );
xnor ( n8233 , n8222 , n8232 );
buf ( n8234 , n8233 );
and ( n8235 , n8194 , n8234 );
not ( n8236 , n8194 );
not ( n8237 , n8234 );
and ( n8238 , n8236 , n8237 );
nor ( n8239 , n8235 , n8238 );
not ( n8240 , n8239 );
and ( n8241 , n8144 , n8240 );
and ( n8242 , n8143 , n8239 );
nor ( n8243 , n8241 , n8242 );
not ( n8244 , n8243 );
buf ( n8245 , n4604 );
buf ( n8246 , n4605 );
not ( n8247 , n8246 );
buf ( n8248 , n4606 );
buf ( n8249 , n8248 );
and ( n8250 , n8247 , n8249 );
not ( n8251 , n8247 );
not ( n8252 , n8248 );
and ( n8253 , n8251 , n8252 );
nor ( n8254 , n8250 , n8253 );
xor ( n8255 , n8245 , n8254 );
buf ( n8256 , n4607 );
buf ( n8257 , n4608 );
buf ( n8258 , n8257 );
xor ( n8259 , n8256 , n8258 );
buf ( n8260 , n6770 );
buf ( n8261 , n4609 );
nand ( n8262 , n8260 , n8261 );
xnor ( n8263 , n8259 , n8262 );
xnor ( n8264 , n8255 , n8263 );
not ( n8265 , n8264 );
buf ( n8266 , n4610 );
nand ( n8267 , n7067 , n8266 );
buf ( n8268 , n4611 );
buf ( n8269 , n8268 );
and ( n8270 , n8267 , n8269 );
not ( n8271 , n8267 );
not ( n8272 , n8268 );
and ( n8273 , n8271 , n8272 );
nor ( n8274 , n8270 , n8273 );
buf ( n8275 , n8274 );
not ( n8276 , n8275 );
and ( n8277 , n8265 , n8276 );
and ( n8278 , n8264 , n8275 );
nor ( n8279 , n8277 , n8278 );
buf ( n8280 , n4612 );
nand ( n8281 , n7293 , n8280 );
buf ( n8282 , n4613 );
buf ( n8283 , n8282 );
and ( n8284 , n8281 , n8283 );
not ( n8285 , n8281 );
not ( n8286 , n8282 );
and ( n8287 , n8285 , n8286 );
nor ( n8288 , n8284 , n8287 );
xor ( n8289 , n7227 , n8288 );
buf ( n8290 , n4614 );
nand ( n8291 , n7258 , n8290 );
buf ( n8292 , n4615 );
not ( n8293 , n8292 );
and ( n8294 , n8291 , n8293 );
not ( n8295 , n8291 );
buf ( n8296 , n8292 );
and ( n8297 , n8295 , n8296 );
nor ( n8298 , n8294 , n8297 );
xnor ( n8299 , n8289 , n8298 );
not ( n8300 , n8299 );
buf ( n8301 , n4616 );
not ( n8302 , n8301 );
buf ( n8303 , n4617 );
buf ( n8304 , n8303 );
and ( n8305 , n8302 , n8304 );
not ( n8306 , n8302 );
not ( n8307 , n8303 );
and ( n8308 , n8306 , n8307 );
nor ( n8309 , n8305 , n8308 );
not ( n8310 , n8309 );
and ( n8311 , n8300 , n8310 );
and ( n8312 , n8299 , n8309 );
nor ( n8313 , n8311 , n8312 );
buf ( n8314 , n8313 );
and ( n8315 , n8279 , n8314 );
not ( n8316 , n8279 );
not ( n8317 , n8313 );
and ( n8318 , n8316 , n8317 );
nor ( n8319 , n8315 , n8318 );
not ( n8320 , n8319 );
not ( n8321 , n6792 );
buf ( n8322 , n6513 );
buf ( n8323 , n8322 );
buf ( n8324 , n4618 );
nand ( n8325 , n8323 , n8324 );
buf ( n8326 , n4619 );
not ( n8327 , n8326 );
and ( n8328 , n8325 , n8327 );
not ( n8329 , n8325 );
buf ( n8330 , n8326 );
and ( n8331 , n8329 , n8330 );
nor ( n8332 , n8328 , n8331 );
not ( n8333 , n8332 );
not ( n8334 , n6839 );
or ( n8335 , n8333 , n8334 );
not ( n8336 , n8332 );
nand ( n8337 , n8336 , n6844 );
nand ( n8338 , n8335 , n8337 );
not ( n8339 , n8338 );
or ( n8340 , n8321 , n8339 );
or ( n8341 , n8338 , n6792 );
nand ( n8342 , n8340 , n8341 );
nand ( n8343 , n8320 , n8342 );
buf ( n8344 , n4620 );
not ( n8345 , n8344 );
buf ( n8346 , n4621 );
buf ( n8347 , n8346 );
not ( n8348 , n8347 );
buf ( n8349 , n4622 );
not ( n8350 , n8349 );
not ( n8351 , n8350 );
or ( n8352 , n8348 , n8351 );
not ( n8353 , n8346 );
buf ( n8354 , n8349 );
nand ( n8355 , n8353 , n8354 );
nand ( n8356 , n8352 , n8355 );
buf ( n8357 , n4623 );
not ( n8358 , n8357 );
and ( n8359 , n8356 , n8358 );
not ( n8360 , n8356 );
buf ( n8361 , n8357 );
and ( n8362 , n8360 , n8361 );
nor ( n8363 , n8359 , n8362 );
buf ( n8364 , n6718 );
buf ( n8365 , n4624 );
nand ( n8366 , n8364 , n8365 );
buf ( n8367 , n4625 );
buf ( n8368 , n8367 );
and ( n8369 , n8366 , n8368 );
not ( n8370 , n8366 );
not ( n8371 , n8367 );
and ( n8372 , n8370 , n8371 );
nor ( n8373 , n8369 , n8372 );
xor ( n8374 , n8363 , n8373 );
buf ( n8375 , n8069 );
buf ( n8376 , n4626 );
nand ( n8377 , n8375 , n8376 );
buf ( n8378 , n4627 );
not ( n8379 , n8378 );
and ( n8380 , n8377 , n8379 );
not ( n8381 , n8377 );
buf ( n8382 , n8378 );
and ( n8383 , n8381 , n8382 );
nor ( n8384 , n8380 , n8383 );
xnor ( n8385 , n8374 , n8384 );
not ( n8386 , n8385 );
or ( n8387 , n8345 , n8386 );
not ( n8388 , n8344 );
not ( n8389 , n8373 );
not ( n8390 , n8384 );
or ( n8391 , n8389 , n8390 );
or ( n8392 , n8373 , n8384 );
nand ( n8393 , n8391 , n8392 );
not ( n8394 , n8363 );
and ( n8395 , n8393 , n8394 );
not ( n8396 , n8393 );
and ( n8397 , n8396 , n8363 );
nor ( n8398 , n8395 , n8397 );
nand ( n8399 , n8388 , n8398 );
nand ( n8400 , n8387 , n8399 );
buf ( n8401 , n4628 );
buf ( n8402 , n8401 );
not ( n8403 , n8402 );
buf ( n8404 , n4629 );
not ( n8405 , n8404 );
not ( n8406 , n8405 );
or ( n8407 , n8403 , n8406 );
not ( n8408 , n8401 );
buf ( n8409 , n8404 );
nand ( n8410 , n8408 , n8409 );
nand ( n8411 , n8407 , n8410 );
buf ( n8412 , n4630 );
not ( n8413 , n8412 );
and ( n8414 , n8411 , n8413 );
not ( n8415 , n8411 );
buf ( n8416 , n8412 );
and ( n8417 , n8415 , n8416 );
nor ( n8418 , n8414 , n8417 );
buf ( n8419 , n4631 );
nand ( n8420 , n7107 , n8419 );
buf ( n8421 , n4632 );
buf ( n8422 , n8421 );
and ( n8423 , n8420 , n8422 );
not ( n8424 , n8420 );
not ( n8425 , n8421 );
and ( n8426 , n8424 , n8425 );
nor ( n8427 , n8423 , n8426 );
xor ( n8428 , n8418 , n8427 );
buf ( n8429 , n4633 );
nand ( n8430 , n7912 , n8429 );
buf ( n8431 , n4634 );
buf ( n8432 , n8431 );
and ( n8433 , n8430 , n8432 );
not ( n8434 , n8430 );
not ( n8435 , n8431 );
and ( n8436 , n8434 , n8435 );
nor ( n8437 , n8433 , n8436 );
xor ( n8438 , n8428 , n8437 );
buf ( n8439 , n8438 );
not ( n8440 , n8439 );
and ( n8441 , n8400 , n8440 );
not ( n8442 , n8400 );
and ( n8443 , n8442 , n8439 );
nor ( n8444 , n8441 , n8443 );
not ( n8445 , n8444 );
and ( n8446 , n8343 , n8445 );
not ( n8447 , n8343 );
and ( n8448 , n8447 , n8444 );
nor ( n8449 , n8446 , n8448 );
not ( n8450 , n8449 );
or ( n8451 , n8244 , n8450 );
or ( n8452 , n8449 , n8243 );
nand ( n8453 , n8451 , n8452 );
buf ( n8454 , n6513 );
buf ( n8455 , n8454 );
buf ( n8456 , n4635 );
nand ( n8457 , n8455 , n8456 );
buf ( n8458 , n4636 );
buf ( n8459 , n8458 );
and ( n8460 , n8457 , n8459 );
not ( n8461 , n8457 );
not ( n8462 , n8458 );
and ( n8463 , n8461 , n8462 );
nor ( n8464 , n8460 , n8463 );
not ( n8465 , n8464 );
buf ( n8466 , n4637 );
buf ( n8467 , n8466 );
not ( n8468 , n8467 );
buf ( n8469 , n4638 );
not ( n8470 , n8469 );
not ( n8471 , n8470 );
or ( n8472 , n8468 , n8471 );
not ( n8473 , n8466 );
buf ( n8474 , n8469 );
nand ( n8475 , n8473 , n8474 );
nand ( n8476 , n8472 , n8475 );
buf ( n8477 , n4639 );
buf ( n8478 , n8477 );
and ( n8479 , n8476 , n8478 );
not ( n8480 , n8476 );
not ( n8481 , n8477 );
and ( n8482 , n8480 , n8481 );
nor ( n8483 , n8479 , n8482 );
buf ( n8484 , n4640 );
nand ( n8485 , n6916 , n8484 );
buf ( n8486 , n4641 );
buf ( n8487 , n8486 );
and ( n8488 , n8485 , n8487 );
not ( n8489 , n8485 );
not ( n8490 , n8486 );
and ( n8491 , n8489 , n8490 );
nor ( n8492 , n8488 , n8491 );
xor ( n8493 , n8483 , n8492 );
buf ( n8494 , n4642 );
nand ( n8495 , n6927 , n8494 );
buf ( n8496 , n4643 );
buf ( n8497 , n8496 );
and ( n8498 , n8495 , n8497 );
not ( n8499 , n8495 );
not ( n8500 , n8496 );
and ( n8501 , n8499 , n8500 );
nor ( n8502 , n8498 , n8501 );
not ( n8503 , n8502 );
xnor ( n8504 , n8493 , n8503 );
not ( n8505 , n8504 );
or ( n8506 , n8465 , n8505 );
or ( n8507 , n8504 , n8464 );
nand ( n8508 , n8506 , n8507 );
buf ( n8509 , n4644 );
buf ( n8510 , n8509 );
not ( n8511 , n8510 );
buf ( n8512 , n4645 );
not ( n8513 , n8512 );
not ( n8514 , n8513 );
or ( n8515 , n8511 , n8514 );
not ( n8516 , n8509 );
buf ( n8517 , n8512 );
nand ( n8518 , n8516 , n8517 );
nand ( n8519 , n8515 , n8518 );
buf ( n8520 , n4646 );
not ( n8521 , n8520 );
and ( n8522 , n8519 , n8521 );
not ( n8523 , n8519 );
buf ( n8524 , n8520 );
and ( n8525 , n8523 , n8524 );
nor ( n8526 , n8522 , n8525 );
buf ( n8527 , n4647 );
nand ( n8528 , n6770 , n8527 );
buf ( n8529 , n4648 );
buf ( n8530 , n8529 );
and ( n8531 , n8528 , n8530 );
not ( n8532 , n8528 );
not ( n8533 , n8529 );
and ( n8534 , n8532 , n8533 );
nor ( n8535 , n8531 , n8534 );
xor ( n8536 , n8526 , n8535 );
buf ( n8537 , n8068 );
buf ( n8538 , n4649 );
nand ( n8539 , n8537 , n8538 );
buf ( n8540 , n4650 );
not ( n8541 , n8540 );
and ( n8542 , n8539 , n8541 );
not ( n8543 , n8539 );
buf ( n8544 , n8540 );
and ( n8545 , n8543 , n8544 );
nor ( n8546 , n8542 , n8545 );
xnor ( n8547 , n8536 , n8546 );
buf ( n8548 , n8547 );
not ( n8549 , n8548 );
and ( n8550 , n8508 , n8549 );
not ( n8551 , n8508 );
and ( n8552 , n8551 , n8548 );
nor ( n8553 , n8550 , n8552 );
not ( n8554 , n8553 );
buf ( n8555 , n4651 );
nand ( n8556 , n6557 , n8555 );
buf ( n8557 , n4652 );
buf ( n8558 , n8557 );
and ( n8559 , n8556 , n8558 );
not ( n8560 , n8556 );
not ( n8561 , n8557 );
and ( n8562 , n8560 , n8561 );
nor ( n8563 , n8559 , n8562 );
buf ( n8564 , n8563 );
not ( n8565 , n8564 );
not ( n8566 , n7802 );
or ( n8567 , n8565 , n8566 );
buf ( n8568 , n7801 );
not ( n8569 , n8568 );
or ( n8570 , n8569 , n8564 );
nand ( n8571 , n8567 , n8570 );
not ( n8572 , n8571 );
not ( n8573 , n7833 );
and ( n8574 , n8572 , n8573 );
and ( n8575 , n8571 , n7830 );
nor ( n8576 , n8574 , n8575 );
not ( n8577 , n8576 );
nand ( n8578 , n8554 , n8577 );
buf ( n8579 , n4653 );
buf ( n8580 , n8579 );
not ( n8581 , n8580 );
buf ( n8582 , n4654 );
buf ( n8583 , n8582 );
not ( n8584 , n8583 );
not ( n8585 , n6954 );
or ( n8586 , n8584 , n8585 );
not ( n8587 , n8582 );
buf ( n8588 , n6953 );
nand ( n8589 , n8587 , n8588 );
nand ( n8590 , n8586 , n8589 );
buf ( n8591 , n4655 );
not ( n8592 , n8591 );
and ( n8593 , n8590 , n8592 );
not ( n8594 , n8590 );
buf ( n8595 , n8591 );
and ( n8596 , n8594 , n8595 );
nor ( n8597 , n8593 , n8596 );
buf ( n8598 , n4656 );
nand ( n8599 , n7107 , n8598 );
buf ( n8600 , n4657 );
buf ( n8601 , n8600 );
and ( n8602 , n8599 , n8601 );
not ( n8603 , n8599 );
not ( n8604 , n8600 );
and ( n8605 , n8603 , n8604 );
nor ( n8606 , n8602 , n8605 );
xor ( n8607 , n8597 , n8606 );
buf ( n8608 , n6815 );
buf ( n8609 , n4658 );
nand ( n8610 , n8608 , n8609 );
buf ( n8611 , n4659 );
not ( n8612 , n8611 );
and ( n8613 , n8610 , n8612 );
not ( n8614 , n8610 );
buf ( n8615 , n8611 );
and ( n8616 , n8614 , n8615 );
nor ( n8617 , n8613 , n8616 );
xnor ( n8618 , n8607 , n8617 );
buf ( n8619 , n8618 );
buf ( n8620 , n8619 );
not ( n8621 , n8620 );
or ( n8622 , n8581 , n8621 );
or ( n8623 , n8620 , n8580 );
nand ( n8624 , n8622 , n8623 );
buf ( n8625 , n4660 );
buf ( n8626 , n8625 );
not ( n8627 , n8626 );
buf ( n8628 , n4661 );
not ( n8629 , n8628 );
not ( n8630 , n8629 );
or ( n8631 , n8627 , n8630 );
not ( n8632 , n8625 );
buf ( n8633 , n8628 );
nand ( n8634 , n8632 , n8633 );
nand ( n8635 , n8631 , n8634 );
buf ( n8636 , n4662 );
not ( n8637 , n8636 );
and ( n8638 , n8635 , n8637 );
not ( n8639 , n8635 );
buf ( n8640 , n8636 );
and ( n8641 , n8639 , n8640 );
nor ( n8642 , n8638 , n8641 );
buf ( n8643 , n4663 );
nand ( n8644 , n6927 , n8643 );
buf ( n8645 , n4664 );
buf ( n8646 , n8645 );
and ( n8647 , n8644 , n8646 );
not ( n8648 , n8644 );
not ( n8649 , n8645 );
and ( n8650 , n8648 , n8649 );
nor ( n8651 , n8647 , n8650 );
xor ( n8652 , n8642 , n8651 );
buf ( n8653 , n4665 );
nand ( n8654 , n8455 , n8653 );
buf ( n8655 , n4666 );
buf ( n8656 , n8655 );
and ( n8657 , n8654 , n8656 );
not ( n8658 , n8654 );
not ( n8659 , n8655 );
and ( n8660 , n8658 , n8659 );
nor ( n8661 , n8657 , n8660 );
xnor ( n8662 , n8652 , n8661 );
not ( n8663 , n8662 );
xor ( n8664 , n8624 , n8663 );
and ( n8665 , n8578 , n8664 );
not ( n8666 , n8578 );
not ( n8667 , n8664 );
and ( n8668 , n8666 , n8667 );
nor ( n8669 , n8665 , n8668 );
and ( n8670 , n8453 , n8669 );
not ( n8671 , n8453 );
not ( n8672 , n8669 );
and ( n8673 , n8671 , n8672 );
nor ( n8674 , n8670 , n8673 );
buf ( n8675 , n6871 );
buf ( n8676 , n4667 );
nand ( n8677 , n8675 , n8676 );
buf ( n8678 , n4668 );
not ( n8679 , n8678 );
and ( n8680 , n8677 , n8679 );
not ( n8681 , n8677 );
buf ( n8682 , n8678 );
and ( n8683 , n8681 , n8682 );
nor ( n8684 , n8680 , n8683 );
buf ( n8685 , n4669 );
buf ( n8686 , n8685 );
not ( n8687 , n8686 );
buf ( n8688 , n4670 );
not ( n8689 , n8688 );
not ( n8690 , n8689 );
or ( n8691 , n8687 , n8690 );
not ( n8692 , n8685 );
buf ( n8693 , n8688 );
nand ( n8694 , n8692 , n8693 );
nand ( n8695 , n8691 , n8694 );
buf ( n8696 , n4671 );
buf ( n8697 , n8696 );
and ( n8698 , n8695 , n8697 );
not ( n8699 , n8695 );
not ( n8700 , n8696 );
and ( n8701 , n8699 , n8700 );
nor ( n8702 , n8698 , n8701 );
buf ( n8703 , n4672 );
nand ( n8704 , n8176 , n8703 );
buf ( n8705 , n4673 );
buf ( n8706 , n8705 );
and ( n8707 , n8704 , n8706 );
not ( n8708 , n8704 );
not ( n8709 , n8705 );
and ( n8710 , n8708 , n8709 );
nor ( n8711 , n8707 , n8710 );
xor ( n8712 , n8702 , n8711 );
buf ( n8713 , n4674 );
nand ( n8714 , n6558 , n8713 );
buf ( n8715 , n4675 );
not ( n8716 , n8715 );
and ( n8717 , n8714 , n8716 );
not ( n8718 , n8714 );
buf ( n8719 , n8715 );
and ( n8720 , n8718 , n8719 );
nor ( n8721 , n8717 , n8720 );
xnor ( n8722 , n8712 , n8721 );
buf ( n8723 , n8722 );
not ( n8724 , n8723 );
xor ( n8725 , n8684 , n8724 );
buf ( n8726 , n4676 );
not ( n8727 , n8726 );
buf ( n8728 , n4677 );
buf ( n8729 , n8728 );
and ( n8730 , n8727 , n8729 );
not ( n8731 , n8727 );
not ( n8732 , n8728 );
and ( n8733 , n8731 , n8732 );
nor ( n8734 , n8730 , n8733 );
not ( n8735 , n8734 );
buf ( n8736 , n4678 );
buf ( n8737 , n4679 );
nand ( n8738 , n7698 , n8737 );
buf ( n8739 , n4680 );
buf ( n8740 , n8739 );
and ( n8741 , n8738 , n8740 );
not ( n8742 , n8738 );
not ( n8743 , n8739 );
and ( n8744 , n8742 , n8743 );
nor ( n8745 , n8741 , n8744 );
xor ( n8746 , n8736 , n8745 );
buf ( n8747 , n4681 );
nand ( n8748 , n6828 , n8747 );
buf ( n8749 , n4682 );
not ( n8750 , n8749 );
and ( n8751 , n8748 , n8750 );
not ( n8752 , n8748 );
buf ( n8753 , n8749 );
and ( n8754 , n8752 , n8753 );
nor ( n8755 , n8751 , n8754 );
xnor ( n8756 , n8746 , n8755 );
not ( n8757 , n8756 );
or ( n8758 , n8735 , n8757 );
or ( n8759 , n8756 , n8734 );
nand ( n8760 , n8758 , n8759 );
buf ( n8761 , n8760 );
not ( n8762 , n8761 );
xnor ( n8763 , n8725 , n8762 );
buf ( n8764 , n4683 );
buf ( n8765 , n4684 );
buf ( n8766 , n8765 );
not ( n8767 , n8766 );
buf ( n8768 , n4685 );
not ( n8769 , n8768 );
not ( n8770 , n8769 );
or ( n8771 , n8767 , n8770 );
not ( n8772 , n8765 );
buf ( n8773 , n8768 );
nand ( n8774 , n8772 , n8773 );
nand ( n8775 , n8771 , n8774 );
xor ( n8776 , n8764 , n8775 );
buf ( n8777 , n4686 );
not ( n8778 , n8777 );
buf ( n8779 , n4687 );
xor ( n8780 , n8778 , n8779 );
buf ( n8781 , n6827 );
buf ( n8782 , n4688 );
nand ( n8783 , n8781 , n8782 );
xnor ( n8784 , n8780 , n8783 );
xnor ( n8785 , n8776 , n8784 );
buf ( n8786 , n8785 );
not ( n8787 , n8786 );
buf ( n8788 , n4689 );
nand ( n8789 , n7606 , n8788 );
buf ( n8790 , n4690 );
buf ( n8791 , n8790 );
and ( n8792 , n8789 , n8791 );
not ( n8793 , n8789 );
not ( n8794 , n8790 );
and ( n8795 , n8793 , n8794 );
nor ( n8796 , n8792 , n8795 );
buf ( n8797 , n8796 );
not ( n8798 , n8797 );
and ( n8799 , n8787 , n8798 );
and ( n8800 , n8786 , n8797 );
nor ( n8801 , n8799 , n8800 );
buf ( n8802 , n4691 );
buf ( n8803 , n8802 );
not ( n8804 , n8803 );
buf ( n8805 , n4692 );
not ( n8806 , n8805 );
not ( n8807 , n8806 );
or ( n8808 , n8804 , n8807 );
not ( n8809 , n8802 );
buf ( n8810 , n8805 );
nand ( n8811 , n8809 , n8810 );
nand ( n8812 , n8808 , n8811 );
not ( n8813 , n8812 );
buf ( n8814 , n4693 );
not ( n8815 , n8814 );
buf ( n8816 , n4694 );
nand ( n8817 , n6815 , n8816 );
not ( n8818 , n8817 );
buf ( n8819 , n4695 );
not ( n8820 , n8819 );
and ( n8821 , n8818 , n8820 );
nand ( n8822 , n8537 , n8816 );
and ( n8823 , n8822 , n8819 );
nor ( n8824 , n8821 , n8823 );
xor ( n8825 , n8815 , n8824 );
buf ( n8826 , n4696 );
nand ( n8827 , n7247 , n8826 );
not ( n8828 , n8827 );
buf ( n8829 , n4697 );
not ( n8830 , n8829 );
and ( n8831 , n8828 , n8830 );
nand ( n8832 , n8375 , n8826 );
and ( n8833 , n8832 , n8829 );
nor ( n8834 , n8831 , n8833 );
xnor ( n8835 , n8825 , n8834 );
not ( n8836 , n8835 );
not ( n8837 , n8836 );
or ( n8838 , n8813 , n8837 );
not ( n8839 , n8812 );
nand ( n8840 , n8839 , n8835 );
nand ( n8841 , n8838 , n8840 );
buf ( n8842 , n8841 );
not ( n8843 , n8842 );
and ( n8844 , n8801 , n8843 );
not ( n8845 , n8801 );
and ( n8846 , n8845 , n8842 );
nor ( n8847 , n8844 , n8846 );
nand ( n8848 , n8763 , n8847 );
buf ( n8849 , n4698 );
buf ( n8850 , n8849 );
not ( n8851 , n8850 );
buf ( n8852 , n4699 );
not ( n8853 , n8852 );
not ( n8854 , n8853 );
or ( n8855 , n8851 , n8854 );
not ( n8856 , n8849 );
buf ( n8857 , n8852 );
nand ( n8858 , n8856 , n8857 );
nand ( n8859 , n8855 , n8858 );
buf ( n8860 , n4700 );
buf ( n8861 , n8860 );
and ( n8862 , n8859 , n8861 );
not ( n8863 , n8859 );
not ( n8864 , n8860 );
and ( n8865 , n8863 , n8864 );
nor ( n8866 , n8862 , n8865 );
buf ( n8867 , n4701 );
nand ( n8868 , n7107 , n8867 );
buf ( n8869 , n4702 );
buf ( n8870 , n8869 );
and ( n8871 , n8868 , n8870 );
not ( n8872 , n8868 );
not ( n8873 , n8869 );
and ( n8874 , n8872 , n8873 );
nor ( n8875 , n8871 , n8874 );
xor ( n8876 , n8866 , n8875 );
buf ( n8877 , n4703 );
nand ( n8878 , n7355 , n8877 );
buf ( n8879 , n4704 );
buf ( n8880 , n8879 );
and ( n8881 , n8878 , n8880 );
not ( n8882 , n8878 );
not ( n8883 , n8879 );
and ( n8884 , n8882 , n8883 );
nor ( n8885 , n8881 , n8884 );
not ( n8886 , n8885 );
xnor ( n8887 , n8876 , n8886 );
not ( n8888 , n8887 );
buf ( n8889 , n4705 );
buf ( n8890 , n8889 );
nor ( n8891 , n8888 , n8890 );
not ( n8892 , n8891 );
nand ( n8893 , n8888 , n8890 );
nand ( n8894 , n8892 , n8893 );
buf ( n8895 , n4706 );
buf ( n8896 , n4707 );
not ( n8897 , n8896 );
buf ( n8898 , n4708 );
buf ( n8899 , n8898 );
and ( n8900 , n8897 , n8899 );
not ( n8901 , n8897 );
not ( n8902 , n8898 );
and ( n8903 , n8901 , n8902 );
nor ( n8904 , n8900 , n8903 );
xor ( n8905 , n8895 , n8904 );
buf ( n8906 , n4709 );
buf ( n8907 , n8906 );
buf ( n8908 , n4710 );
xor ( n8909 , n8907 , n8908 );
buf ( n8910 , n4711 );
nand ( n8911 , n6719 , n8910 );
xnor ( n8912 , n8909 , n8911 );
xnor ( n8913 , n8905 , n8912 );
and ( n8914 , n8894 , n8913 );
not ( n8915 , n8894 );
not ( n8916 , n8913 );
and ( n8917 , n8915 , n8916 );
nor ( n8918 , n8914 , n8917 );
not ( n8919 , n8918 );
and ( n8920 , n8848 , n8919 );
not ( n8921 , n8848 );
and ( n8922 , n8921 , n8918 );
nor ( n8923 , n8920 , n8922 );
not ( n8924 , n8923 );
buf ( n8925 , n4712 );
nand ( n8926 , n7787 , n8925 );
buf ( n8927 , n4713 );
buf ( n8928 , n8927 );
and ( n8929 , n8926 , n8928 );
not ( n8930 , n8926 );
not ( n8931 , n8927 );
and ( n8932 , n8930 , n8931 );
nor ( n8933 , n8929 , n8932 );
buf ( n8934 , n8933 );
not ( n8935 , n8934 );
buf ( n8936 , n4714 );
buf ( n8937 , n8936 );
not ( n8938 , n8937 );
buf ( n8939 , n4715 );
not ( n8940 , n8939 );
not ( n8941 , n8940 );
or ( n8942 , n8938 , n8941 );
not ( n8943 , n8936 );
buf ( n8944 , n8939 );
nand ( n8945 , n8943 , n8944 );
nand ( n8946 , n8942 , n8945 );
buf ( n8947 , n4716 );
buf ( n8948 , n8947 );
and ( n8949 , n8946 , n8948 );
not ( n8950 , n8946 );
not ( n8951 , n8947 );
and ( n8952 , n8950 , n8951 );
nor ( n8953 , n8949 , n8952 );
buf ( n8954 , n8322 );
buf ( n8955 , n4717 );
nand ( n8956 , n8954 , n8955 );
buf ( n8957 , n4718 );
buf ( n8958 , n8957 );
and ( n8959 , n8956 , n8958 );
not ( n8960 , n8956 );
not ( n8961 , n8957 );
and ( n8962 , n8960 , n8961 );
nor ( n8963 , n8959 , n8962 );
buf ( n8964 , n8963 );
xor ( n8965 , n8953 , n8964 );
buf ( n8966 , n6827 );
buf ( n8967 , n4719 );
nand ( n8968 , n8966 , n8967 );
buf ( n8969 , n4720 );
not ( n8970 , n8969 );
and ( n8971 , n8968 , n8970 );
not ( n8972 , n8968 );
buf ( n8973 , n8969 );
and ( n8974 , n8972 , n8973 );
nor ( n8975 , n8971 , n8974 );
buf ( n8976 , n8975 );
xnor ( n8977 , n8965 , n8976 );
buf ( n8978 , n8977 );
not ( n8979 , n8978 );
or ( n8980 , n8935 , n8979 );
or ( n8981 , n8978 , n8934 );
nand ( n8982 , n8980 , n8981 );
xor ( n8983 , n7518 , n7537 );
not ( n8984 , n7527 );
xnor ( n8985 , n8983 , n8984 );
buf ( n8986 , n8985 );
and ( n8987 , n8982 , n8986 );
not ( n8988 , n8982 );
and ( n8989 , n8988 , n7540 );
nor ( n8990 , n8987 , n8989 );
not ( n8991 , n8298 );
buf ( n8992 , n7270 );
not ( n8993 , n8992 );
or ( n8994 , n8991 , n8993 );
not ( n8995 , n8298 );
not ( n8996 , n8992 );
nand ( n8997 , n8995 , n8996 );
nand ( n8998 , n8994 , n8997 );
and ( n8999 , n8998 , n7315 );
not ( n9000 , n8998 );
not ( n9001 , n7315 );
and ( n9002 , n9000 , n9001 );
nor ( n9003 , n8999 , n9002 );
and ( n9004 , n8990 , n9003 );
buf ( n9005 , n4721 );
buf ( n9006 , n9005 );
buf ( n9007 , n4722 );
buf ( n9008 , n9007 );
not ( n9009 , n9008 );
buf ( n9010 , n4723 );
not ( n9011 , n9010 );
not ( n9012 , n9011 );
or ( n9013 , n9009 , n9012 );
not ( n9014 , n9007 );
buf ( n9015 , n9010 );
nand ( n9016 , n9014 , n9015 );
nand ( n9017 , n9013 , n9016 );
buf ( n9018 , n4724 );
buf ( n9019 , n9018 );
and ( n9020 , n9017 , n9019 );
not ( n9021 , n9017 );
not ( n9022 , n9018 );
and ( n9023 , n9021 , n9022 );
nor ( n9024 , n9020 , n9023 );
buf ( n9025 , n4725 );
nand ( n9026 , n8124 , n9025 );
buf ( n9027 , n4726 );
buf ( n9028 , n9027 );
and ( n9029 , n9026 , n9028 );
not ( n9030 , n9026 );
not ( n9031 , n9027 );
and ( n9032 , n9030 , n9031 );
nor ( n9033 , n9029 , n9032 );
xor ( n9034 , n9024 , n9033 );
buf ( n9035 , n4727 );
nand ( n9036 , n7202 , n9035 );
buf ( n9037 , n4728 );
not ( n9038 , n9037 );
and ( n9039 , n9036 , n9038 );
not ( n9040 , n9036 );
buf ( n9041 , n9037 );
and ( n9042 , n9040 , n9041 );
nor ( n9043 , n9039 , n9042 );
buf ( n9044 , n9043 );
xnor ( n9045 , n9034 , n9044 );
buf ( n9046 , n9045 );
xor ( n9047 , n9006 , n9046 );
buf ( n9048 , n4729 );
not ( n9049 , n9048 );
buf ( n9050 , n4730 );
not ( n9051 , n9050 );
buf ( n9052 , n4731 );
buf ( n9053 , n9052 );
nand ( n9054 , n9051 , n9053 );
not ( n9055 , n9052 );
buf ( n9056 , n9050 );
nand ( n9057 , n9055 , n9056 );
and ( n9058 , n9054 , n9057 );
xor ( n9059 , n9049 , n9058 );
buf ( n9060 , n4732 );
buf ( n9061 , n4733 );
xor ( n9062 , n9060 , n9061 );
buf ( n9063 , n4734 );
nand ( n9064 , n7569 , n9063 );
xnor ( n9065 , n9062 , n9064 );
xnor ( n9066 , n9059 , n9065 );
buf ( n9067 , n9066 );
xnor ( n9068 , n9047 , n9067 );
not ( n9069 , n9068 );
and ( n9070 , n9004 , n9069 );
not ( n9071 , n9004 );
and ( n9072 , n9071 , n9068 );
nor ( n9073 , n9070 , n9072 );
not ( n9074 , n9073 );
and ( n9075 , n8924 , n9074 );
and ( n9076 , n8923 , n9073 );
nor ( n9077 , n9075 , n9076 );
and ( n9078 , n8674 , n9077 );
not ( n9079 , n8674 );
not ( n9080 , n9077 );
and ( n9081 , n9079 , n9080 );
nor ( n9082 , n9078 , n9081 );
buf ( n9083 , n9082 );
and ( n9084 , n7959 , n9083 );
not ( n9085 , n7959 );
not ( n9086 , n9077 );
not ( n9087 , n8674 );
or ( n9088 , n9086 , n9087 );
not ( n9089 , n8674 );
nand ( n9090 , n9089 , n9080 );
nand ( n9091 , n9088 , n9090 );
buf ( n9092 , n9091 );
and ( n9093 , n9085 , n9092 );
nor ( n9094 , n9084 , n9093 );
not ( n9095 , n9094 );
buf ( n9096 , n4735 );
buf ( n9097 , n9096 );
buf ( n9098 , n4736 );
buf ( n9099 , n9098 );
not ( n9100 , n9099 );
buf ( n9101 , n4737 );
not ( n9102 , n9101 );
not ( n9103 , n9102 );
or ( n9104 , n9100 , n9103 );
not ( n9105 , n9098 );
buf ( n9106 , n9101 );
nand ( n9107 , n9105 , n9106 );
nand ( n9108 , n9104 , n9107 );
buf ( n9109 , n4738 );
not ( n9110 , n9109 );
and ( n9111 , n9108 , n9110 );
not ( n9112 , n9108 );
buf ( n9113 , n9109 );
and ( n9114 , n9112 , n9113 );
nor ( n9115 , n9111 , n9114 );
buf ( n9116 , n4739 );
nand ( n9117 , n7698 , n9116 );
buf ( n9118 , n4740 );
buf ( n9119 , n9118 );
and ( n9120 , n9117 , n9119 );
not ( n9121 , n9117 );
not ( n9122 , n9118 );
and ( n9123 , n9121 , n9122 );
nor ( n9124 , n9120 , n9123 );
xor ( n9125 , n9115 , n9124 );
buf ( n9126 , n4741 );
nand ( n9127 , n8781 , n9126 );
buf ( n9128 , n4742 );
buf ( n9129 , n9128 );
and ( n9130 , n9127 , n9129 );
not ( n9131 , n9127 );
not ( n9132 , n9128 );
and ( n9133 , n9131 , n9132 );
nor ( n9134 , n9130 , n9133 );
xnor ( n9135 , n9125 , n9134 );
buf ( n9136 , n9135 );
not ( n9137 , n9136 );
and ( n9138 , n9097 , n9137 );
not ( n9139 , n9097 );
and ( n9140 , n9139 , n9136 );
or ( n9141 , n9138 , n9140 );
buf ( n9142 , n4743 );
buf ( n9143 , n9142 );
not ( n9144 , n9143 );
buf ( n9145 , n4744 );
not ( n9146 , n9145 );
not ( n9147 , n9146 );
or ( n9148 , n9144 , n9147 );
not ( n9149 , n9142 );
buf ( n9150 , n9145 );
nand ( n9151 , n9149 , n9150 );
nand ( n9152 , n9148 , n9151 );
buf ( n9153 , n4745 );
not ( n9154 , n9153 );
and ( n9155 , n9152 , n9154 );
not ( n9156 , n9152 );
buf ( n9157 , n9153 );
and ( n9158 , n9156 , n9157 );
nor ( n9159 , n9155 , n9158 );
buf ( n9160 , n6556 );
buf ( n9161 , n4746 );
nand ( n9162 , n9160 , n9161 );
buf ( n9163 , n4747 );
buf ( n9164 , n9163 );
and ( n9165 , n9162 , n9164 );
not ( n9166 , n9162 );
not ( n9167 , n9163 );
and ( n9168 , n9166 , n9167 );
nor ( n9169 , n9165 , n9168 );
xor ( n9170 , n9159 , n9169 );
buf ( n9171 , n4748 );
nand ( n9172 , n7355 , n9171 );
buf ( n9173 , n4749 );
buf ( n9174 , n9173 );
and ( n9175 , n9172 , n9174 );
not ( n9176 , n9172 );
not ( n9177 , n9173 );
and ( n9178 , n9176 , n9177 );
nor ( n9179 , n9175 , n9178 );
xor ( n9180 , n9170 , n9179 );
buf ( n9181 , n9180 );
and ( n9182 , n9141 , n9181 );
not ( n9183 , n9141 );
not ( n9184 , n9181 );
and ( n9185 , n9183 , n9184 );
nor ( n9186 , n9182 , n9185 );
not ( n9187 , n9186 );
buf ( n9188 , n4750 );
nand ( n9189 , n8032 , n9188 );
buf ( n9190 , n4751 );
buf ( n9191 , n9190 );
and ( n9192 , n9189 , n9191 );
not ( n9193 , n9189 );
not ( n9194 , n9190 );
and ( n9195 , n9193 , n9194 );
nor ( n9196 , n9192 , n9195 );
not ( n9197 , n9196 );
buf ( n9198 , n4752 );
buf ( n9199 , n9198 );
not ( n9200 , n9199 );
buf ( n9201 , n4753 );
not ( n9202 , n9201 );
not ( n9203 , n9202 );
or ( n9204 , n9200 , n9203 );
not ( n9205 , n9198 );
buf ( n9206 , n9201 );
nand ( n9207 , n9205 , n9206 );
nand ( n9208 , n9204 , n9207 );
buf ( n9209 , n4754 );
buf ( n9210 , n9209 );
and ( n9211 , n9208 , n9210 );
not ( n9212 , n9208 );
not ( n9213 , n9209 );
and ( n9214 , n9212 , n9213 );
nor ( n9215 , n9211 , n9214 );
buf ( n9216 , n4755 );
nand ( n9217 , n6604 , n9216 );
buf ( n9218 , n4756 );
not ( n9219 , n9218 );
and ( n9220 , n9217 , n9219 );
not ( n9221 , n9217 );
buf ( n9222 , n9218 );
and ( n9223 , n9221 , n9222 );
nor ( n9224 , n9220 , n9223 );
xor ( n9225 , n9215 , n9224 );
buf ( n9226 , n4757 );
nand ( n9227 , n6647 , n9226 );
buf ( n9228 , n4758 );
not ( n9229 , n9228 );
and ( n9230 , n9227 , n9229 );
not ( n9231 , n9227 );
buf ( n9232 , n9228 );
and ( n9233 , n9231 , n9232 );
nor ( n9234 , n9230 , n9233 );
xnor ( n9235 , n9225 , n9234 );
not ( n9236 , n9235 );
not ( n9237 , n9236 );
or ( n9238 , n9197 , n9237 );
or ( n9239 , n9236 , n9196 );
nand ( n9240 , n9238 , n9239 );
not ( n9241 , n9240 );
not ( n9242 , n9241 );
buf ( n9243 , n4759 );
not ( n9244 , n9243 );
buf ( n9245 , n4760 );
buf ( n9246 , n9245 );
not ( n9247 , n9246 );
buf ( n9248 , n4761 );
not ( n9249 , n9248 );
not ( n9250 , n9249 );
or ( n9251 , n9247 , n9250 );
not ( n9252 , n9245 );
buf ( n9253 , n9248 );
nand ( n9254 , n9252 , n9253 );
nand ( n9255 , n9251 , n9254 );
xor ( n9256 , n9244 , n9255 );
not ( n9257 , n8051 );
buf ( n9258 , n4762 );
nand ( n9259 , n6577 , n9258 );
buf ( n9260 , n4763 );
buf ( n9261 , n9260 );
and ( n9262 , n9259 , n9261 );
not ( n9263 , n9259 );
not ( n9264 , n9260 );
and ( n9265 , n9263 , n9264 );
nor ( n9266 , n9262 , n9265 );
not ( n9267 , n9266 );
or ( n9268 , n9257 , n9267 );
or ( n9269 , n9266 , n8051 );
nand ( n9270 , n9268 , n9269 );
xnor ( n9271 , n9256 , n9270 );
buf ( n9272 , n9271 );
not ( n9273 , n9272 );
or ( n9274 , n9242 , n9273 );
buf ( n9275 , n9243 );
xor ( n9276 , n9275 , n9255 );
xnor ( n9277 , n9276 , n9270 );
nand ( n9278 , n9277 , n9240 );
nand ( n9279 , n9274 , n9278 );
buf ( n9280 , n4764 );
not ( n9281 , n9280 );
buf ( n9282 , n4765 );
buf ( n9283 , n9282 );
not ( n9284 , n9283 );
buf ( n9285 , n4766 );
not ( n9286 , n9285 );
not ( n9287 , n9286 );
or ( n9288 , n9284 , n9287 );
not ( n9289 , n9282 );
buf ( n9290 , n9285 );
nand ( n9291 , n9289 , n9290 );
nand ( n9292 , n9288 , n9291 );
buf ( n9293 , n4767 );
not ( n9294 , n9293 );
and ( n9295 , n9292 , n9294 );
not ( n9296 , n9292 );
buf ( n9297 , n9293 );
and ( n9298 , n9296 , n9297 );
nor ( n9299 , n9295 , n9298 );
buf ( n9300 , n4768 );
nand ( n9301 , n6927 , n9300 );
buf ( n9302 , n4769 );
buf ( n9303 , n9302 );
and ( n9304 , n9301 , n9303 );
not ( n9305 , n9301 );
not ( n9306 , n9302 );
and ( n9307 , n9305 , n9306 );
nor ( n9308 , n9304 , n9307 );
xor ( n9309 , n9299 , n9308 );
buf ( n9310 , n7013 );
buf ( n9311 , n4770 );
nand ( n9312 , n9310 , n9311 );
buf ( n9313 , n4771 );
not ( n9314 , n9313 );
and ( n9315 , n9312 , n9314 );
not ( n9316 , n9312 );
buf ( n9317 , n9313 );
and ( n9318 , n9316 , n9317 );
nor ( n9319 , n9315 , n9318 );
xnor ( n9320 , n9309 , n9319 );
not ( n9321 , n9320 );
not ( n9322 , n9321 );
not ( n9323 , n9322 );
or ( n9324 , n9281 , n9323 );
not ( n9325 , n9280 );
nand ( n9326 , n9325 , n9321 );
nand ( n9327 , n9324 , n9326 );
buf ( n9328 , n4772 );
nand ( n9329 , n8364 , n9328 );
buf ( n9330 , n4773 );
buf ( n9331 , n9330 );
and ( n9332 , n9329 , n9331 );
not ( n9333 , n9329 );
not ( n9334 , n9330 );
and ( n9335 , n9333 , n9334 );
nor ( n9336 , n9332 , n9335 );
not ( n9337 , n9336 );
buf ( n9338 , n4774 );
nand ( n9339 , n6770 , n9338 );
buf ( n9340 , n4775 );
not ( n9341 , n9340 );
and ( n9342 , n9339 , n9341 );
not ( n9343 , n9339 );
buf ( n9344 , n9340 );
and ( n9345 , n9343 , n9344 );
nor ( n9346 , n9342 , n9345 );
not ( n9347 , n9346 );
or ( n9348 , n9337 , n9347 );
or ( n9349 , n9336 , n9346 );
nand ( n9350 , n9348 , n9349 );
buf ( n9351 , n4776 );
buf ( n9352 , n9351 );
not ( n9353 , n9352 );
buf ( n9354 , n4777 );
not ( n9355 , n9354 );
not ( n9356 , n9355 );
or ( n9357 , n9353 , n9356 );
not ( n9358 , n9351 );
buf ( n9359 , n9354 );
nand ( n9360 , n9358 , n9359 );
nand ( n9361 , n9357 , n9360 );
buf ( n9362 , n4778 );
not ( n9363 , n9362 );
and ( n9364 , n9361 , n9363 );
not ( n9365 , n9361 );
buf ( n9366 , n9362 );
and ( n9367 , n9365 , n9366 );
nor ( n9368 , n9364 , n9367 );
not ( n9369 , n9368 );
and ( n9370 , n9350 , n9369 );
not ( n9371 , n9350 );
and ( n9372 , n9371 , n9368 );
nor ( n9373 , n9370 , n9372 );
not ( n9374 , n9373 );
and ( n9375 , n9327 , n9374 );
not ( n9376 , n9327 );
not ( n9377 , n9374 );
and ( n9378 , n9376 , n9377 );
nor ( n9379 , n9375 , n9378 );
nor ( n9380 , n9279 , n9379 );
not ( n9381 , n9380 );
or ( n9382 , n9187 , n9381 );
or ( n9383 , n9380 , n9186 );
nand ( n9384 , n9382 , n9383 );
not ( n9385 , n9384 );
nand ( n9386 , n9186 , n9279 );
not ( n9387 , n9386 );
buf ( n9388 , n4779 );
buf ( n9389 , n9388 );
not ( n9390 , n9389 );
buf ( n9391 , n4780 );
buf ( n9392 , n9391 );
not ( n9393 , n9392 );
buf ( n9394 , n4781 );
not ( n9395 , n9394 );
not ( n9396 , n9395 );
or ( n9397 , n9393 , n9396 );
not ( n9398 , n9391 );
buf ( n9399 , n9394 );
nand ( n9400 , n9398 , n9399 );
nand ( n9401 , n9397 , n9400 );
buf ( n9402 , n4782 );
not ( n9403 , n9402 );
and ( n9404 , n9401 , n9403 );
not ( n9405 , n9401 );
buf ( n9406 , n9402 );
and ( n9407 , n9405 , n9406 );
nor ( n9408 , n9404 , n9407 );
xor ( n9409 , n9408 , n8796 );
buf ( n9410 , n4783 );
nand ( n9411 , n6605 , n9410 );
buf ( n9412 , n4784 );
buf ( n9413 , n9412 );
and ( n9414 , n9411 , n9413 );
not ( n9415 , n9411 );
not ( n9416 , n9412 );
and ( n9417 , n9415 , n9416 );
nor ( n9418 , n9414 , n9417 );
xor ( n9419 , n9409 , n9418 );
not ( n9420 , n9419 );
or ( n9421 , n9390 , n9420 );
or ( n9422 , n9419 , n9389 );
nand ( n9423 , n9421 , n9422 );
buf ( n9424 , n4785 );
buf ( n9425 , n9424 );
not ( n9426 , n9425 );
buf ( n9427 , n4786 );
not ( n9428 , n9427 );
not ( n9429 , n9428 );
or ( n9430 , n9426 , n9429 );
not ( n9431 , n9424 );
buf ( n9432 , n9427 );
nand ( n9433 , n9431 , n9432 );
nand ( n9434 , n9430 , n9433 );
buf ( n9435 , n4787 );
not ( n9436 , n9435 );
and ( n9437 , n9434 , n9436 );
not ( n9438 , n9434 );
buf ( n9439 , n9435 );
and ( n9440 , n9438 , n9439 );
nor ( n9441 , n9437 , n9440 );
buf ( n9442 , n4788 );
nand ( n9443 , n8124 , n9442 );
buf ( n9444 , n4789 );
not ( n9445 , n9444 );
and ( n9446 , n9443 , n9445 );
not ( n9447 , n9443 );
buf ( n9448 , n9444 );
and ( n9449 , n9447 , n9448 );
nor ( n9450 , n9446 , n9449 );
xor ( n9451 , n9441 , n9450 );
buf ( n9452 , n4790 );
nand ( n9453 , n6816 , n9452 );
buf ( n9454 , n4791 );
not ( n9455 , n9454 );
and ( n9456 , n9453 , n9455 );
not ( n9457 , n9453 );
buf ( n9458 , n9454 );
and ( n9459 , n9457 , n9458 );
nor ( n9460 , n9456 , n9459 );
xnor ( n9461 , n9451 , n9460 );
buf ( n9462 , n9461 );
and ( n9463 , n9423 , n9462 );
not ( n9464 , n9423 );
not ( n9465 , n9462 );
and ( n9466 , n9464 , n9465 );
nor ( n9467 , n9463 , n9466 );
not ( n9468 , n9467 );
and ( n9469 , n9387 , n9468 );
buf ( n9470 , n9279 );
nand ( n9471 , n9186 , n9470 );
and ( n9472 , n9471 , n9467 );
nor ( n9473 , n9469 , n9472 );
not ( n9474 , n9473 );
buf ( n9475 , n4792 );
buf ( n9476 , n9475 );
not ( n9477 , n9476 );
buf ( n9478 , n4793 );
not ( n9479 , n9478 );
not ( n9480 , n9479 );
or ( n9481 , n9477 , n9480 );
not ( n9482 , n9475 );
buf ( n9483 , n9478 );
nand ( n9484 , n9482 , n9483 );
nand ( n9485 , n9481 , n9484 );
buf ( n9486 , n4794 );
buf ( n9487 , n9486 );
and ( n9488 , n9485 , n9487 );
not ( n9489 , n9485 );
not ( n9490 , n9486 );
and ( n9491 , n9489 , n9490 );
nor ( n9492 , n9488 , n9491 );
buf ( n9493 , n4795 );
nand ( n9494 , n7563 , n9493 );
buf ( n9495 , n4796 );
buf ( n9496 , n9495 );
and ( n9497 , n9494 , n9496 );
not ( n9498 , n9494 );
not ( n9499 , n9495 );
and ( n9500 , n9498 , n9499 );
nor ( n9501 , n9497 , n9500 );
xor ( n9502 , n9492 , n9501 );
buf ( n9503 , n4797 );
nand ( n9504 , n8223 , n9503 );
buf ( n9505 , n4798 );
not ( n9506 , n9505 );
and ( n9507 , n9504 , n9506 );
not ( n9508 , n9504 );
buf ( n9509 , n9505 );
and ( n9510 , n9508 , n9509 );
nor ( n9511 , n9507 , n9510 );
xnor ( n9512 , n9502 , n9511 );
not ( n9513 , n9512 );
not ( n9514 , n9513 );
buf ( n9515 , n4799 );
not ( n9516 , n9515 );
and ( n9517 , n9514 , n9516 );
buf ( n9518 , n9512 );
not ( n9519 , n9518 );
and ( n9520 , n9519 , n9515 );
nor ( n9521 , n9517 , n9520 );
buf ( n9522 , n4800 );
buf ( n9523 , n9522 );
not ( n9524 , n9523 );
buf ( n9525 , n4801 );
not ( n9526 , n9525 );
not ( n9527 , n9526 );
or ( n9528 , n9524 , n9527 );
not ( n9529 , n9522 );
buf ( n9530 , n9525 );
nand ( n9531 , n9529 , n9530 );
nand ( n9532 , n9528 , n9531 );
buf ( n9533 , n4802 );
not ( n9534 , n9533 );
and ( n9535 , n9532 , n9534 );
not ( n9536 , n9532 );
buf ( n9537 , n9533 );
and ( n9538 , n9536 , n9537 );
nor ( n9539 , n9535 , n9538 );
not ( n9540 , n9539 );
buf ( n9541 , n4803 );
nand ( n9542 , n6604 , n9541 );
buf ( n9543 , n4804 );
xor ( n9544 , n9542 , n9543 );
xor ( n9545 , n9540 , n9544 );
buf ( n9546 , n4805 );
nand ( n9547 , n7569 , n9546 );
buf ( n9548 , n4806 );
buf ( n9549 , n9548 );
and ( n9550 , n9547 , n9549 );
not ( n9551 , n9547 );
not ( n9552 , n9548 );
and ( n9553 , n9551 , n9552 );
nor ( n9554 , n9550 , n9553 );
xnor ( n9555 , n9545 , n9554 );
not ( n9556 , n9555 );
not ( n9557 , n9556 );
and ( n9558 , n9521 , n9557 );
not ( n9559 , n9521 );
xor ( n9560 , n9539 , n9544 );
xnor ( n9561 , n9560 , n9554 );
buf ( n9562 , n9561 );
and ( n9563 , n9559 , n9562 );
nor ( n9564 , n9558 , n9563 );
not ( n9565 , n9564 );
buf ( n9566 , n4807 );
nand ( n9567 , n7868 , n9566 );
buf ( n9568 , n4808 );
not ( n9569 , n9568 );
and ( n9570 , n9567 , n9569 );
not ( n9571 , n9567 );
buf ( n9572 , n9568 );
and ( n9573 , n9571 , n9572 );
nor ( n9574 , n9570 , n9573 );
buf ( n9575 , n9574 );
not ( n9576 , n9575 );
buf ( n9577 , n4809 );
buf ( n9578 , n4810 );
buf ( n9579 , n9578 );
not ( n9580 , n9579 );
buf ( n9581 , n4811 );
not ( n9582 , n9581 );
not ( n9583 , n9582 );
or ( n9584 , n9580 , n9583 );
not ( n9585 , n9578 );
buf ( n9586 , n9581 );
nand ( n9587 , n9585 , n9586 );
nand ( n9588 , n9584 , n9587 );
xor ( n9589 , n9577 , n9588 );
buf ( n9590 , n4812 );
buf ( n9591 , n4813 );
not ( n9592 , n9591 );
xor ( n9593 , n9590 , n9592 );
buf ( n9594 , n4814 );
nand ( n9595 , n8323 , n9594 );
xnor ( n9596 , n9593 , n9595 );
xnor ( n9597 , n9589 , n9596 );
not ( n9598 , n9597 );
not ( n9599 , n9598 );
or ( n9600 , n9576 , n9599 );
not ( n9601 , n9575 );
nand ( n9602 , n9601 , n9597 );
nand ( n9603 , n9600 , n9602 );
buf ( n9604 , n4815 );
buf ( n9605 , n9604 );
not ( n9606 , n9605 );
buf ( n9607 , n4816 );
not ( n9608 , n9607 );
not ( n9609 , n9608 );
or ( n9610 , n9606 , n9609 );
not ( n9611 , n9604 );
buf ( n9612 , n9607 );
nand ( n9613 , n9611 , n9612 );
nand ( n9614 , n9610 , n9613 );
buf ( n9615 , n4817 );
buf ( n9616 , n9615 );
and ( n9617 , n9614 , n9616 );
not ( n9618 , n9614 );
not ( n9619 , n9615 );
and ( n9620 , n9618 , n9619 );
nor ( n9621 , n9617 , n9620 );
buf ( n9622 , n4818 );
nand ( n9623 , n8781 , n9622 );
buf ( n9624 , n4819 );
buf ( n9625 , n9624 );
and ( n9626 , n9623 , n9625 );
not ( n9627 , n9623 );
not ( n9628 , n9624 );
and ( n9629 , n9627 , n9628 );
nor ( n9630 , n9626 , n9629 );
xor ( n9631 , n9621 , n9630 );
buf ( n9632 , n4820 );
nand ( n9633 , n6828 , n9632 );
buf ( n9634 , n4821 );
buf ( n9635 , n9634 );
and ( n9636 , n9633 , n9635 );
not ( n9637 , n9633 );
not ( n9638 , n9634 );
and ( n9639 , n9637 , n9638 );
nor ( n9640 , n9636 , n9639 );
not ( n9641 , n9640 );
xnor ( n9642 , n9631 , n9641 );
not ( n9643 , n9642 );
not ( n9644 , n9643 );
and ( n9645 , n9603 , n9644 );
not ( n9646 , n9603 );
xor ( n9647 , n9621 , n9640 );
not ( n9648 , n9630 );
xor ( n9649 , n9647 , n9648 );
buf ( n9650 , n9649 );
and ( n9651 , n9646 , n9650 );
nor ( n9652 , n9645 , n9651 );
nand ( n9653 , n9565 , n9652 );
buf ( n9654 , n4822 );
buf ( n9655 , n9654 );
not ( n9656 , n9655 );
buf ( n9657 , n4823 );
buf ( n9658 , n9657 );
not ( n9659 , n9658 );
buf ( n9660 , n4824 );
not ( n9661 , n9660 );
not ( n9662 , n9661 );
or ( n9663 , n9659 , n9662 );
not ( n9664 , n9657 );
buf ( n9665 , n9660 );
nand ( n9666 , n9664 , n9665 );
nand ( n9667 , n9663 , n9666 );
buf ( n9668 , n4825 );
buf ( n9669 , n9668 );
and ( n9670 , n9667 , n9669 );
not ( n9671 , n9667 );
not ( n9672 , n9668 );
and ( n9673 , n9671 , n9672 );
nor ( n9674 , n9670 , n9673 );
buf ( n9675 , n4826 );
nand ( n9676 , n8124 , n9675 );
buf ( n9677 , n4827 );
buf ( n9678 , n9677 );
and ( n9679 , n9676 , n9678 );
not ( n9680 , n9676 );
not ( n9681 , n9677 );
and ( n9682 , n9680 , n9681 );
nor ( n9683 , n9679 , n9682 );
xor ( n9684 , n9674 , n9683 );
buf ( n9685 , n4828 );
nand ( n9686 , n8375 , n9685 );
buf ( n9687 , n4829 );
not ( n9688 , n9687 );
and ( n9689 , n9686 , n9688 );
not ( n9690 , n9686 );
buf ( n9691 , n9687 );
and ( n9692 , n9690 , n9691 );
nor ( n9693 , n9689 , n9692 );
xnor ( n9694 , n9684 , n9693 );
not ( n9695 , n9694 );
not ( n9696 , n9695 );
or ( n9697 , n9656 , n9696 );
not ( n9698 , n9655 );
nand ( n9699 , n9698 , n9694 );
nand ( n9700 , n9697 , n9699 );
not ( n9701 , n9700 );
buf ( n9702 , n4830 );
buf ( n9703 , n9702 );
not ( n9704 , n9703 );
buf ( n9705 , n4831 );
not ( n9706 , n9705 );
not ( n9707 , n9706 );
or ( n9708 , n9704 , n9707 );
not ( n9709 , n9702 );
buf ( n9710 , n9705 );
nand ( n9711 , n9709 , n9710 );
nand ( n9712 , n9708 , n9711 );
not ( n9713 , n9712 );
xor ( n9714 , n6476 , n9713 );
buf ( n9715 , n4832 );
not ( n9716 , n9715 );
buf ( n9717 , n4833 );
nand ( n9718 , n8966 , n9717 );
buf ( n9719 , n4834 );
buf ( n9720 , n9719 );
and ( n9721 , n9718 , n9720 );
not ( n9722 , n9718 );
not ( n9723 , n9719 );
and ( n9724 , n9722 , n9723 );
nor ( n9725 , n9721 , n9724 );
not ( n9726 , n9725 );
or ( n9727 , n9716 , n9726 );
or ( n9728 , n9725 , n9715 );
nand ( n9729 , n9727 , n9728 );
xnor ( n9730 , n9714 , n9729 );
buf ( n9731 , n9730 );
not ( n9732 , n9731 );
and ( n9733 , n9701 , n9732 );
and ( n9734 , n9731 , n9700 );
nor ( n9735 , n9733 , n9734 );
and ( n9736 , n9653 , n9735 );
not ( n9737 , n9653 );
not ( n9738 , n9735 );
and ( n9739 , n9737 , n9738 );
nor ( n9740 , n9736 , n9739 );
not ( n9741 , n9740 );
or ( n9742 , n9474 , n9741 );
or ( n9743 , n9740 , n9473 );
nand ( n9744 , n9742 , n9743 );
buf ( n9745 , n4835 );
buf ( n9746 , n9745 );
not ( n9747 , n9746 );
buf ( n9748 , n4836 );
buf ( n9749 , n9748 );
not ( n9750 , n9749 );
buf ( n9751 , n4837 );
not ( n9752 , n9751 );
not ( n9753 , n9752 );
or ( n9754 , n9750 , n9753 );
not ( n9755 , n9748 );
buf ( n9756 , n9751 );
nand ( n9757 , n9755 , n9756 );
nand ( n9758 , n9754 , n9757 );
buf ( n9759 , n4838 );
not ( n9760 , n9759 );
and ( n9761 , n9758 , n9760 );
not ( n9762 , n9758 );
buf ( n9763 , n9759 );
and ( n9764 , n9762 , n9763 );
nor ( n9765 , n9761 , n9764 );
buf ( n9766 , n4839 );
nand ( n9767 , n6927 , n9766 );
buf ( n9768 , n4840 );
buf ( n9769 , n9768 );
and ( n9770 , n9767 , n9769 );
not ( n9771 , n9767 );
not ( n9772 , n9768 );
and ( n9773 , n9771 , n9772 );
nor ( n9774 , n9770 , n9773 );
xor ( n9775 , n9765 , n9774 );
buf ( n9776 , n4841 );
nand ( n9777 , n9310 , n9776 );
buf ( n9778 , n4842 );
not ( n9779 , n9778 );
and ( n9780 , n9777 , n9779 );
not ( n9781 , n9777 );
buf ( n9782 , n9778 );
and ( n9783 , n9781 , n9782 );
nor ( n9784 , n9780 , n9783 );
xnor ( n9785 , n9775 , n9784 );
not ( n9786 , n9785 );
or ( n9787 , n9747 , n9786 );
buf ( n9788 , n9785 );
or ( n9789 , n9788 , n9746 );
nand ( n9790 , n9787 , n9789 );
not ( n9791 , n9790 );
not ( n9792 , n9791 );
buf ( n9793 , n4843 );
not ( n9794 , n9793 );
buf ( n9795 , n4844 );
buf ( n9796 , n9795 );
and ( n9797 , n9794 , n9796 );
not ( n9798 , n9794 );
not ( n9799 , n9795 );
and ( n9800 , n9798 , n9799 );
nor ( n9801 , n9797 , n9800 );
buf ( n9802 , n4845 );
nand ( n9803 , n9160 , n9802 );
buf ( n9804 , n4846 );
buf ( n9805 , n9804 );
and ( n9806 , n9803 , n9805 );
not ( n9807 , n9803 );
not ( n9808 , n9804 );
and ( n9809 , n9807 , n9808 );
nor ( n9810 , n9806 , n9809 );
not ( n9811 , n9810 );
buf ( n9812 , n8322 );
buf ( n9813 , n4847 );
nand ( n9814 , n9812 , n9813 );
buf ( n9815 , n4848 );
not ( n9816 , n9815 );
and ( n9817 , n9814 , n9816 );
not ( n9818 , n9814 );
buf ( n9819 , n9815 );
and ( n9820 , n9818 , n9819 );
nor ( n9821 , n9817 , n9820 );
not ( n9822 , n9821 );
or ( n9823 , n9811 , n9822 );
not ( n9824 , n9821 );
not ( n9825 , n9810 );
nand ( n9826 , n9824 , n9825 );
nand ( n9827 , n9823 , n9826 );
buf ( n9828 , n4849 );
not ( n9829 , n9828 );
and ( n9830 , n9827 , n9829 );
not ( n9831 , n9827 );
buf ( n9832 , n9828 );
and ( n9833 , n9831 , n9832 );
nor ( n9834 , n9830 , n9833 );
not ( n9835 , n9834 );
and ( n9836 , n9801 , n9835 );
not ( n9837 , n9801 );
and ( n9838 , n9837 , n9834 );
nor ( n9839 , n9836 , n9838 );
not ( n9840 , n9839 );
not ( n9841 , n9840 );
or ( n9842 , n9792 , n9841 );
xor ( n9843 , n9829 , n9801 );
xnor ( n9844 , n9843 , n9827 );
nand ( n9845 , n9844 , n9790 );
nand ( n9846 , n9842 , n9845 );
not ( n9847 , n9846 );
buf ( n9848 , n4850 );
nand ( n9849 , n8124 , n9848 );
buf ( n9850 , n4851 );
xor ( n9851 , n9849 , n9850 );
not ( n9852 , n9851 );
buf ( n9853 , n4852 );
nand ( n9854 , n7606 , n9853 );
buf ( n9855 , n4853 );
buf ( n9856 , n9855 );
and ( n9857 , n9854 , n9856 );
not ( n9858 , n9854 );
not ( n9859 , n9855 );
and ( n9860 , n9858 , n9859 );
nor ( n9861 , n9857 , n9860 );
not ( n9862 , n9861 );
buf ( n9863 , n4854 );
nand ( n9864 , n7344 , n9863 );
buf ( n9865 , n4855 );
not ( n9866 , n9865 );
and ( n9867 , n9864 , n9866 );
not ( n9868 , n9864 );
buf ( n9869 , n9865 );
and ( n9870 , n9868 , n9869 );
nor ( n9871 , n9867 , n9870 );
not ( n9872 , n9871 );
or ( n9873 , n9862 , n9872 );
or ( n9874 , n9861 , n9871 );
nand ( n9875 , n9873 , n9874 );
buf ( n9876 , n4856 );
buf ( n9877 , n9876 );
not ( n9878 , n9877 );
buf ( n9879 , n4857 );
not ( n9880 , n9879 );
not ( n9881 , n9880 );
or ( n9882 , n9878 , n9881 );
not ( n9883 , n9876 );
buf ( n9884 , n9879 );
nand ( n9885 , n9883 , n9884 );
nand ( n9886 , n9882 , n9885 );
buf ( n9887 , n4858 );
not ( n9888 , n9887 );
and ( n9889 , n9886 , n9888 );
not ( n9890 , n9886 );
buf ( n9891 , n9887 );
and ( n9892 , n9890 , n9891 );
nor ( n9893 , n9889 , n9892 );
not ( n9894 , n9893 );
and ( n9895 , n9875 , n9894 );
not ( n9896 , n9875 );
and ( n9897 , n9896 , n9893 );
nor ( n9898 , n9895 , n9897 );
not ( n9899 , n9898 );
or ( n9900 , n9852 , n9899 );
or ( n9901 , n9898 , n9851 );
nand ( n9902 , n9900 , n9901 );
buf ( n9903 , n4859 );
buf ( n9904 , n9903 );
not ( n9905 , n9904 );
buf ( n9906 , n4860 );
not ( n9907 , n9906 );
not ( n9908 , n9907 );
or ( n9909 , n9905 , n9908 );
not ( n9910 , n9903 );
buf ( n9911 , n9906 );
nand ( n9912 , n9910 , n9911 );
nand ( n9913 , n9909 , n9912 );
buf ( n9914 , n4861 );
buf ( n9915 , n9914 );
and ( n9916 , n9913 , n9915 );
not ( n9917 , n9913 );
not ( n9918 , n9914 );
and ( n9919 , n9917 , n9918 );
nor ( n9920 , n9916 , n9919 );
buf ( n9921 , n4862 );
nand ( n9922 , n7787 , n9921 );
buf ( n9923 , n4863 );
buf ( n9924 , n9923 );
and ( n9925 , n9922 , n9924 );
not ( n9926 , n9922 );
not ( n9927 , n9923 );
and ( n9928 , n9926 , n9927 );
nor ( n9929 , n9925 , n9928 );
xor ( n9930 , n9920 , n9929 );
buf ( n9931 , n4864 );
nand ( n9932 , n7247 , n9931 );
buf ( n9933 , n4865 );
buf ( n9934 , n9933 );
and ( n9935 , n9932 , n9934 );
not ( n9936 , n9932 );
not ( n9937 , n9933 );
and ( n9938 , n9936 , n9937 );
nor ( n9939 , n9935 , n9938 );
xnor ( n9940 , n9930 , n9939 );
not ( n9941 , n9940 );
not ( n9942 , n9941 );
and ( n9943 , n9902 , n9942 );
not ( n9944 , n9902 );
and ( n9945 , n9944 , n9941 );
nor ( n9946 , n9943 , n9945 );
not ( n9947 , n9946 );
nand ( n9948 , n9847 , n9947 );
buf ( n9949 , n4866 );
buf ( n9950 , n9949 );
buf ( n9951 , n4867 );
buf ( n9952 , n9951 );
not ( n9953 , n9952 );
buf ( n9954 , n4868 );
not ( n9955 , n9954 );
not ( n9956 , n9955 );
or ( n9957 , n9953 , n9956 );
not ( n9958 , n9951 );
buf ( n9959 , n9954 );
nand ( n9960 , n9958 , n9959 );
nand ( n9961 , n9957 , n9960 );
buf ( n9962 , n4869 );
buf ( n9963 , n9962 );
and ( n9964 , n9961 , n9963 );
not ( n9965 , n9961 );
not ( n9966 , n9962 );
and ( n9967 , n9965 , n9966 );
nor ( n9968 , n9964 , n9967 );
not ( n9969 , n9968 );
buf ( n9970 , n4870 );
nand ( n9971 , n7698 , n9970 );
buf ( n9972 , n4871 );
buf ( n9973 , n9972 );
and ( n9974 , n9971 , n9973 );
not ( n9975 , n9971 );
not ( n9976 , n9972 );
and ( n9977 , n9975 , n9976 );
nor ( n9978 , n9974 , n9977 );
xor ( n9979 , n9969 , n9978 );
buf ( n9980 , n4872 );
nand ( n9981 , n7569 , n9980 );
buf ( n9982 , n4873 );
buf ( n9983 , n9982 );
and ( n9984 , n9981 , n9983 );
not ( n9985 , n9981 );
not ( n9986 , n9982 );
and ( n9987 , n9985 , n9986 );
nor ( n9988 , n9984 , n9987 );
xnor ( n9989 , n9979 , n9988 );
buf ( n9990 , n9989 );
xor ( n9991 , n9950 , n9990 );
buf ( n9992 , n4874 );
not ( n9993 , n9992 );
buf ( n9994 , n4875 );
not ( n9995 , n9994 );
buf ( n9996 , n4876 );
buf ( n9997 , n9996 );
and ( n9998 , n9995 , n9997 );
not ( n9999 , n9995 );
not ( n10000 , n9996 );
and ( n10001 , n9999 , n10000 );
nor ( n10002 , n9998 , n10001 );
xor ( n10003 , n9993 , n10002 );
buf ( n10004 , n4877 );
buf ( n10005 , n4878 );
xor ( n10006 , n10004 , n10005 );
buf ( n10007 , n4879 );
nand ( n10008 , n6558 , n10007 );
xnor ( n10009 , n10006 , n10008 );
xnor ( n10010 , n10003 , n10009 );
buf ( n10011 , n10010 );
xnor ( n10012 , n9991 , n10011 );
not ( n10013 , n10012 );
and ( n10014 , n9948 , n10013 );
not ( n10015 , n9948 );
and ( n10016 , n10015 , n10012 );
nor ( n10017 , n10014 , n10016 );
not ( n10018 , n10017 );
and ( n10019 , n9744 , n10018 );
not ( n10020 , n9744 );
and ( n10021 , n10020 , n10017 );
nor ( n10022 , n10019 , n10021 );
not ( n10023 , n10022 );
buf ( n10024 , n4880 );
buf ( n10025 , n10024 );
not ( n10026 , n10025 );
not ( n10027 , n8963 );
not ( n10028 , n8975 );
or ( n10029 , n10027 , n10028 );
or ( n10030 , n8963 , n8975 );
nand ( n10031 , n10029 , n10030 );
not ( n10032 , n8953 );
and ( n10033 , n10031 , n10032 );
not ( n10034 , n10031 );
and ( n10035 , n10034 , n8953 );
nor ( n10036 , n10033 , n10035 );
buf ( n10037 , n10036 );
not ( n10038 , n10037 );
or ( n10039 , n10026 , n10038 );
not ( n10040 , n10025 );
nand ( n10041 , n10040 , n8978 );
nand ( n10042 , n10039 , n10041 );
and ( n10043 , n10042 , n8986 );
not ( n10044 , n10042 );
and ( n10045 , n10044 , n7540 );
nor ( n10046 , n10043 , n10045 );
not ( n10047 , n10046 );
buf ( n10048 , n4881 );
buf ( n10049 , n10048 );
not ( n10050 , n10049 );
buf ( n10051 , n4882 );
buf ( n10052 , n10051 );
not ( n10053 , n10052 );
buf ( n10054 , n4883 );
not ( n10055 , n10054 );
not ( n10056 , n10055 );
or ( n10057 , n10053 , n10056 );
not ( n10058 , n10051 );
buf ( n10059 , n10054 );
nand ( n10060 , n10058 , n10059 );
nand ( n10061 , n10057 , n10060 );
buf ( n10062 , n4884 );
buf ( n10063 , n10062 );
and ( n10064 , n10061 , n10063 );
not ( n10065 , n10061 );
not ( n10066 , n10062 );
and ( n10067 , n10065 , n10066 );
nor ( n10068 , n10064 , n10067 );
buf ( n10069 , n4885 );
nand ( n10070 , n6502 , n10069 );
buf ( n10071 , n4886 );
buf ( n10072 , n10071 );
and ( n10073 , n10070 , n10072 );
not ( n10074 , n10070 );
not ( n10075 , n10071 );
and ( n10076 , n10074 , n10075 );
nor ( n10077 , n10073 , n10076 );
xor ( n10078 , n10068 , n10077 );
buf ( n10079 , n4887 );
nand ( n10080 , n8125 , n10079 );
buf ( n10081 , n4888 );
not ( n10082 , n10081 );
and ( n10083 , n10080 , n10082 );
not ( n10084 , n10080 );
buf ( n10085 , n10081 );
and ( n10086 , n10084 , n10085 );
nor ( n10087 , n10083 , n10086 );
xnor ( n10088 , n10078 , n10087 );
buf ( n10089 , n10088 );
not ( n10090 , n10089 );
not ( n10091 , n10090 );
or ( n10092 , n10050 , n10091 );
not ( n10093 , n10048 );
nand ( n10094 , n10089 , n10093 );
nand ( n10095 , n10092 , n10094 );
buf ( n10096 , n4889 );
buf ( n10097 , n10096 );
buf ( n10098 , n4890 );
buf ( n10099 , n10098 );
not ( n10100 , n10099 );
buf ( n10101 , n4891 );
not ( n10102 , n10101 );
not ( n10103 , n10102 );
or ( n10104 , n10100 , n10103 );
not ( n10105 , n10098 );
buf ( n10106 , n10101 );
nand ( n10107 , n10105 , n10106 );
nand ( n10108 , n10104 , n10107 );
xor ( n10109 , n10097 , n10108 );
buf ( n10110 , n4892 );
not ( n10111 , n10110 );
buf ( n10112 , n4893 );
nand ( n10113 , n7355 , n10112 );
buf ( n10114 , n4894 );
buf ( n10115 , n10114 );
and ( n10116 , n10113 , n10115 );
not ( n10117 , n10113 );
not ( n10118 , n10114 );
and ( n10119 , n10117 , n10118 );
nor ( n10120 , n10116 , n10119 );
not ( n10121 , n10120 );
or ( n10122 , n10111 , n10121 );
or ( n10123 , n10120 , n10110 );
nand ( n10124 , n10122 , n10123 );
xnor ( n10125 , n10109 , n10124 );
buf ( n10126 , n10125 );
buf ( n10127 , n10126 );
xnor ( n10128 , n10095 , n10127 );
not ( n10129 , n10128 );
buf ( n10130 , n9064 );
not ( n10131 , n10130 );
not ( n10132 , n9061 );
and ( n10133 , n10131 , n10132 );
and ( n10134 , n10130 , n9061 );
nor ( n10135 , n10133 , n10134 );
not ( n10136 , n10135 );
buf ( n10137 , n4895 );
buf ( n10138 , n10137 );
not ( n10139 , n10138 );
buf ( n10140 , n4896 );
not ( n10141 , n10140 );
not ( n10142 , n10141 );
or ( n10143 , n10139 , n10142 );
not ( n10144 , n10137 );
buf ( n10145 , n10140 );
nand ( n10146 , n10144 , n10145 );
nand ( n10147 , n10143 , n10146 );
buf ( n10148 , n4897 );
buf ( n10149 , n10148 );
and ( n10150 , n10147 , n10149 );
not ( n10151 , n10147 );
not ( n10152 , n10148 );
and ( n10153 , n10151 , n10152 );
nor ( n10154 , n10150 , n10153 );
buf ( n10155 , n4898 );
nand ( n10156 , n6828 , n10155 );
buf ( n10157 , n4899 );
buf ( n10158 , n10157 );
and ( n10159 , n10156 , n10158 );
not ( n10160 , n10156 );
not ( n10161 , n10157 );
and ( n10162 , n10160 , n10161 );
nor ( n10163 , n10159 , n10162 );
xor ( n10164 , n10154 , n10163 );
buf ( n10165 , n7013 );
buf ( n10166 , n4900 );
nand ( n10167 , n10165 , n10166 );
buf ( n10168 , n4901 );
buf ( n10169 , n10168 );
and ( n10170 , n10167 , n10169 );
not ( n10171 , n10167 );
not ( n10172 , n10168 );
and ( n10173 , n10171 , n10172 );
nor ( n10174 , n10170 , n10173 );
xor ( n10175 , n10164 , n10174 );
not ( n10176 , n10175 );
or ( n10177 , n10136 , n10176 );
or ( n10178 , n10175 , n10135 );
nand ( n10179 , n10177 , n10178 );
not ( n10180 , n10179 );
buf ( n10181 , n4902 );
nand ( n10182 , n6916 , n10181 );
buf ( n10183 , n4903 );
buf ( n10184 , n10183 );
and ( n10185 , n10182 , n10184 );
not ( n10186 , n10182 );
not ( n10187 , n10183 );
and ( n10188 , n10186 , n10187 );
nor ( n10189 , n10185 , n10188 );
not ( n10190 , n10189 );
buf ( n10191 , n4904 );
nand ( n10192 , n8966 , n10191 );
buf ( n10193 , n4905 );
not ( n10194 , n10193 );
and ( n10195 , n10192 , n10194 );
not ( n10196 , n10192 );
buf ( n10197 , n10193 );
and ( n10198 , n10196 , n10197 );
nor ( n10199 , n10195 , n10198 );
not ( n10200 , n10199 );
or ( n10201 , n10190 , n10200 );
or ( n10202 , n10189 , n10199 );
nand ( n10203 , n10201 , n10202 );
buf ( n10204 , n4906 );
buf ( n10205 , n10204 );
not ( n10206 , n10205 );
buf ( n10207 , n4907 );
not ( n10208 , n10207 );
not ( n10209 , n10208 );
or ( n10210 , n10206 , n10209 );
not ( n10211 , n10204 );
buf ( n10212 , n10207 );
nand ( n10213 , n10211 , n10212 );
nand ( n10214 , n10210 , n10213 );
buf ( n10215 , n4908 );
buf ( n10216 , n10215 );
and ( n10217 , n10214 , n10216 );
not ( n10218 , n10214 );
not ( n10219 , n10215 );
and ( n10220 , n10218 , n10219 );
nor ( n10221 , n10217 , n10220 );
not ( n10222 , n10221 );
and ( n10223 , n10203 , n10222 );
not ( n10224 , n10203 );
and ( n10225 , n10224 , n10221 );
nor ( n10226 , n10223 , n10225 );
buf ( n10227 , n10226 );
buf ( n10228 , n10227 );
not ( n10229 , n10228 );
and ( n10230 , n10180 , n10229 );
and ( n10231 , n10179 , n10227 );
nor ( n10232 , n10230 , n10231 );
not ( n10233 , n10232 );
nand ( n10234 , n10129 , n10233 );
not ( n10235 , n10234 );
or ( n10236 , n10047 , n10235 );
or ( n10237 , n10046 , n10234 );
nand ( n10238 , n10236 , n10237 );
not ( n10239 , n7896 );
buf ( n10240 , n4909 );
buf ( n10241 , n10240 );
not ( n10242 , n10241 );
buf ( n10243 , n4910 );
not ( n10244 , n10243 );
not ( n10245 , n10244 );
or ( n10246 , n10242 , n10245 );
not ( n10247 , n10240 );
buf ( n10248 , n10243 );
nand ( n10249 , n10247 , n10248 );
nand ( n10250 , n10246 , n10249 );
not ( n10251 , n10250 );
buf ( n10252 , n4911 );
buf ( n10253 , n4912 );
xor ( n10254 , n10252 , n10253 );
buf ( n10255 , n4913 );
nand ( n10256 , n6577 , n10255 );
buf ( n10257 , n4914 );
not ( n10258 , n10257 );
and ( n10259 , n10256 , n10258 );
not ( n10260 , n10256 );
buf ( n10261 , n10257 );
and ( n10262 , n10260 , n10261 );
nor ( n10263 , n10259 , n10262 );
xnor ( n10264 , n10254 , n10263 );
not ( n10265 , n10264 );
or ( n10266 , n10251 , n10265 );
not ( n10267 , n10264 );
not ( n10268 , n10250 );
nand ( n10269 , n10267 , n10268 );
nand ( n10270 , n10266 , n10269 );
buf ( n10271 , n10270 );
not ( n10272 , n10271 );
or ( n10273 , n10239 , n10272 );
or ( n10274 , n10271 , n7896 );
nand ( n10275 , n10273 , n10274 );
buf ( n10276 , n4915 );
buf ( n10277 , n4916 );
nand ( n10278 , n8537 , n10277 );
buf ( n10279 , n4917 );
buf ( n10280 , n10279 );
and ( n10281 , n10278 , n10280 );
not ( n10282 , n10278 );
not ( n10283 , n10279 );
and ( n10284 , n10282 , n10283 );
nor ( n10285 , n10281 , n10284 );
xor ( n10286 , n10276 , n10285 );
buf ( n10287 , n4918 );
nand ( n10288 , n9310 , n10287 );
buf ( n10289 , n4919 );
not ( n10290 , n10289 );
and ( n10291 , n10288 , n10290 );
not ( n10292 , n10288 );
buf ( n10293 , n10289 );
and ( n10294 , n10292 , n10293 );
nor ( n10295 , n10291 , n10294 );
xnor ( n10296 , n10286 , n10295 );
not ( n10297 , n10296 );
buf ( n10298 , n4920 );
not ( n10299 , n10298 );
buf ( n10300 , n4921 );
buf ( n10301 , n10300 );
and ( n10302 , n10299 , n10301 );
not ( n10303 , n10299 );
not ( n10304 , n10300 );
and ( n10305 , n10303 , n10304 );
nor ( n10306 , n10302 , n10305 );
not ( n10307 , n10306 );
and ( n10308 , n10297 , n10307 );
and ( n10309 , n10296 , n10306 );
nor ( n10310 , n10308 , n10309 );
buf ( n10311 , n10310 );
and ( n10312 , n10275 , n10311 );
not ( n10313 , n10275 );
not ( n10314 , n10311 );
and ( n10315 , n10313 , n10314 );
nor ( n10316 , n10312 , n10315 );
buf ( n10317 , n4922 );
buf ( n10318 , n4923 );
nand ( n10319 , n9160 , n10318 );
buf ( n10320 , n4924 );
buf ( n10321 , n10320 );
and ( n10322 , n10319 , n10321 );
not ( n10323 , n10319 );
not ( n10324 , n10320 );
and ( n10325 , n10323 , n10324 );
nor ( n10326 , n10322 , n10325 );
xor ( n10327 , n10317 , n10326 );
buf ( n10328 , n4925 );
nand ( n10329 , n6605 , n10328 );
buf ( n10330 , n4926 );
not ( n10331 , n10330 );
and ( n10332 , n10329 , n10331 );
not ( n10333 , n10329 );
buf ( n10334 , n10330 );
and ( n10335 , n10333 , n10334 );
nor ( n10336 , n10332 , n10335 );
xnor ( n10337 , n10327 , n10336 );
not ( n10338 , n10337 );
buf ( n10339 , n4927 );
not ( n10340 , n10339 );
not ( n10341 , n10340 );
buf ( n10342 , n4928 );
not ( n10343 , n10342 );
and ( n10344 , n10341 , n10343 );
and ( n10345 , n10342 , n10340 );
nor ( n10346 , n10344 , n10345 );
not ( n10347 , n10346 );
and ( n10348 , n10338 , n10347 );
and ( n10349 , n10337 , n10346 );
nor ( n10350 , n10348 , n10349 );
buf ( n10351 , n10350 );
not ( n10352 , n10351 );
not ( n10353 , n9648 );
buf ( n10354 , n4929 );
buf ( n10355 , n10354 );
not ( n10356 , n10355 );
buf ( n10357 , n4930 );
not ( n10358 , n10357 );
not ( n10359 , n10358 );
or ( n10360 , n10356 , n10359 );
not ( n10361 , n10354 );
buf ( n10362 , n10357 );
nand ( n10363 , n10361 , n10362 );
nand ( n10364 , n10360 , n10363 );
buf ( n10365 , n4931 );
not ( n10366 , n10365 );
and ( n10367 , n10364 , n10366 );
not ( n10368 , n10364 );
buf ( n10369 , n10365 );
and ( n10370 , n10368 , n10369 );
nor ( n10371 , n10367 , n10370 );
buf ( n10372 , n6718 );
buf ( n10373 , n4932 );
nand ( n10374 , n10372 , n10373 );
buf ( n10375 , n4933 );
buf ( n10376 , n10375 );
and ( n10377 , n10374 , n10376 );
not ( n10378 , n10374 );
not ( n10379 , n10375 );
and ( n10380 , n10378 , n10379 );
nor ( n10381 , n10377 , n10380 );
xor ( n10382 , n10371 , n10381 );
buf ( n10383 , n6927 );
buf ( n10384 , n4934 );
nand ( n10385 , n10383 , n10384 );
buf ( n10386 , n4935 );
buf ( n10387 , n10386 );
and ( n10388 , n10385 , n10387 );
not ( n10389 , n10385 );
not ( n10390 , n10386 );
and ( n10391 , n10389 , n10390 );
nor ( n10392 , n10388 , n10391 );
xnor ( n10393 , n10382 , n10392 );
not ( n10394 , n10393 );
not ( n10395 , n10394 );
or ( n10396 , n10353 , n10395 );
not ( n10397 , n9648 );
buf ( n10398 , n10393 );
nand ( n10399 , n10397 , n10398 );
nand ( n10400 , n10396 , n10399 );
not ( n10401 , n10400 );
and ( n10402 , n10352 , n10401 );
and ( n10403 , n10351 , n10400 );
nor ( n10404 , n10402 , n10403 );
not ( n10405 , n10404 );
nand ( n10406 , n10316 , n10405 );
not ( n10407 , n10406 );
buf ( n10408 , n6590 );
not ( n10409 , n10408 );
not ( n10410 , n8548 );
or ( n10411 , n10409 , n10410 );
or ( n10412 , n8548 , n10408 );
nand ( n10413 , n10411 , n10412 );
buf ( n10414 , n4936 );
buf ( n10415 , n10414 );
not ( n10416 , n10415 );
buf ( n10417 , n4937 );
not ( n10418 , n10417 );
not ( n10419 , n10418 );
or ( n10420 , n10416 , n10419 );
not ( n10421 , n10414 );
buf ( n10422 , n10417 );
nand ( n10423 , n10421 , n10422 );
nand ( n10424 , n10420 , n10423 );
buf ( n10425 , n4938 );
not ( n10426 , n10425 );
and ( n10427 , n10424 , n10426 );
not ( n10428 , n10424 );
buf ( n10429 , n10425 );
and ( n10430 , n10428 , n10429 );
nor ( n10431 , n10427 , n10430 );
buf ( n10432 , n4939 );
nand ( n10433 , n10372 , n10432 );
buf ( n10434 , n4940 );
buf ( n10435 , n10434 );
and ( n10436 , n10433 , n10435 );
not ( n10437 , n10433 );
not ( n10438 , n10434 );
and ( n10439 , n10437 , n10438 );
nor ( n10440 , n10436 , n10439 );
xor ( n10441 , n10431 , n10440 );
xnor ( n10442 , n10441 , n8274 );
buf ( n10443 , n10442 );
and ( n10444 , n10413 , n10443 );
not ( n10445 , n10413 );
not ( n10446 , n10442 );
buf ( n10447 , n10446 );
and ( n10448 , n10445 , n10447 );
nor ( n10449 , n10444 , n10448 );
not ( n10450 , n10449 );
and ( n10451 , n10407 , n10450 );
and ( n10452 , n10406 , n10449 );
nor ( n10453 , n10451 , n10452 );
and ( n10454 , n10238 , n10453 );
not ( n10455 , n10238 );
not ( n10456 , n10453 );
and ( n10457 , n10455 , n10456 );
nor ( n10458 , n10454 , n10457 );
not ( n10459 , n10458 );
not ( n10460 , n10459 );
and ( n10461 , n10023 , n10460 );
and ( n10462 , n10459 , n10022 );
nor ( n10463 , n10461 , n10462 );
not ( n10464 , n10463 );
or ( n10465 , n9385 , n10464 );
not ( n10466 , n9384 );
not ( n10467 , n10459 );
not ( n10468 , n10022 );
or ( n10469 , n10467 , n10468 );
not ( n10470 , n10022 );
nand ( n10471 , n10470 , n10458 );
nand ( n10472 , n10469 , n10471 );
nand ( n10473 , n10466 , n10472 );
nand ( n10474 , n10465 , n10473 );
buf ( n10475 , n4941 );
nand ( n10476 , n7912 , n10475 );
buf ( n10477 , n4942 );
buf ( n10478 , n10477 );
and ( n10479 , n10476 , n10478 );
not ( n10480 , n10476 );
not ( n10481 , n10477 );
and ( n10482 , n10480 , n10481 );
nor ( n10483 , n10479 , n10482 );
not ( n10484 , n10483 );
not ( n10485 , n10089 );
or ( n10486 , n10484 , n10485 );
or ( n10487 , n10089 , n10483 );
nand ( n10488 , n10486 , n10487 );
not ( n10489 , n10488 );
not ( n10490 , n10489 );
not ( n10491 , n10125 );
not ( n10492 , n10491 );
or ( n10493 , n10490 , n10492 );
nand ( n10494 , n10126 , n10488 );
nand ( n10495 , n10493 , n10494 );
not ( n10496 , n10495 );
buf ( n10497 , n4943 );
buf ( n10498 , n10497 );
not ( n10499 , n10498 );
buf ( n10500 , n4944 );
not ( n10501 , n10500 );
not ( n10502 , n10501 );
or ( n10503 , n10499 , n10502 );
not ( n10504 , n10497 );
buf ( n10505 , n10500 );
nand ( n10506 , n10504 , n10505 );
nand ( n10507 , n10503 , n10506 );
buf ( n10508 , n4945 );
buf ( n10509 , n10508 );
and ( n10510 , n10507 , n10509 );
not ( n10511 , n10507 );
not ( n10512 , n10508 );
and ( n10513 , n10511 , n10512 );
nor ( n10514 , n10510 , n10513 );
buf ( n10515 , n4946 );
nand ( n10516 , n7197 , n10515 );
buf ( n10517 , n4947 );
buf ( n10518 , n10517 );
and ( n10519 , n10516 , n10518 );
not ( n10520 , n10516 );
not ( n10521 , n10517 );
and ( n10522 , n10520 , n10521 );
nor ( n10523 , n10519 , n10522 );
xor ( n10524 , n10514 , n10523 );
buf ( n10525 , n4948 );
nand ( n10526 , n8537 , n10525 );
buf ( n10527 , n4949 );
buf ( n10528 , n10527 );
and ( n10529 , n10526 , n10528 );
not ( n10530 , n10526 );
not ( n10531 , n10527 );
and ( n10532 , n10530 , n10531 );
nor ( n10533 , n10529 , n10532 );
xor ( n10534 , n10524 , n10533 );
not ( n10535 , n10534 );
not ( n10536 , n10535 );
buf ( n10537 , n4950 );
buf ( n10538 , n10537 );
not ( n10539 , n10538 );
and ( n10540 , n10536 , n10539 );
not ( n10541 , n10534 );
and ( n10542 , n10541 , n10538 );
nor ( n10543 , n10540 , n10542 );
not ( n10544 , n9950 );
buf ( n10545 , n4951 );
not ( n10546 , n10545 );
not ( n10547 , n10546 );
or ( n10548 , n10544 , n10547 );
not ( n10549 , n9949 );
buf ( n10550 , n10545 );
nand ( n10551 , n10549 , n10550 );
nand ( n10552 , n10548 , n10551 );
buf ( n10553 , n4952 );
not ( n10554 , n10553 );
and ( n10555 , n10552 , n10554 );
not ( n10556 , n10552 );
buf ( n10557 , n10553 );
and ( n10558 , n10556 , n10557 );
nor ( n10559 , n10555 , n10558 );
buf ( n10560 , n4953 );
nand ( n10561 , n6719 , n10560 );
buf ( n10562 , n4954 );
buf ( n10563 , n10562 );
and ( n10564 , n10561 , n10563 );
not ( n10565 , n10561 );
not ( n10566 , n10562 );
and ( n10567 , n10565 , n10566 );
nor ( n10568 , n10564 , n10567 );
xor ( n10569 , n10559 , n10568 );
buf ( n10570 , n7355 );
buf ( n10571 , n4955 );
nand ( n10572 , n10570 , n10571 );
buf ( n10573 , n4956 );
not ( n10574 , n10573 );
and ( n10575 , n10572 , n10574 );
not ( n10576 , n10572 );
buf ( n10577 , n10573 );
and ( n10578 , n10576 , n10577 );
nor ( n10579 , n10575 , n10578 );
xnor ( n10580 , n10569 , n10579 );
buf ( n10581 , n10580 );
and ( n10582 , n10543 , n10581 );
not ( n10583 , n10543 );
not ( n10584 , n10568 );
xor ( n10585 , n10559 , n10584 );
xnor ( n10586 , n10585 , n10579 );
buf ( n10587 , n10586 );
and ( n10588 , n10583 , n10587 );
nor ( n10589 , n10582 , n10588 );
nand ( n10590 , n10496 , n10589 );
not ( n10591 , n10590 );
buf ( n10592 , n4957 );
buf ( n10593 , n10592 );
not ( n10594 , n10593 );
buf ( n10595 , n4958 );
not ( n10596 , n10595 );
not ( n10597 , n10596 );
or ( n10598 , n10594 , n10597 );
not ( n10599 , n10592 );
buf ( n10600 , n10595 );
nand ( n10601 , n10599 , n10600 );
nand ( n10602 , n10598 , n10601 );
not ( n10603 , n10602 );
not ( n10604 , n7759 );
xor ( n10605 , n10604 , n8563 );
buf ( n10606 , n4959 );
nand ( n10607 , n8537 , n10606 );
buf ( n10608 , n4960 );
buf ( n10609 , n10608 );
and ( n10610 , n10607 , n10609 );
not ( n10611 , n10607 );
not ( n10612 , n10608 );
and ( n10613 , n10611 , n10612 );
nor ( n10614 , n10610 , n10613 );
xnor ( n10615 , n10605 , n10614 );
xor ( n10616 , n10603 , n10615 );
not ( n10617 , n10616 );
buf ( n10618 , n4961 );
nand ( n10619 , n6719 , n10618 );
buf ( n10620 , n4962 );
buf ( n10621 , n10620 );
and ( n10622 , n10619 , n10621 );
not ( n10623 , n10619 );
not ( n10624 , n10620 );
and ( n10625 , n10623 , n10624 );
nor ( n10626 , n10622 , n10625 );
buf ( n10627 , n10626 );
not ( n10628 , n10627 );
buf ( n10629 , n4963 );
buf ( n10630 , n10629 );
not ( n10631 , n10630 );
buf ( n10632 , n4964 );
not ( n10633 , n10632 );
not ( n10634 , n10633 );
or ( n10635 , n10631 , n10634 );
not ( n10636 , n10629 );
buf ( n10637 , n10632 );
nand ( n10638 , n10636 , n10637 );
nand ( n10639 , n10635 , n10638 );
buf ( n10640 , n4965 );
not ( n10641 , n10640 );
and ( n10642 , n10639 , n10641 );
not ( n10643 , n10639 );
buf ( n10644 , n10640 );
and ( n10645 , n10643 , n10644 );
nor ( n10646 , n10642 , n10645 );
buf ( n10647 , n4966 );
nand ( n10648 , n6577 , n10647 );
buf ( n10649 , n4967 );
buf ( n10650 , n10649 );
and ( n10651 , n10648 , n10650 );
not ( n10652 , n10648 );
not ( n10653 , n10649 );
and ( n10654 , n10652 , n10653 );
nor ( n10655 , n10651 , n10654 );
xor ( n10656 , n10646 , n10655 );
buf ( n10657 , n4968 );
nand ( n10658 , n6770 , n10657 );
buf ( n10659 , n4969 );
buf ( n10660 , n10659 );
and ( n10661 , n10658 , n10660 );
not ( n10662 , n10658 );
not ( n10663 , n10659 );
and ( n10664 , n10662 , n10663 );
nor ( n10665 , n10661 , n10664 );
xnor ( n10666 , n10656 , n10665 );
not ( n10667 , n10666 );
or ( n10668 , n10628 , n10667 );
or ( n10669 , n10666 , n10627 );
nand ( n10670 , n10668 , n10669 );
not ( n10671 , n10670 );
and ( n10672 , n10617 , n10671 );
not ( n10673 , n10602 );
not ( n10674 , n10615 );
not ( n10675 , n10674 );
or ( n10676 , n10673 , n10675 );
nand ( n10677 , n10615 , n10603 );
nand ( n10678 , n10676 , n10677 );
not ( n10679 , n10678 );
and ( n10680 , n10679 , n10670 );
nor ( n10681 , n10672 , n10680 );
not ( n10682 , n10681 );
not ( n10683 , n10682 );
and ( n10684 , n10591 , n10683 );
and ( n10685 , n10590 , n10682 );
nor ( n10686 , n10684 , n10685 );
not ( n10687 , n10686 );
not ( n10688 , n9839 );
buf ( n10689 , n4970 );
nand ( n10690 , n10372 , n10689 );
buf ( n10691 , n4971 );
xor ( n10692 , n10690 , n10691 );
buf ( n10693 , n10692 );
not ( n10694 , n10693 );
not ( n10695 , n9785 );
not ( n10696 , n10695 );
or ( n10697 , n10694 , n10696 );
or ( n10698 , n10695 , n10693 );
nand ( n10699 , n10697 , n10698 );
not ( n10700 , n10699 );
and ( n10701 , n10688 , n10700 );
and ( n10702 , n9839 , n10699 );
nor ( n10703 , n10701 , n10702 );
buf ( n10704 , n4972 );
buf ( n10705 , n10704 );
not ( n10706 , n10705 );
buf ( n10707 , n4973 );
buf ( n10708 , n10707 );
not ( n10709 , n10708 );
buf ( n10710 , n4974 );
not ( n10711 , n10710 );
not ( n10712 , n10711 );
or ( n10713 , n10709 , n10712 );
not ( n10714 , n10707 );
buf ( n10715 , n10710 );
nand ( n10716 , n10714 , n10715 );
nand ( n10717 , n10713 , n10716 );
buf ( n10718 , n4975 );
not ( n10719 , n10718 );
and ( n10720 , n10717 , n10719 );
not ( n10721 , n10717 );
buf ( n10722 , n10718 );
and ( n10723 , n10721 , n10722 );
nor ( n10724 , n10720 , n10723 );
buf ( n10725 , n4976 );
nand ( n10726 , n7013 , n10725 );
buf ( n10727 , n4977 );
buf ( n10728 , n10727 );
and ( n10729 , n10726 , n10728 );
not ( n10730 , n10726 );
not ( n10731 , n10727 );
and ( n10732 , n10730 , n10731 );
nor ( n10733 , n10729 , n10732 );
xor ( n10734 , n10724 , n10733 );
buf ( n10735 , n4978 );
nand ( n10736 , n6605 , n10735 );
buf ( n10737 , n4979 );
not ( n10738 , n10737 );
and ( n10739 , n10736 , n10738 );
not ( n10740 , n10736 );
buf ( n10741 , n10737 );
and ( n10742 , n10740 , n10741 );
nor ( n10743 , n10739 , n10742 );
xnor ( n10744 , n10734 , n10743 );
not ( n10745 , n10744 );
or ( n10746 , n10706 , n10745 );
not ( n10747 , n10724 );
xor ( n10748 , n10747 , n10733 );
xnor ( n10749 , n10748 , n10743 );
not ( n10750 , n10704 );
nand ( n10751 , n10749 , n10750 );
nand ( n10752 , n10746 , n10751 );
not ( n10753 , n10752 );
not ( n10754 , n9067 );
or ( n10755 , n10753 , n10754 );
or ( n10756 , n9067 , n10752 );
nand ( n10757 , n10755 , n10756 );
buf ( n10758 , n4980 );
nand ( n10759 , n8454 , n10758 );
buf ( n10760 , n4981 );
buf ( n10761 , n10760 );
and ( n10762 , n10759 , n10761 );
not ( n10763 , n10759 );
not ( n10764 , n10760 );
and ( n10765 , n10763 , n10764 );
nor ( n10766 , n10762 , n10765 );
not ( n10767 , n10766 );
not ( n10768 , n8504 );
or ( n10769 , n10767 , n10768 );
or ( n10770 , n8504 , n10766 );
nand ( n10771 , n10769 , n10770 );
not ( n10772 , n10771 );
not ( n10773 , n8547 );
not ( n10774 , n10773 );
not ( n10775 , n10774 );
and ( n10776 , n10772 , n10775 );
and ( n10777 , n10771 , n10774 );
nor ( n10778 , n10776 , n10777 );
nand ( n10779 , n10757 , n10778 );
xor ( n10780 , n10703 , n10779 );
not ( n10781 , n10780 );
or ( n10782 , n10687 , n10781 );
or ( n10783 , n10780 , n10686 );
nand ( n10784 , n10782 , n10783 );
buf ( n10785 , n8721 );
buf ( n10786 , n4982 );
buf ( n10787 , n10786 );
not ( n10788 , n10787 );
buf ( n10789 , n4983 );
not ( n10790 , n10789 );
not ( n10791 , n10790 );
or ( n10792 , n10788 , n10791 );
not ( n10793 , n10786 );
buf ( n10794 , n10789 );
nand ( n10795 , n10793 , n10794 );
nand ( n10796 , n10792 , n10795 );
buf ( n10797 , n4984 );
buf ( n10798 , n10797 );
and ( n10799 , n10796 , n10798 );
not ( n10800 , n10796 );
not ( n10801 , n10797 );
and ( n10802 , n10800 , n10801 );
nor ( n10803 , n10799 , n10802 );
buf ( n10804 , n4985 );
nand ( n10805 , n6828 , n10804 );
buf ( n10806 , n4986 );
buf ( n10807 , n10806 );
and ( n10808 , n10805 , n10807 );
not ( n10809 , n10805 );
not ( n10810 , n10806 );
and ( n10811 , n10809 , n10810 );
nor ( n10812 , n10808 , n10811 );
xor ( n10813 , n10803 , n10812 );
buf ( n10814 , n4987 );
nand ( n10815 , n7344 , n10814 );
buf ( n10816 , n4988 );
buf ( n10817 , n10816 );
and ( n10818 , n10815 , n10817 );
not ( n10819 , n10815 );
not ( n10820 , n10816 );
and ( n10821 , n10819 , n10820 );
nor ( n10822 , n10818 , n10821 );
not ( n10823 , n10822 );
xnor ( n10824 , n10813 , n10823 );
not ( n10825 , n10824 );
not ( n10826 , n10825 );
xor ( n10827 , n10785 , n10826 );
buf ( n10828 , n4989 );
buf ( n10829 , n10828 );
buf ( n10830 , n4990 );
buf ( n10831 , n10830 );
not ( n10832 , n10831 );
buf ( n10833 , n4991 );
not ( n10834 , n10833 );
not ( n10835 , n10834 );
or ( n10836 , n10832 , n10835 );
not ( n10837 , n10830 );
buf ( n10838 , n10833 );
nand ( n10839 , n10837 , n10838 );
nand ( n10840 , n10836 , n10839 );
xor ( n10841 , n10829 , n10840 );
buf ( n10842 , n4992 );
buf ( n10843 , n10842 );
buf ( n10844 , n4993 );
xor ( n10845 , n10843 , n10844 );
buf ( n10846 , n4994 );
nand ( n10847 , n7569 , n10846 );
xnor ( n10848 , n10845 , n10847 );
xnor ( n10849 , n10841 , n10848 );
not ( n10850 , n10849 );
not ( n10851 , n10850 );
xnor ( n10852 , n10827 , n10851 );
not ( n10853 , n10852 );
buf ( n10854 , n4995 );
buf ( n10855 , n10854 );
not ( n10856 , n10855 );
not ( n10857 , n8619 );
or ( n10858 , n10856 , n10857 );
not ( n10859 , n8620 );
not ( n10860 , n10854 );
nand ( n10861 , n10859 , n10860 );
nand ( n10862 , n10858 , n10861 );
not ( n10863 , n10862 );
buf ( n10864 , n8662 );
not ( n10865 , n10864 );
not ( n10866 , n10865 );
and ( n10867 , n10863 , n10866 );
and ( n10868 , n10862 , n10865 );
nor ( n10869 , n10867 , n10868 );
not ( n10870 , n10869 );
nand ( n10871 , n10853 , n10870 );
buf ( n10872 , n4996 );
not ( n10873 , n10872 );
buf ( n10874 , n8176 );
buf ( n10875 , n4997 );
nand ( n10876 , n10874 , n10875 );
buf ( n10877 , n10876 );
not ( n10878 , n10877 );
or ( n10879 , n10873 , n10878 );
or ( n10880 , n10877 , n10872 );
nand ( n10881 , n10879 , n10880 );
not ( n10882 , n10881 );
buf ( n10883 , n4998 );
buf ( n10884 , n10883 );
not ( n10885 , n10884 );
buf ( n10886 , n4999 );
not ( n10887 , n10886 );
not ( n10888 , n10887 );
or ( n10889 , n10885 , n10888 );
not ( n10890 , n10883 );
buf ( n10891 , n10886 );
nand ( n10892 , n10890 , n10891 );
nand ( n10893 , n10889 , n10892 );
buf ( n10894 , n5000 );
buf ( n10895 , n10894 );
and ( n10896 , n10893 , n10895 );
not ( n10897 , n10893 );
not ( n10898 , n10894 );
and ( n10899 , n10897 , n10898 );
nor ( n10900 , n10896 , n10899 );
buf ( n10901 , n5001 );
nand ( n10902 , n7293 , n10901 );
buf ( n10903 , n5002 );
buf ( n10904 , n10903 );
and ( n10905 , n10902 , n10904 );
not ( n10906 , n10902 );
not ( n10907 , n10903 );
and ( n10908 , n10906 , n10907 );
nor ( n10909 , n10905 , n10908 );
xor ( n10910 , n10900 , n10909 );
xnor ( n10911 , n10910 , n9196 );
buf ( n10912 , n10911 );
not ( n10913 , n10912 );
or ( n10914 , n10882 , n10913 );
not ( n10915 , n10881 );
not ( n10916 , n10911 );
nand ( n10917 , n10915 , n10916 );
nand ( n10918 , n10914 , n10917 );
buf ( n10919 , n5003 );
buf ( n10920 , n10919 );
not ( n10921 , n10920 );
buf ( n10922 , n5004 );
not ( n10923 , n10922 );
not ( n10924 , n10923 );
or ( n10925 , n10921 , n10924 );
not ( n10926 , n10919 );
buf ( n10927 , n10922 );
nand ( n10928 , n10926 , n10927 );
nand ( n10929 , n10925 , n10928 );
buf ( n10930 , n5005 );
buf ( n10931 , n10930 );
and ( n10932 , n10929 , n10931 );
not ( n10933 , n10929 );
not ( n10934 , n10930 );
and ( n10935 , n10933 , n10934 );
nor ( n10936 , n10932 , n10935 );
buf ( n10937 , n5006 );
nand ( n10938 , n7202 , n10937 );
buf ( n10939 , n5007 );
buf ( n10940 , n10939 );
and ( n10941 , n10938 , n10940 );
not ( n10942 , n10938 );
not ( n10943 , n10939 );
and ( n10944 , n10942 , n10943 );
nor ( n10945 , n10941 , n10944 );
xor ( n10946 , n10936 , n10945 );
buf ( n10947 , n9160 );
buf ( n10948 , n5008 );
nand ( n10949 , n10947 , n10948 );
buf ( n10950 , n5009 );
buf ( n10951 , n10950 );
and ( n10952 , n10949 , n10951 );
not ( n10953 , n10949 );
not ( n10954 , n10950 );
and ( n10955 , n10953 , n10954 );
nor ( n10956 , n10952 , n10955 );
xnor ( n10957 , n10946 , n10956 );
buf ( n10958 , n10957 );
buf ( n10959 , n10958 );
not ( n10960 , n10959 );
and ( n10961 , n10918 , n10960 );
not ( n10962 , n10918 );
and ( n10963 , n10962 , n10959 );
nor ( n10964 , n10961 , n10963 );
buf ( n10965 , n10964 );
not ( n10966 , n10965 );
and ( n10967 , n10871 , n10966 );
not ( n10968 , n10871 );
and ( n10969 , n10968 , n10965 );
nor ( n10970 , n10967 , n10969 );
and ( n10971 , n10784 , n10970 );
not ( n10972 , n10784 );
not ( n10973 , n10970 );
and ( n10974 , n10972 , n10973 );
nor ( n10975 , n10971 , n10974 );
not ( n10976 , n10975 );
not ( n10977 , n10976 );
buf ( n10978 , n5010 );
not ( n10979 , n9655 );
buf ( n10980 , n5011 );
not ( n10981 , n10980 );
not ( n10982 , n10981 );
or ( n10983 , n10979 , n10982 );
not ( n10984 , n9654 );
buf ( n10985 , n10980 );
nand ( n10986 , n10984 , n10985 );
nand ( n10987 , n10983 , n10986 );
buf ( n10988 , n5012 );
buf ( n10989 , n10988 );
and ( n10990 , n10987 , n10989 );
not ( n10991 , n10987 );
not ( n10992 , n10988 );
and ( n10993 , n10991 , n10992 );
nor ( n10994 , n10990 , n10993 );
buf ( n10995 , n5013 );
nand ( n10996 , n6634 , n10995 );
buf ( n10997 , n5014 );
buf ( n10998 , n10997 );
and ( n10999 , n10996 , n10998 );
not ( n11000 , n10996 );
not ( n11001 , n10997 );
and ( n11002 , n11000 , n11001 );
nor ( n11003 , n10999 , n11002 );
xor ( n11004 , n10994 , n11003 );
buf ( n11005 , n5015 );
nand ( n11006 , n7247 , n11005 );
buf ( n11007 , n5016 );
buf ( n11008 , n11007 );
and ( n11009 , n11006 , n11008 );
not ( n11010 , n11006 );
not ( n11011 , n11007 );
and ( n11012 , n11010 , n11011 );
nor ( n11013 , n11009 , n11012 );
not ( n11014 , n11013 );
xnor ( n11015 , n11004 , n11014 );
xor ( n11016 , n10978 , n11015 );
buf ( n11017 , n5017 );
buf ( n11018 , n11017 );
not ( n11019 , n11018 );
buf ( n11020 , n5018 );
not ( n11021 , n11020 );
not ( n11022 , n11021 );
or ( n11023 , n11019 , n11022 );
not ( n11024 , n11017 );
buf ( n11025 , n11020 );
nand ( n11026 , n11024 , n11025 );
nand ( n11027 , n11023 , n11026 );
buf ( n11028 , n5019 );
buf ( n11029 , n11028 );
and ( n11030 , n11027 , n11029 );
not ( n11031 , n11027 );
not ( n11032 , n11028 );
and ( n11033 , n11031 , n11032 );
nor ( n11034 , n11030 , n11033 );
buf ( n11035 , n5020 );
nand ( n11036 , n7107 , n11035 );
buf ( n11037 , n5021 );
buf ( n11038 , n11037 );
and ( n11039 , n11036 , n11038 );
not ( n11040 , n11036 );
not ( n11041 , n11037 );
and ( n11042 , n11040 , n11041 );
nor ( n11043 , n11039 , n11042 );
xor ( n11044 , n11034 , n11043 );
buf ( n11045 , n5022 );
nand ( n11046 , n8675 , n11045 );
buf ( n11047 , n5023 );
buf ( n11048 , n11047 );
and ( n11049 , n11046 , n11048 );
not ( n11050 , n11046 );
not ( n11051 , n11047 );
and ( n11052 , n11050 , n11051 );
nor ( n11053 , n11049 , n11052 );
xnor ( n11054 , n11044 , n11053 );
not ( n11055 , n11054 );
xnor ( n11056 , n11016 , n11055 );
not ( n11057 , n11056 );
not ( n11058 , n11057 );
buf ( n11059 , n5024 );
buf ( n11060 , n11059 );
not ( n11061 , n11060 );
buf ( n11062 , n5025 );
not ( n11063 , n11062 );
buf ( n11064 , n5026 );
buf ( n11065 , n11064 );
not ( n11066 , n11065 );
buf ( n11067 , n5027 );
not ( n11068 , n11067 );
not ( n11069 , n11068 );
or ( n11070 , n11066 , n11069 );
not ( n11071 , n11064 );
buf ( n11072 , n11067 );
nand ( n11073 , n11071 , n11072 );
nand ( n11074 , n11070 , n11073 );
xor ( n11075 , n11063 , n11074 );
buf ( n11076 , n5028 );
buf ( n11077 , n5029 );
xor ( n11078 , n11076 , n11077 );
buf ( n11079 , n5030 );
nand ( n11080 , n7197 , n11079 );
xnor ( n11081 , n11078 , n11080 );
xor ( n11082 , n11075 , n11081 );
not ( n11083 , n11082 );
or ( n11084 , n11061 , n11083 );
or ( n11085 , n11082 , n11060 );
nand ( n11086 , n11084 , n11085 );
not ( n11087 , n11086 );
not ( n11088 , n6937 );
not ( n11089 , n11088 );
not ( n11090 , n11089 );
and ( n11091 , n11087 , n11090 );
and ( n11092 , n11086 , n11089 );
nor ( n11093 , n11091 , n11092 );
not ( n11094 , n11093 );
nand ( n11095 , n11058 , n11094 );
not ( n11096 , n11095 );
not ( n11097 , n8079 );
not ( n11098 , n6730 );
or ( n11099 , n11097 , n11098 );
or ( n11100 , n6730 , n8079 );
nand ( n11101 , n11099 , n11100 );
not ( n11102 , n11101 );
xor ( n11103 , n6668 , n6677 );
xnor ( n11104 , n11103 , n6684 );
not ( n11105 , n11104 );
not ( n11106 , n11105 );
or ( n11107 , n11102 , n11106 );
not ( n11108 , n6685 );
or ( n11109 , n11108 , n11101 );
nand ( n11110 , n11107 , n11109 );
buf ( n11111 , n11110 );
not ( n11112 , n11111 );
and ( n11113 , n11096 , n11112 );
and ( n11114 , n11095 , n11111 );
nor ( n11115 , n11113 , n11114 );
not ( n11116 , n11115 );
buf ( n11117 , n10392 );
not ( n11118 , n11117 );
not ( n11119 , n7808 );
xor ( n11120 , n11119 , n7820 );
xor ( n11121 , n11120 , n7827 );
not ( n11122 , n11121 );
not ( n11123 , n11122 );
or ( n11124 , n11118 , n11123 );
or ( n11125 , n11122 , n11117 );
nand ( n11126 , n11124 , n11125 );
buf ( n11127 , n5031 );
buf ( n11128 , n11127 );
not ( n11129 , n11128 );
buf ( n11130 , n5032 );
not ( n11131 , n11130 );
not ( n11132 , n11131 );
or ( n11133 , n11129 , n11132 );
not ( n11134 , n11127 );
buf ( n11135 , n11130 );
nand ( n11136 , n11134 , n11135 );
nand ( n11137 , n11133 , n11136 );
not ( n11138 , n9745 );
and ( n11139 , n11137 , n11138 );
not ( n11140 , n11137 );
and ( n11141 , n11140 , n9746 );
nor ( n11142 , n11139 , n11141 );
xor ( n11143 , n11142 , n10692 );
buf ( n11144 , n5033 );
nand ( n11145 , n10570 , n11144 );
buf ( n11146 , n5034 );
not ( n11147 , n11146 );
and ( n11148 , n11145 , n11147 );
not ( n11149 , n11145 );
buf ( n11150 , n11146 );
and ( n11151 , n11149 , n11150 );
nor ( n11152 , n11148 , n11151 );
xnor ( n11153 , n11143 , n11152 );
buf ( n11154 , n11153 );
buf ( n11155 , n11154 );
not ( n11156 , n11155 );
and ( n11157 , n11126 , n11156 );
not ( n11158 , n11126 );
and ( n11159 , n11158 , n11155 );
nor ( n11160 , n11157 , n11159 );
not ( n11161 , n11160 );
not ( n11162 , n9462 );
not ( n11163 , n11162 );
buf ( n11164 , n5035 );
not ( n11165 , n11164 );
buf ( n11166 , n5036 );
nand ( n11167 , n7912 , n11166 );
not ( n11168 , n11167 );
or ( n11169 , n11165 , n11168 );
nand ( n11170 , n8070 , n11166 );
or ( n11171 , n11170 , n11164 );
nand ( n11172 , n11169 , n11171 );
not ( n11173 , n11172 );
not ( n11174 , n9419 );
not ( n11175 , n11174 );
not ( n11176 , n11175 );
or ( n11177 , n11173 , n11176 );
not ( n11178 , n11172 );
nand ( n11179 , n11174 , n11178 );
nand ( n11180 , n11177 , n11179 );
not ( n11181 , n11180 );
or ( n11182 , n11163 , n11181 );
or ( n11183 , n11180 , n9465 );
nand ( n11184 , n11182 , n11183 );
not ( n11185 , n11184 );
buf ( n11186 , n5037 );
buf ( n11187 , n11186 );
not ( n11188 , n11187 );
buf ( n11189 , n5038 );
buf ( n11190 , n11189 );
not ( n11191 , n11190 );
buf ( n11192 , n5039 );
not ( n11193 , n11192 );
not ( n11194 , n11193 );
or ( n11195 , n11191 , n11194 );
not ( n11196 , n11189 );
buf ( n11197 , n11192 );
nand ( n11198 , n11196 , n11197 );
nand ( n11199 , n11195 , n11198 );
buf ( n11200 , n5040 );
not ( n11201 , n11200 );
and ( n11202 , n11199 , n11201 );
not ( n11203 , n11199 );
buf ( n11204 , n11200 );
and ( n11205 , n11203 , n11204 );
nor ( n11206 , n11202 , n11205 );
buf ( n11207 , n5041 );
nand ( n11208 , n6604 , n11207 );
buf ( n11209 , n5042 );
buf ( n11210 , n11209 );
and ( n11211 , n11208 , n11210 );
not ( n11212 , n11208 );
not ( n11213 , n11209 );
and ( n11214 , n11212 , n11213 );
nor ( n11215 , n11211 , n11214 );
xor ( n11216 , n11206 , n11215 );
buf ( n11217 , n5043 );
nand ( n11218 , n8375 , n11217 );
buf ( n11219 , n5044 );
not ( n11220 , n11219 );
and ( n11221 , n11218 , n11220 );
not ( n11222 , n11218 );
buf ( n11223 , n11219 );
and ( n11224 , n11222 , n11223 );
nor ( n11225 , n11221 , n11224 );
xnor ( n11226 , n11216 , n11225 );
not ( n11227 , n11226 );
not ( n11228 , n11227 );
not ( n11229 , n11228 );
or ( n11230 , n11188 , n11229 );
not ( n11231 , n11187 );
nand ( n11232 , n11231 , n11227 );
nand ( n11233 , n11230 , n11232 );
buf ( n11234 , n5045 );
buf ( n11235 , n11234 );
not ( n11236 , n11235 );
buf ( n11237 , n5046 );
not ( n11238 , n11237 );
not ( n11239 , n11238 );
or ( n11240 , n11236 , n11239 );
not ( n11241 , n11234 );
buf ( n11242 , n11237 );
nand ( n11243 , n11241 , n11242 );
nand ( n11244 , n11240 , n11243 );
buf ( n11245 , n5047 );
buf ( n11246 , n11245 );
and ( n11247 , n11244 , n11246 );
not ( n11248 , n11244 );
not ( n11249 , n11245 );
and ( n11250 , n11248 , n11249 );
nor ( n11251 , n11247 , n11250 );
buf ( n11252 , n5048 );
nand ( n11253 , n8454 , n11252 );
buf ( n11254 , n5049 );
buf ( n11255 , n11254 );
and ( n11256 , n11253 , n11255 );
not ( n11257 , n11253 );
not ( n11258 , n11254 );
and ( n11259 , n11257 , n11258 );
nor ( n11260 , n11256 , n11259 );
xor ( n11261 , n11251 , n11260 );
buf ( n11262 , n5050 );
nand ( n11263 , n9310 , n11262 );
buf ( n11264 , n5051 );
buf ( n11265 , n11264 );
and ( n11266 , n11263 , n11265 );
not ( n11267 , n11263 );
not ( n11268 , n11264 );
and ( n11269 , n11267 , n11268 );
nor ( n11270 , n11266 , n11269 );
xnor ( n11271 , n11261 , n11270 );
buf ( n11272 , n11271 );
and ( n11273 , n11233 , n11272 );
not ( n11274 , n11233 );
not ( n11275 , n11272 );
and ( n11276 , n11274 , n11275 );
nor ( n11277 , n11273 , n11276 );
not ( n11278 , n11277 );
nand ( n11279 , n11185 , n11278 );
not ( n11280 , n11279 );
or ( n11281 , n11161 , n11280 );
or ( n11282 , n11279 , n11160 );
nand ( n11283 , n11281 , n11282 );
not ( n11284 , n11283 );
and ( n11285 , n11116 , n11284 );
and ( n11286 , n11115 , n11283 );
nor ( n11287 , n11285 , n11286 );
not ( n11288 , n11287 );
not ( n11289 , n11288 );
and ( n11290 , n10977 , n11289 );
and ( n11291 , n10976 , n11288 );
nor ( n11292 , n11290 , n11291 );
buf ( n11293 , n11292 );
and ( n11294 , n10474 , n11293 );
not ( n11295 , n10474 );
not ( n11296 , n11287 );
not ( n11297 , n10975 );
or ( n11298 , n11296 , n11297 );
not ( n11299 , n11287 );
nand ( n11300 , n11299 , n10976 );
nand ( n11301 , n11298 , n11300 );
buf ( n11302 , n11301 );
and ( n11303 , n11295 , n11302 );
nor ( n11304 , n11294 , n11303 );
xor ( n11305 , n8245 , n8254 );
xnor ( n11306 , n11305 , n8263 );
buf ( n11307 , n11306 );
not ( n11308 , n8517 );
buf ( n11309 , n5052 );
buf ( n11310 , n11309 );
not ( n11311 , n11310 );
buf ( n11312 , n5053 );
not ( n11313 , n11312 );
not ( n11314 , n11313 );
or ( n11315 , n11311 , n11314 );
not ( n11316 , n11309 );
buf ( n11317 , n11312 );
nand ( n11318 , n11316 , n11317 );
nand ( n11319 , n11315 , n11318 );
buf ( n11320 , n5054 );
buf ( n11321 , n11320 );
and ( n11322 , n11319 , n11321 );
not ( n11323 , n11319 );
not ( n11324 , n11320 );
and ( n11325 , n11323 , n11324 );
nor ( n11326 , n11322 , n11325 );
buf ( n11327 , n5055 );
nand ( n11328 , n7202 , n11327 );
buf ( n11329 , n5056 );
not ( n11330 , n11329 );
and ( n11331 , n11328 , n11330 );
not ( n11332 , n11328 );
buf ( n11333 , n11329 );
and ( n11334 , n11332 , n11333 );
nor ( n11335 , n11331 , n11334 );
xor ( n11336 , n11326 , n11335 );
buf ( n11337 , n7606 );
buf ( n11338 , n5057 );
nand ( n11339 , n11337 , n11338 );
buf ( n11340 , n5058 );
not ( n11341 , n11340 );
and ( n11342 , n11339 , n11341 );
not ( n11343 , n11339 );
buf ( n11344 , n11340 );
and ( n11345 , n11343 , n11344 );
nor ( n11346 , n11342 , n11345 );
xnor ( n11347 , n11336 , n11346 );
buf ( n11348 , n11347 );
not ( n11349 , n11348 );
or ( n11350 , n11308 , n11349 );
or ( n11351 , n11348 , n8517 );
nand ( n11352 , n11350 , n11351 );
and ( n11353 , n11307 , n11352 );
not ( n11354 , n11307 );
not ( n11355 , n11352 );
and ( n11356 , n11354 , n11355 );
nor ( n11357 , n11353 , n11356 );
buf ( n11358 , n5059 );
nand ( n11359 , n10947 , n11358 );
buf ( n11360 , n5060 );
not ( n11361 , n11360 );
and ( n11362 , n11359 , n11361 );
not ( n11363 , n11359 );
buf ( n11364 , n11360 );
and ( n11365 , n11363 , n11364 );
nor ( n11366 , n11362 , n11365 );
not ( n11367 , n11366 );
buf ( n11368 , n5061 );
buf ( n11369 , n11368 );
not ( n11370 , n11369 );
not ( n11371 , n6845 );
or ( n11372 , n11370 , n11371 );
not ( n11373 , n11368 );
nand ( n11374 , n11373 , n6795 );
nand ( n11375 , n11372 , n11374 );
buf ( n11376 , n5062 );
buf ( n11377 , n11376 );
and ( n11378 , n11375 , n11377 );
not ( n11379 , n11375 );
not ( n11380 , n11376 );
and ( n11381 , n11379 , n11380 );
nor ( n11382 , n11378 , n11381 );
buf ( n11383 , n5063 );
nand ( n11384 , n6927 , n11383 );
buf ( n11385 , n5064 );
buf ( n11386 , n11385 );
and ( n11387 , n11384 , n11386 );
not ( n11388 , n11384 );
not ( n11389 , n11385 );
and ( n11390 , n11388 , n11389 );
nor ( n11391 , n11387 , n11390 );
xor ( n11392 , n11382 , n11391 );
xor ( n11393 , n11392 , n8332 );
buf ( n11394 , n11393 );
not ( n11395 , n11394 );
or ( n11396 , n11367 , n11395 );
or ( n11397 , n11366 , n11394 );
nand ( n11398 , n11396 , n11397 );
buf ( n11399 , n5065 );
buf ( n11400 , n11399 );
not ( n11401 , n11400 );
buf ( n11402 , n5066 );
not ( n11403 , n11402 );
not ( n11404 , n11403 );
or ( n11405 , n11401 , n11404 );
not ( n11406 , n11399 );
buf ( n11407 , n11402 );
nand ( n11408 , n11406 , n11407 );
nand ( n11409 , n11405 , n11408 );
buf ( n11410 , n5067 );
not ( n11411 , n11410 );
and ( n11412 , n11409 , n11411 );
not ( n11413 , n11409 );
buf ( n11414 , n11410 );
and ( n11415 , n11413 , n11414 );
nor ( n11416 , n11412 , n11415 );
buf ( n11417 , n5068 );
nand ( n11418 , n9812 , n11417 );
buf ( n11419 , n5069 );
buf ( n11420 , n11419 );
and ( n11421 , n11418 , n11420 );
not ( n11422 , n11418 );
not ( n11423 , n11419 );
and ( n11424 , n11422 , n11423 );
nor ( n11425 , n11421 , n11424 );
xor ( n11426 , n11416 , n11425 );
buf ( n11427 , n5070 );
nand ( n11428 , n11337 , n11427 );
buf ( n11429 , n5071 );
not ( n11430 , n11429 );
and ( n11431 , n11428 , n11430 );
not ( n11432 , n11428 );
buf ( n11433 , n11429 );
and ( n11434 , n11432 , n11433 );
nor ( n11435 , n11431 , n11434 );
xnor ( n11436 , n11426 , n11435 );
buf ( n11437 , n11436 );
buf ( n11438 , n11437 );
and ( n11439 , n11398 , n11438 );
not ( n11440 , n11398 );
not ( n11441 , n11438 );
and ( n11442 , n11440 , n11441 );
nor ( n11443 , n11439 , n11442 );
nand ( n11444 , n11357 , n11443 );
not ( n11445 , n11444 );
buf ( n11446 , n5072 );
nand ( n11447 , n6515 , n11446 );
buf ( n11448 , n5073 );
buf ( n11449 , n11448 );
and ( n11450 , n11447 , n11449 );
not ( n11451 , n11447 );
not ( n11452 , n11448 );
and ( n11453 , n11451 , n11452 );
nor ( n11454 , n11450 , n11453 );
not ( n11455 , n11454 );
not ( n11456 , n11455 );
not ( n11457 , n7411 );
or ( n11458 , n11456 , n11457 );
not ( n11459 , n11455 );
not ( n11460 , n7411 );
nand ( n11461 , n11459 , n11460 );
nand ( n11462 , n11458 , n11461 );
buf ( n11463 , n5074 );
buf ( n11464 , n11463 );
not ( n11465 , n11464 );
buf ( n11466 , n5075 );
not ( n11467 , n11466 );
not ( n11468 , n11467 );
or ( n11469 , n11465 , n11468 );
not ( n11470 , n11463 );
buf ( n11471 , n11466 );
nand ( n11472 , n11470 , n11471 );
nand ( n11473 , n11469 , n11472 );
buf ( n11474 , n5076 );
not ( n11475 , n11474 );
and ( n11476 , n11473 , n11475 );
not ( n11477 , n11473 );
buf ( n11478 , n11474 );
and ( n11479 , n11477 , n11478 );
nor ( n11480 , n11476 , n11479 );
buf ( n11481 , n5077 );
nand ( n11482 , n7787 , n11481 );
buf ( n11483 , n5078 );
not ( n11484 , n11483 );
and ( n11485 , n11482 , n11484 );
not ( n11486 , n11482 );
buf ( n11487 , n11483 );
and ( n11488 , n11486 , n11487 );
nor ( n11489 , n11485 , n11488 );
xor ( n11490 , n11480 , n11489 );
buf ( n11491 , n5079 );
nand ( n11492 , n7247 , n11491 );
buf ( n11493 , n5080 );
buf ( n11494 , n11493 );
and ( n11495 , n11492 , n11494 );
not ( n11496 , n11492 );
not ( n11497 , n11493 );
and ( n11498 , n11496 , n11497 );
nor ( n11499 , n11495 , n11498 );
xor ( n11500 , n11490 , n11499 );
not ( n11501 , n11500 );
buf ( n11502 , n11501 );
not ( n11503 , n11502 );
and ( n11504 , n11462 , n11503 );
not ( n11505 , n11462 );
not ( n11506 , n11500 );
buf ( n11507 , n11506 );
not ( n11508 , n11507 );
not ( n11509 , n11508 );
and ( n11510 , n11505 , n11509 );
nor ( n11511 , n11504 , n11510 );
not ( n11512 , n11511 );
not ( n11513 , n11512 );
not ( n11514 , n11513 );
and ( n11515 , n11445 , n11514 );
and ( n11516 , n11444 , n11513 );
nor ( n11517 , n11515 , n11516 );
not ( n11518 , n11517 );
not ( n11519 , n11518 );
buf ( n11520 , n5081 );
nand ( n11521 , n8675 , n11520 );
buf ( n11522 , n5082 );
not ( n11523 , n11522 );
and ( n11524 , n11521 , n11523 );
not ( n11525 , n11521 );
buf ( n11526 , n11522 );
and ( n11527 , n11525 , n11526 );
nor ( n11528 , n11524 , n11527 );
buf ( n11529 , n5083 );
buf ( n11530 , n5084 );
not ( n11531 , n11530 );
nand ( n11532 , n11531 , n7324 );
not ( n11533 , n7323 );
buf ( n11534 , n11530 );
nand ( n11535 , n11533 , n11534 );
and ( n11536 , n11532 , n11535 );
xor ( n11537 , n11529 , n11536 );
buf ( n11538 , n5085 );
buf ( n11539 , n5086 );
xor ( n11540 , n11538 , n11539 );
buf ( n11541 , n5087 );
nand ( n11542 , n7709 , n11541 );
xnor ( n11543 , n11540 , n11542 );
xnor ( n11544 , n11537 , n11543 );
xor ( n11545 , n11528 , n11544 );
buf ( n11546 , n5088 );
buf ( n11547 , n11546 );
not ( n11548 , n11547 );
buf ( n11549 , n5089 );
not ( n11550 , n11549 );
not ( n11551 , n11550 );
or ( n11552 , n11548 , n11551 );
not ( n11553 , n11546 );
buf ( n11554 , n11549 );
nand ( n11555 , n11553 , n11554 );
nand ( n11556 , n11552 , n11555 );
buf ( n11557 , n5090 );
not ( n11558 , n11557 );
and ( n11559 , n11556 , n11558 );
not ( n11560 , n11556 );
buf ( n11561 , n11557 );
and ( n11562 , n11560 , n11561 );
nor ( n11563 , n11559 , n11562 );
xor ( n11564 , n11563 , n11454 );
buf ( n11565 , n5091 );
nand ( n11566 , n6647 , n11565 );
buf ( n11567 , n5092 );
buf ( n11568 , n11567 );
and ( n11569 , n11566 , n11568 );
not ( n11570 , n11566 );
not ( n11571 , n11567 );
and ( n11572 , n11570 , n11571 );
nor ( n11573 , n11569 , n11572 );
not ( n11574 , n11573 );
xnor ( n11575 , n11564 , n11574 );
xnor ( n11576 , n11545 , n11575 );
not ( n11577 , n11576 );
not ( n11578 , n7466 );
buf ( n11579 , n5093 );
buf ( n11580 , n11579 );
not ( n11581 , n11580 );
buf ( n11582 , n5094 );
not ( n11583 , n11582 );
not ( n11584 , n11583 );
or ( n11585 , n11581 , n11584 );
not ( n11586 , n11579 );
buf ( n11587 , n11582 );
nand ( n11588 , n11586 , n11587 );
nand ( n11589 , n11585 , n11588 );
not ( n11590 , n9005 );
and ( n11591 , n11589 , n11590 );
not ( n11592 , n11589 );
and ( n11593 , n11592 , n9006 );
nor ( n11594 , n11591 , n11593 );
buf ( n11595 , n5095 );
nand ( n11596 , n6633 , n11595 );
buf ( n11597 , n5096 );
buf ( n11598 , n11597 );
and ( n11599 , n11596 , n11598 );
not ( n11600 , n11596 );
not ( n11601 , n11597 );
and ( n11602 , n11600 , n11601 );
nor ( n11603 , n11599 , n11602 );
xor ( n11604 , n11594 , n11603 );
buf ( n11605 , n5097 );
nand ( n11606 , n8781 , n11605 );
buf ( n11607 , n5098 );
not ( n11608 , n11607 );
and ( n11609 , n11606 , n11608 );
not ( n11610 , n11606 );
buf ( n11611 , n11607 );
and ( n11612 , n11610 , n11611 );
nor ( n11613 , n11609 , n11612 );
xnor ( n11614 , n11604 , n11613 );
not ( n11615 , n11614 );
not ( n11616 , n11615 );
or ( n11617 , n11578 , n11616 );
or ( n11618 , n11615 , n7466 );
nand ( n11619 , n11617 , n11618 );
buf ( n11620 , n9235 );
and ( n11621 , n11619 , n11620 );
not ( n11622 , n11619 );
not ( n11623 , n11620 );
and ( n11624 , n11622 , n11623 );
nor ( n11625 , n11621 , n11624 );
not ( n11626 , n11625 );
nand ( n11627 , n11577 , n11626 );
buf ( n11628 , n5099 );
not ( n11629 , n11628 );
buf ( n11630 , n5100 );
nand ( n11631 , n7293 , n11630 );
buf ( n11632 , n5101 );
buf ( n11633 , n11632 );
and ( n11634 , n11631 , n11633 );
not ( n11635 , n11631 );
not ( n11636 , n11632 );
and ( n11637 , n11635 , n11636 );
nor ( n11638 , n11634 , n11637 );
not ( n11639 , n11638 );
buf ( n11640 , n5102 );
nand ( n11641 , n8070 , n11640 );
buf ( n11642 , n5103 );
not ( n11643 , n11642 );
and ( n11644 , n11641 , n11643 );
not ( n11645 , n11641 );
buf ( n11646 , n11642 );
and ( n11647 , n11645 , n11646 );
nor ( n11648 , n11644 , n11647 );
not ( n11649 , n11648 );
or ( n11650 , n11639 , n11649 );
or ( n11651 , n11638 , n11648 );
nand ( n11652 , n11650 , n11651 );
buf ( n11653 , n5104 );
buf ( n11654 , n11653 );
not ( n11655 , n11654 );
buf ( n11656 , n5105 );
not ( n11657 , n11656 );
not ( n11658 , n11657 );
or ( n11659 , n11655 , n11658 );
not ( n11660 , n11653 );
buf ( n11661 , n11656 );
nand ( n11662 , n11660 , n11661 );
nand ( n11663 , n11659 , n11662 );
buf ( n11664 , n5106 );
buf ( n11665 , n11664 );
and ( n11666 , n11663 , n11665 );
not ( n11667 , n11663 );
not ( n11668 , n11664 );
and ( n11669 , n11667 , n11668 );
nor ( n11670 , n11666 , n11669 );
not ( n11671 , n11670 );
xor ( n11672 , n11652 , n11671 );
not ( n11673 , n11672 );
or ( n11674 , n11629 , n11673 );
or ( n11675 , n11672 , n11628 );
nand ( n11676 , n11674 , n11675 );
not ( n11677 , n11676 );
buf ( n11678 , n5107 );
nand ( n11679 , n8781 , n11678 );
buf ( n11680 , n5108 );
buf ( n11681 , n11680 );
and ( n11682 , n11679 , n11681 );
not ( n11683 , n11679 );
not ( n11684 , n11680 );
and ( n11685 , n11683 , n11684 );
nor ( n11686 , n11682 , n11685 );
not ( n11687 , n11686 );
buf ( n11688 , n7293 );
buf ( n11689 , n5109 );
nand ( n11690 , n11688 , n11689 );
buf ( n11691 , n5110 );
not ( n11692 , n11691 );
and ( n11693 , n11690 , n11692 );
not ( n11694 , n11690 );
buf ( n11695 , n11691 );
and ( n11696 , n11694 , n11695 );
nor ( n11697 , n11693 , n11696 );
not ( n11698 , n11697 );
or ( n11699 , n11687 , n11698 );
or ( n11700 , n11686 , n11697 );
nand ( n11701 , n11699 , n11700 );
buf ( n11702 , n5111 );
buf ( n11703 , n11702 );
not ( n11704 , n11703 );
buf ( n11705 , n5112 );
not ( n11706 , n11705 );
not ( n11707 , n11706 );
or ( n11708 , n11704 , n11707 );
not ( n11709 , n11702 );
buf ( n11710 , n11705 );
nand ( n11711 , n11709 , n11710 );
nand ( n11712 , n11708 , n11711 );
buf ( n11713 , n5113 );
not ( n11714 , n11713 );
and ( n11715 , n11712 , n11714 );
not ( n11716 , n11712 );
buf ( n11717 , n11713 );
and ( n11718 , n11716 , n11717 );
nor ( n11719 , n11715 , n11718 );
and ( n11720 , n11701 , n11719 );
not ( n11721 , n11701 );
not ( n11722 , n11719 );
and ( n11723 , n11721 , n11722 );
nor ( n11724 , n11720 , n11723 );
not ( n11725 , n11724 );
and ( n11726 , n11677 , n11725 );
buf ( n11727 , n11724 );
and ( n11728 , n11676 , n11727 );
nor ( n11729 , n11726 , n11728 );
not ( n11730 , n11729 );
xnor ( n11731 , n11627 , n11730 );
not ( n11732 , n11731 );
not ( n11733 , n11732 );
buf ( n11734 , n5114 );
buf ( n11735 , n5115 );
buf ( n11736 , n11735 );
not ( n11737 , n11736 );
buf ( n11738 , n5116 );
not ( n11739 , n11738 );
not ( n11740 , n11739 );
or ( n11741 , n11737 , n11740 );
not ( n11742 , n11735 );
buf ( n11743 , n11738 );
nand ( n11744 , n11742 , n11743 );
nand ( n11745 , n11741 , n11744 );
xor ( n11746 , n11734 , n11745 );
buf ( n11747 , n5117 );
buf ( n11748 , n5118 );
buf ( n11749 , n11748 );
xor ( n11750 , n11747 , n11749 );
buf ( n11751 , n5119 );
nand ( n11752 , n8675 , n11751 );
xnor ( n11753 , n11750 , n11752 );
not ( n11754 , n11753 );
xnor ( n11755 , n11746 , n11754 );
not ( n11756 , n11755 );
not ( n11757 , n7313 );
not ( n11758 , n11757 );
buf ( n11759 , n5120 );
nand ( n11760 , n8124 , n11759 );
buf ( n11761 , n5121 );
buf ( n11762 , n11761 );
and ( n11763 , n11760 , n11762 );
not ( n11764 , n11760 );
not ( n11765 , n11761 );
and ( n11766 , n11764 , n11765 );
nor ( n11767 , n11763 , n11766 );
buf ( n11768 , n11767 );
not ( n11769 , n11768 );
and ( n11770 , n11758 , n11769 );
and ( n11771 , n11757 , n11768 );
nor ( n11772 , n11770 , n11771 );
not ( n11773 , n11772 );
or ( n11774 , n11756 , n11773 );
buf ( n11775 , n11755 );
or ( n11776 , n11775 , n11772 );
nand ( n11777 , n11774 , n11776 );
not ( n11778 , n11777 );
buf ( n11779 , n5122 );
buf ( n11780 , n11779 );
not ( n11781 , n11780 );
buf ( n11782 , n5123 );
not ( n11783 , n11782 );
not ( n11784 , n11783 );
or ( n11785 , n11781 , n11784 );
not ( n11786 , n11779 );
buf ( n11787 , n11782 );
nand ( n11788 , n11786 , n11787 );
nand ( n11789 , n11785 , n11788 );
buf ( n11790 , n5124 );
buf ( n11791 , n11790 );
and ( n11792 , n11789 , n11791 );
not ( n11793 , n11789 );
not ( n11794 , n11790 );
and ( n11795 , n11793 , n11794 );
nor ( n11796 , n11792 , n11795 );
buf ( n11797 , n5125 );
buf ( n11798 , n5126 );
buf ( n11799 , n11798 );
not ( n11800 , n11799 );
buf ( n11801 , n5127 );
nand ( n11802 , n7912 , n11801 );
not ( n11803 , n11802 );
or ( n11804 , n11800 , n11803 );
not ( n11805 , n11798 );
nand ( n11806 , n6927 , n11805 , n11801 );
nand ( n11807 , n11804 , n11806 );
xor ( n11808 , n11797 , n11807 );
buf ( n11809 , n5128 );
nand ( n11810 , n7107 , n11809 );
buf ( n11811 , n5129 );
not ( n11812 , n11811 );
and ( n11813 , n11810 , n11812 );
not ( n11814 , n11810 );
buf ( n11815 , n11811 );
and ( n11816 , n11814 , n11815 );
nor ( n11817 , n11813 , n11816 );
xnor ( n11818 , n11808 , n11817 );
not ( n11819 , n11818 );
xor ( n11820 , n11796 , n11819 );
not ( n11821 , n11060 );
buf ( n11822 , n5130 );
not ( n11823 , n11822 );
not ( n11824 , n11823 );
or ( n11825 , n11821 , n11824 );
not ( n11826 , n11059 );
buf ( n11827 , n11822 );
nand ( n11828 , n11826 , n11827 );
nand ( n11829 , n11825 , n11828 );
buf ( n11830 , n5131 );
not ( n11831 , n11830 );
and ( n11832 , n11829 , n11831 );
not ( n11833 , n11829 );
buf ( n11834 , n11830 );
and ( n11835 , n11833 , n11834 );
nor ( n11836 , n11832 , n11835 );
buf ( n11837 , n5132 );
nand ( n11838 , n6828 , n11837 );
buf ( n11839 , n5133 );
buf ( n11840 , n11839 );
and ( n11841 , n11838 , n11840 );
not ( n11842 , n11838 );
not ( n11843 , n11839 );
and ( n11844 , n11842 , n11843 );
nor ( n11845 , n11841 , n11844 );
xor ( n11846 , n11836 , n11845 );
buf ( n11847 , n8954 );
buf ( n11848 , n5134 );
nand ( n11849 , n11847 , n11848 );
buf ( n11850 , n5135 );
not ( n11851 , n11850 );
and ( n11852 , n11849 , n11851 );
not ( n11853 , n11849 );
buf ( n11854 , n11850 );
and ( n11855 , n11853 , n11854 );
nor ( n11856 , n11852 , n11855 );
xnor ( n11857 , n11846 , n11856 );
not ( n11858 , n11857 );
xnor ( n11859 , n11820 , n11858 );
not ( n11860 , n11859 );
nand ( n11861 , n11778 , n11860 );
buf ( n11862 , n5136 );
buf ( n11863 , n11862 );
not ( n11864 , n11863 );
not ( n11865 , n11226 );
or ( n11866 , n11864 , n11865 );
or ( n11867 , n11226 , n11863 );
nand ( n11868 , n11866 , n11867 );
xor ( n11869 , n11868 , n11271 );
not ( n11870 , n11869 );
and ( n11871 , n11861 , n11870 );
not ( n11872 , n11861 );
and ( n11873 , n11872 , n11869 );
nor ( n11874 , n11871 , n11873 );
not ( n11875 , n11874 );
not ( n11876 , n11875 );
or ( n11877 , n11733 , n11876 );
nand ( n11878 , n11874 , n11731 );
nand ( n11879 , n11877 , n11878 );
buf ( n11880 , n5137 );
nand ( n11881 , n8537 , n11880 );
buf ( n11882 , n5138 );
buf ( n11883 , n11882 );
and ( n11884 , n11881 , n11883 );
not ( n11885 , n11881 );
not ( n11886 , n11882 );
and ( n11887 , n11885 , n11886 );
nor ( n11888 , n11884 , n11887 );
not ( n11889 , n9389 );
buf ( n11890 , n5139 );
not ( n11891 , n11890 );
not ( n11892 , n11891 );
or ( n11893 , n11889 , n11892 );
not ( n11894 , n9388 );
buf ( n11895 , n11890 );
nand ( n11896 , n11894 , n11895 );
nand ( n11897 , n11893 , n11896 );
not ( n11898 , n11897 );
buf ( n11899 , n5140 );
buf ( n11900 , n5141 );
nand ( n11901 , n8069 , n11900 );
not ( n11902 , n11901 );
buf ( n11903 , n5142 );
not ( n11904 , n11903 );
and ( n11905 , n11902 , n11904 );
nand ( n11906 , n7013 , n11900 );
and ( n11907 , n11906 , n11903 );
nor ( n11908 , n11905 , n11907 );
xor ( n11909 , n11899 , n11908 );
xnor ( n11910 , n11909 , n11172 );
not ( n11911 , n11910 );
not ( n11912 , n11911 );
or ( n11913 , n11898 , n11912 );
not ( n11914 , n11897 );
nand ( n11915 , n11910 , n11914 );
nand ( n11916 , n11913 , n11915 );
xor ( n11917 , n11888 , n11916 );
buf ( n11918 , n5143 );
buf ( n11919 , n11918 );
not ( n11920 , n11919 );
buf ( n11921 , n5144 );
not ( n11922 , n11921 );
not ( n11923 , n11922 );
or ( n11924 , n11920 , n11923 );
not ( n11925 , n11918 );
buf ( n11926 , n11921 );
nand ( n11927 , n11925 , n11926 );
nand ( n11928 , n11924 , n11927 );
buf ( n11929 , n5145 );
not ( n11930 , n11929 );
and ( n11931 , n11928 , n11930 );
not ( n11932 , n11928 );
buf ( n11933 , n11929 );
and ( n11934 , n11932 , n11933 );
nor ( n11935 , n11931 , n11934 );
buf ( n11936 , n5146 );
nand ( n11937 , n6770 , n11936 );
buf ( n11938 , n5147 );
buf ( n11939 , n11938 );
and ( n11940 , n11937 , n11939 );
not ( n11941 , n11937 );
not ( n11942 , n11938 );
and ( n11943 , n11941 , n11942 );
nor ( n11944 , n11940 , n11943 );
xor ( n11945 , n11935 , n11944 );
buf ( n11946 , n8454 );
buf ( n11947 , n5148 );
nand ( n11948 , n11946 , n11947 );
buf ( n11949 , n5149 );
not ( n11950 , n11949 );
and ( n11951 , n11948 , n11950 );
not ( n11952 , n11948 );
buf ( n11953 , n11949 );
and ( n11954 , n11952 , n11953 );
nor ( n11955 , n11951 , n11954 );
xnor ( n11956 , n11945 , n11955 );
buf ( n11957 , n11956 );
not ( n11958 , n11957 );
xnor ( n11959 , n11917 , n11958 );
not ( n11960 , n11959 );
buf ( n11961 , n5150 );
nand ( n11962 , n7202 , n11961 );
buf ( n11963 , n5151 );
buf ( n11964 , n11963 );
and ( n11965 , n11962 , n11964 );
not ( n11966 , n11962 );
not ( n11967 , n11963 );
and ( n11968 , n11966 , n11967 );
nor ( n11969 , n11965 , n11968 );
buf ( n11970 , n11969 );
not ( n11971 , n11970 );
not ( n11972 , n11971 );
buf ( n11973 , n5152 );
buf ( n11974 , n11973 );
not ( n11975 , n11974 );
buf ( n11976 , n5153 );
not ( n11977 , n11976 );
not ( n11978 , n11977 );
or ( n11979 , n11975 , n11978 );
not ( n11980 , n11973 );
buf ( n11981 , n11976 );
nand ( n11982 , n11980 , n11981 );
nand ( n11983 , n11979 , n11982 );
buf ( n11984 , n5154 );
buf ( n11985 , n11984 );
and ( n11986 , n11983 , n11985 );
not ( n11987 , n11983 );
not ( n11988 , n11984 );
and ( n11989 , n11987 , n11988 );
nor ( n11990 , n11986 , n11989 );
buf ( n11991 , n5155 );
nand ( n11992 , n7013 , n11991 );
buf ( n11993 , n5156 );
buf ( n11994 , n11993 );
and ( n11995 , n11992 , n11994 );
not ( n11996 , n11992 );
not ( n11997 , n11993 );
and ( n11998 , n11996 , n11997 );
nor ( n11999 , n11995 , n11998 );
xor ( n12000 , n11990 , n11999 );
buf ( n12001 , n5157 );
nand ( n12002 , n8375 , n12001 );
buf ( n12003 , n5158 );
not ( n12004 , n12003 );
and ( n12005 , n12002 , n12004 );
not ( n12006 , n12002 );
buf ( n12007 , n12003 );
and ( n12008 , n12006 , n12007 );
nor ( n12009 , n12005 , n12008 );
xnor ( n12010 , n12000 , n12009 );
buf ( n12011 , n12010 );
not ( n12012 , n12011 );
not ( n12013 , n12012 );
or ( n12014 , n11972 , n12013 );
nand ( n12015 , n12011 , n11970 );
nand ( n12016 , n12014 , n12015 );
not ( n12017 , n12016 );
buf ( n12018 , n5159 );
not ( n12019 , n12018 );
buf ( n12020 , n5160 );
not ( n12021 , n12020 );
buf ( n12022 , n5161 );
buf ( n12023 , n12022 );
nand ( n12024 , n12021 , n12023 );
not ( n12025 , n12022 );
buf ( n12026 , n12020 );
nand ( n12027 , n12025 , n12026 );
and ( n12028 , n12024 , n12027 );
xor ( n12029 , n12019 , n12028 );
buf ( n12030 , n5162 );
buf ( n12031 , n5163 );
buf ( n12032 , n12031 );
xor ( n12033 , n12030 , n12032 );
buf ( n12034 , n5164 );
nand ( n12035 , n6719 , n12034 );
xnor ( n12036 , n12033 , n12035 );
xnor ( n12037 , n12029 , n12036 );
buf ( n12038 , n12037 );
not ( n12039 , n12038 );
and ( n12040 , n12017 , n12039 );
and ( n12041 , n12038 , n12016 );
nor ( n12042 , n12040 , n12041 );
not ( n12043 , n12042 );
nand ( n12044 , n11960 , n12043 );
buf ( n12045 , n5165 );
buf ( n12046 , n12045 );
not ( n12047 , n12046 );
not ( n12048 , n7150 );
buf ( n12049 , n5166 );
not ( n12050 , n12049 );
not ( n12051 , n12050 );
or ( n12052 , n12048 , n12051 );
not ( n12053 , n7149 );
buf ( n12054 , n12049 );
nand ( n12055 , n12053 , n12054 );
nand ( n12056 , n12052 , n12055 );
buf ( n12057 , n5167 );
buf ( n12058 , n12057 );
and ( n12059 , n12056 , n12058 );
not ( n12060 , n12056 );
not ( n12061 , n12057 );
and ( n12062 , n12060 , n12061 );
nor ( n12063 , n12059 , n12062 );
buf ( n12064 , n5168 );
nand ( n12065 , n7014 , n12064 );
buf ( n12066 , n5169 );
not ( n12067 , n12066 );
and ( n12068 , n12065 , n12067 );
not ( n12069 , n12065 );
buf ( n12070 , n12066 );
and ( n12071 , n12069 , n12070 );
nor ( n12072 , n12068 , n12071 );
xor ( n12073 , n12063 , n12072 );
buf ( n12074 , n5170 );
nand ( n12075 , n8223 , n12074 );
buf ( n12076 , n5171 );
not ( n12077 , n12076 );
and ( n12078 , n12075 , n12077 );
not ( n12079 , n12075 );
buf ( n12080 , n12076 );
and ( n12081 , n12079 , n12080 );
nor ( n12082 , n12078 , n12081 );
xnor ( n12083 , n12073 , n12082 );
not ( n12084 , n12083 );
or ( n12085 , n12047 , n12084 );
not ( n12086 , n12083 );
not ( n12087 , n12086 );
or ( n12088 , n12087 , n12046 );
nand ( n12089 , n12085 , n12088 );
buf ( n12090 , n5172 );
buf ( n12091 , n12090 );
not ( n12092 , n12091 );
buf ( n12093 , n5173 );
not ( n12094 , n12093 );
not ( n12095 , n12094 );
or ( n12096 , n12092 , n12095 );
not ( n12097 , n12090 );
buf ( n12098 , n12093 );
nand ( n12099 , n12097 , n12098 );
nand ( n12100 , n12096 , n12099 );
buf ( n12101 , n5174 );
buf ( n12102 , n12101 );
and ( n12103 , n12100 , n12102 );
not ( n12104 , n12100 );
not ( n12105 , n12101 );
and ( n12106 , n12104 , n12105 );
nor ( n12107 , n12103 , n12106 );
buf ( n12108 , n5175 );
nand ( n12109 , n6502 , n12108 );
buf ( n12110 , n5176 );
buf ( n12111 , n12110 );
and ( n12112 , n12109 , n12111 );
not ( n12113 , n12109 );
not ( n12114 , n12110 );
and ( n12115 , n12113 , n12114 );
nor ( n12116 , n12112 , n12115 );
xor ( n12117 , n12107 , n12116 );
buf ( n12118 , n5177 );
nand ( n12119 , n8675 , n12118 );
buf ( n12120 , n5178 );
not ( n12121 , n12120 );
and ( n12122 , n12119 , n12121 );
not ( n12123 , n12119 );
buf ( n12124 , n12120 );
and ( n12125 , n12123 , n12124 );
nor ( n12126 , n12122 , n12125 );
xor ( n12127 , n12117 , n12126 );
buf ( n12128 , n12127 );
and ( n12129 , n12089 , n12128 );
not ( n12130 , n12089 );
not ( n12131 , n12128 );
and ( n12132 , n12130 , n12131 );
nor ( n12133 , n12129 , n12132 );
and ( n12134 , n12044 , n12133 );
not ( n12135 , n12044 );
not ( n12136 , n12133 );
and ( n12137 , n12135 , n12136 );
nor ( n12138 , n12134 , n12137 );
and ( n12139 , n11879 , n12138 );
not ( n12140 , n11879 );
not ( n12141 , n12138 );
and ( n12142 , n12140 , n12141 );
nor ( n12143 , n12139 , n12142 );
not ( n12144 , n12143 );
not ( n12145 , n12144 );
not ( n12146 , n11443 );
nand ( n12147 , n11512 , n12146 );
not ( n12148 , n12147 );
not ( n12149 , n11154 );
xor ( n12150 , n10369 , n12149 );
xor ( n12151 , n12150 , n7833 );
not ( n12152 , n12151 );
not ( n12153 , n12152 );
or ( n12154 , n12148 , n12153 );
or ( n12155 , n12152 , n12147 );
nand ( n12156 , n12154 , n12155 );
not ( n12157 , n12156 );
not ( n12158 , n12157 );
buf ( n12159 , n5179 );
nand ( n12160 , n6927 , n12159 );
buf ( n12161 , n5180 );
buf ( n12162 , n12161 );
and ( n12163 , n12160 , n12162 );
not ( n12164 , n12160 );
not ( n12165 , n12161 );
and ( n12166 , n12164 , n12165 );
nor ( n12167 , n12163 , n12166 );
buf ( n12168 , n5181 );
buf ( n12169 , n12168 );
not ( n12170 , n12169 );
buf ( n12171 , n5182 );
not ( n12172 , n12171 );
not ( n12173 , n12172 );
or ( n12174 , n12170 , n12173 );
not ( n12175 , n12168 );
buf ( n12176 , n12171 );
nand ( n12177 , n12175 , n12176 );
nand ( n12178 , n12174 , n12177 );
buf ( n12179 , n5183 );
buf ( n12180 , n12179 );
and ( n12181 , n12178 , n12180 );
not ( n12182 , n12178 );
not ( n12183 , n12179 );
and ( n12184 , n12182 , n12183 );
nor ( n12185 , n12181 , n12184 );
not ( n12186 , n12185 );
buf ( n12187 , n5184 );
nand ( n12188 , n6646 , n12187 );
buf ( n12189 , n5185 );
buf ( n12190 , n12189 );
and ( n12191 , n12188 , n12190 );
not ( n12192 , n12188 );
not ( n12193 , n12189 );
and ( n12194 , n12192 , n12193 );
nor ( n12195 , n12191 , n12194 );
xor ( n12196 , n12186 , n12195 );
buf ( n12197 , n5186 );
nand ( n12198 , n6816 , n12197 );
buf ( n12199 , n5187 );
not ( n12200 , n12199 );
and ( n12201 , n12198 , n12200 );
not ( n12202 , n12198 );
buf ( n12203 , n12199 );
and ( n12204 , n12202 , n12203 );
nor ( n12205 , n12201 , n12204 );
xnor ( n12206 , n12196 , n12205 );
xor ( n12207 , n12167 , n12206 );
buf ( n12208 , n5188 );
not ( n12209 , n12208 );
buf ( n12210 , n5189 );
buf ( n12211 , n12210 );
and ( n12212 , n12209 , n12211 );
not ( n12213 , n12209 );
not ( n12214 , n12210 );
and ( n12215 , n12213 , n12214 );
nor ( n12216 , n12212 , n12215 );
not ( n12217 , n12216 );
buf ( n12218 , n5190 );
buf ( n12219 , n5191 );
not ( n12220 , n12219 );
xor ( n12221 , n12218 , n12220 );
buf ( n12222 , n5192 );
nand ( n12223 , n6816 , n12222 );
buf ( n12224 , n5193 );
not ( n12225 , n12224 );
and ( n12226 , n12223 , n12225 );
not ( n12227 , n12223 );
buf ( n12228 , n12224 );
and ( n12229 , n12227 , n12228 );
nor ( n12230 , n12226 , n12229 );
xnor ( n12231 , n12221 , n12230 );
not ( n12232 , n12231 );
or ( n12233 , n12217 , n12232 );
or ( n12234 , n12231 , n12216 );
nand ( n12235 , n12233 , n12234 );
buf ( n12236 , n12235 );
xnor ( n12237 , n12207 , n12236 );
not ( n12238 , n12237 );
buf ( n12239 , n5194 );
not ( n12240 , n12239 );
buf ( n12241 , n5195 );
nand ( n12242 , n7569 , n12241 );
not ( n12243 , n12242 );
or ( n12244 , n12240 , n12243 );
or ( n12245 , n12242 , n12239 );
nand ( n12246 , n12244 , n12245 );
not ( n12247 , n12246 );
buf ( n12248 , n5196 );
buf ( n12249 , n12248 );
not ( n12250 , n12249 );
buf ( n12251 , n5197 );
not ( n12252 , n12251 );
not ( n12253 , n12252 );
or ( n12254 , n12250 , n12253 );
not ( n12255 , n12248 );
buf ( n12256 , n12251 );
nand ( n12257 , n12255 , n12256 );
nand ( n12258 , n12254 , n12257 );
buf ( n12259 , n5198 );
not ( n12260 , n12259 );
and ( n12261 , n12258 , n12260 );
not ( n12262 , n12258 );
buf ( n12263 , n12259 );
and ( n12264 , n12262 , n12263 );
nor ( n12265 , n12261 , n12264 );
buf ( n12266 , n5199 );
nand ( n12267 , n7107 , n12266 );
buf ( n12268 , n5200 );
buf ( n12269 , n12268 );
and ( n12270 , n12267 , n12269 );
not ( n12271 , n12267 );
not ( n12272 , n12268 );
and ( n12273 , n12271 , n12272 );
nor ( n12274 , n12270 , n12273 );
xor ( n12275 , n12265 , n12274 );
buf ( n12276 , n5201 );
nand ( n12277 , n7107 , n12276 );
buf ( n12278 , n5202 );
buf ( n12279 , n12278 );
and ( n12280 , n12277 , n12279 );
not ( n12281 , n12277 );
not ( n12282 , n12278 );
and ( n12283 , n12281 , n12282 );
nor ( n12284 , n12280 , n12283 );
not ( n12285 , n12284 );
xnor ( n12286 , n12275 , n12285 );
buf ( n12287 , n12286 );
not ( n12288 , n12287 );
or ( n12289 , n12247 , n12288 );
or ( n12290 , n12246 , n12286 );
nand ( n12291 , n12289 , n12290 );
not ( n12292 , n8619 );
and ( n12293 , n12291 , n12292 );
not ( n12294 , n12291 );
and ( n12295 , n12294 , n8620 );
nor ( n12296 , n12293 , n12295 );
not ( n12297 , n12296 );
nand ( n12298 , n12238 , n12297 );
not ( n12299 , n12298 );
buf ( n12300 , n5203 );
buf ( n12301 , n12300 );
not ( n12302 , n12301 );
buf ( n12303 , n5204 );
buf ( n12304 , n12303 );
not ( n12305 , n12304 );
buf ( n12306 , n5205 );
not ( n12307 , n12306 );
not ( n12308 , n12307 );
or ( n12309 , n12305 , n12308 );
not ( n12310 , n12303 );
buf ( n12311 , n12306 );
nand ( n12312 , n12310 , n12311 );
nand ( n12313 , n12309 , n12312 );
buf ( n12314 , n5206 );
not ( n12315 , n12314 );
and ( n12316 , n12313 , n12315 );
not ( n12317 , n12313 );
buf ( n12318 , n12314 );
and ( n12319 , n12317 , n12318 );
nor ( n12320 , n12316 , n12319 );
buf ( n12321 , n5207 );
nand ( n12322 , n8176 , n12321 );
buf ( n12323 , n5208 );
buf ( n12324 , n12323 );
and ( n12325 , n12322 , n12324 );
not ( n12326 , n12322 );
not ( n12327 , n12323 );
and ( n12328 , n12326 , n12327 );
nor ( n12329 , n12325 , n12328 );
xor ( n12330 , n12320 , n12329 );
buf ( n12331 , n5209 );
nand ( n12332 , n6916 , n12331 );
buf ( n12333 , n5210 );
buf ( n12334 , n12333 );
and ( n12335 , n12332 , n12334 );
not ( n12336 , n12332 );
not ( n12337 , n12333 );
and ( n12338 , n12336 , n12337 );
nor ( n12339 , n12335 , n12338 );
not ( n12340 , n12339 );
xnor ( n12341 , n12330 , n12340 );
buf ( n12342 , n12341 );
not ( n12343 , n12342 );
or ( n12344 , n12302 , n12343 );
or ( n12345 , n12342 , n12301 );
nand ( n12346 , n12344 , n12345 );
not ( n12347 , n12346 );
buf ( n12348 , n5211 );
not ( n12349 , n12348 );
buf ( n12350 , n5212 );
buf ( n12351 , n12350 );
not ( n12352 , n12351 );
not ( n12353 , n10537 );
not ( n12354 , n12353 );
or ( n12355 , n12352 , n12354 );
not ( n12356 , n12350 );
nand ( n12357 , n12356 , n10538 );
nand ( n12358 , n12355 , n12357 );
xor ( n12359 , n12349 , n12358 );
buf ( n12360 , n5213 );
nand ( n12361 , n8176 , n12360 );
buf ( n12362 , n5214 );
buf ( n12363 , n12362 );
and ( n12364 , n12361 , n12363 );
not ( n12365 , n12361 );
not ( n12366 , n12362 );
and ( n12367 , n12365 , n12366 );
nor ( n12368 , n12364 , n12367 );
not ( n12369 , n12368 );
buf ( n12370 , n5215 );
not ( n12371 , n12370 );
and ( n12372 , n12369 , n12371 );
and ( n12373 , n12368 , n12370 );
nor ( n12374 , n12372 , n12373 );
xor ( n12375 , n12359 , n12374 );
not ( n12376 , n12375 );
not ( n12377 , n12376 );
and ( n12378 , n12347 , n12377 );
buf ( n12379 , n12376 );
and ( n12380 , n12346 , n12379 );
nor ( n12381 , n12378 , n12380 );
not ( n12382 , n12381 );
not ( n12383 , n12382 );
and ( n12384 , n12299 , n12383 );
and ( n12385 , n12298 , n12382 );
nor ( n12386 , n12384 , n12385 );
not ( n12387 , n12386 );
not ( n12388 , n12387 );
or ( n12389 , n12158 , n12388 );
nand ( n12390 , n12386 , n12156 );
nand ( n12391 , n12389 , n12390 );
not ( n12392 , n12391 );
and ( n12393 , n12145 , n12392 );
and ( n12394 , n12144 , n12391 );
nor ( n12395 , n12393 , n12394 );
not ( n12396 , n12395 );
or ( n12397 , n11519 , n12396 );
not ( n12398 , n11518 );
and ( n12399 , n12143 , n12391 );
not ( n12400 , n12143 );
not ( n12401 , n12391 );
and ( n12402 , n12400 , n12401 );
nor ( n12403 , n12399 , n12402 );
nand ( n12404 , n12398 , n12403 );
nand ( n12405 , n12397 , n12404 );
buf ( n12406 , n5216 );
buf ( n12407 , n12406 );
not ( n12408 , n12407 );
buf ( n12409 , n5217 );
buf ( n12410 , n12409 );
not ( n12411 , n12410 );
buf ( n12412 , n5218 );
not ( n12413 , n12412 );
not ( n12414 , n12413 );
or ( n12415 , n12411 , n12414 );
not ( n12416 , n12409 );
buf ( n12417 , n12412 );
nand ( n12418 , n12416 , n12417 );
nand ( n12419 , n12415 , n12418 );
buf ( n12420 , n5219 );
buf ( n12421 , n12420 );
and ( n12422 , n12419 , n12421 );
not ( n12423 , n12419 );
not ( n12424 , n12420 );
and ( n12425 , n12423 , n12424 );
nor ( n12426 , n12422 , n12425 );
buf ( n12427 , n5220 );
nand ( n12428 , n8364 , n12427 );
buf ( n12429 , n5221 );
xor ( n12430 , n12428 , n12429 );
xor ( n12431 , n12426 , n12430 );
buf ( n12432 , n5222 );
nand ( n12433 , n9310 , n12432 );
buf ( n12434 , n5223 );
not ( n12435 , n12434 );
and ( n12436 , n12433 , n12435 );
not ( n12437 , n12433 );
buf ( n12438 , n12434 );
and ( n12439 , n12437 , n12438 );
nor ( n12440 , n12436 , n12439 );
xor ( n12441 , n12431 , n12440 );
buf ( n12442 , n12441 );
not ( n12443 , n12442 );
or ( n12444 , n12408 , n12443 );
or ( n12445 , n12442 , n12407 );
nand ( n12446 , n12444 , n12445 );
not ( n12447 , n12446 );
buf ( n12448 , n5224 );
buf ( n12449 , n5225 );
not ( n12450 , n12449 );
buf ( n12451 , n5226 );
buf ( n12452 , n12451 );
and ( n12453 , n12450 , n12452 );
not ( n12454 , n12450 );
not ( n12455 , n12451 );
and ( n12456 , n12454 , n12455 );
nor ( n12457 , n12453 , n12456 );
xor ( n12458 , n12448 , n12457 );
buf ( n12459 , n5227 );
xor ( n12460 , n12459 , n12239 );
xnor ( n12461 , n12460 , n12242 );
xnor ( n12462 , n12458 , n12461 );
not ( n12463 , n12462 );
not ( n12464 , n12463 );
and ( n12465 , n12447 , n12464 );
not ( n12466 , n12462 );
and ( n12467 , n12446 , n12466 );
nor ( n12468 , n12465 , n12467 );
buf ( n12469 , n5228 );
buf ( n12470 , n12469 );
not ( n12471 , n12470 );
buf ( n12472 , n5229 );
buf ( n12473 , n12472 );
not ( n12474 , n12473 );
buf ( n12475 , n5230 );
not ( n12476 , n12475 );
not ( n12477 , n12476 );
or ( n12478 , n12474 , n12477 );
not ( n12479 , n12472 );
buf ( n12480 , n12475 );
nand ( n12481 , n12479 , n12480 );
nand ( n12482 , n12478 , n12481 );
and ( n12483 , n12482 , n10093 );
not ( n12484 , n12482 );
and ( n12485 , n12484 , n10049 );
nor ( n12486 , n12483 , n12485 );
xor ( n12487 , n12486 , n10483 );
buf ( n12488 , n5231 );
nand ( n12489 , n6558 , n12488 );
buf ( n12490 , n5232 );
not ( n12491 , n12490 );
and ( n12492 , n12489 , n12491 );
not ( n12493 , n12489 );
buf ( n12494 , n12490 );
and ( n12495 , n12493 , n12494 );
nor ( n12496 , n12492 , n12495 );
xnor ( n12497 , n12487 , n12496 );
buf ( n12498 , n12497 );
not ( n12499 , n12498 );
or ( n12500 , n12471 , n12499 );
or ( n12501 , n12498 , n12470 );
nand ( n12502 , n12500 , n12501 );
not ( n12503 , n12502 );
buf ( n12504 , n5233 );
buf ( n12505 , n12504 );
not ( n12506 , n12505 );
buf ( n12507 , n5234 );
not ( n12508 , n12507 );
not ( n12509 , n12508 );
or ( n12510 , n12506 , n12509 );
not ( n12511 , n12504 );
buf ( n12512 , n12507 );
nand ( n12513 , n12511 , n12512 );
nand ( n12514 , n12510 , n12513 );
buf ( n12515 , n5235 );
not ( n12516 , n12515 );
and ( n12517 , n12514 , n12516 );
not ( n12518 , n12514 );
buf ( n12519 , n12515 );
and ( n12520 , n12518 , n12519 );
nor ( n12521 , n12517 , n12520 );
buf ( n12522 , n5236 );
nand ( n12523 , n6770 , n12522 );
buf ( n12524 , n5237 );
buf ( n12525 , n12524 );
and ( n12526 , n12523 , n12525 );
not ( n12527 , n12523 );
not ( n12528 , n12524 );
and ( n12529 , n12527 , n12528 );
nor ( n12530 , n12526 , n12529 );
xor ( n12531 , n12521 , n12530 );
buf ( n12532 , n5238 );
nand ( n12533 , n6719 , n12532 );
buf ( n12534 , n5239 );
not ( n12535 , n12534 );
and ( n12536 , n12533 , n12535 );
not ( n12537 , n12533 );
buf ( n12538 , n12534 );
and ( n12539 , n12537 , n12538 );
nor ( n12540 , n12536 , n12539 );
xor ( n12541 , n12531 , n12540 );
not ( n12542 , n12541 );
buf ( n12543 , n12542 );
not ( n12544 , n12543 );
and ( n12545 , n12503 , n12544 );
buf ( n12546 , n12542 );
and ( n12547 , n12502 , n12546 );
nor ( n12548 , n12545 , n12547 );
not ( n12549 , n12548 );
nand ( n12550 , n12468 , n12549 );
not ( n12551 , n12550 );
not ( n12552 , n6790 );
not ( n12553 , n12552 );
buf ( n12554 , n5240 );
buf ( n12555 , n12554 );
not ( n12556 , n12555 );
buf ( n12557 , n5241 );
not ( n12558 , n12557 );
not ( n12559 , n12558 );
or ( n12560 , n12556 , n12559 );
not ( n12561 , n12554 );
buf ( n12562 , n12557 );
nand ( n12563 , n12561 , n12562 );
nand ( n12564 , n12560 , n12563 );
buf ( n12565 , n5242 );
not ( n12566 , n12565 );
and ( n12567 , n12564 , n12566 );
not ( n12568 , n12564 );
buf ( n12569 , n12565 );
and ( n12570 , n12568 , n12569 );
nor ( n12571 , n12567 , n12570 );
buf ( n12572 , n5243 );
nand ( n12573 , n7912 , n12572 );
buf ( n12574 , n5244 );
buf ( n12575 , n12574 );
and ( n12576 , n12573 , n12575 );
not ( n12577 , n12573 );
not ( n12578 , n12574 );
and ( n12579 , n12577 , n12578 );
nor ( n12580 , n12576 , n12579 );
xor ( n12581 , n12571 , n12580 );
buf ( n12582 , n5245 );
nand ( n12583 , n7912 , n12582 );
buf ( n12584 , n5246 );
buf ( n12585 , n12584 );
and ( n12586 , n12583 , n12585 );
not ( n12587 , n12583 );
not ( n12588 , n12584 );
and ( n12589 , n12587 , n12588 );
nor ( n12590 , n12586 , n12589 );
xnor ( n12591 , n12581 , n12590 );
not ( n12592 , n12591 );
or ( n12593 , n12553 , n12592 );
not ( n12594 , n12591 );
not ( n12595 , n12594 );
or ( n12596 , n12595 , n12552 );
nand ( n12597 , n12593 , n12596 );
buf ( n12598 , n5247 );
buf ( n12599 , n12598 );
not ( n12600 , n12599 );
buf ( n12601 , n5248 );
not ( n12602 , n12601 );
not ( n12603 , n12602 );
or ( n12604 , n12600 , n12603 );
not ( n12605 , n12598 );
buf ( n12606 , n12601 );
nand ( n12607 , n12605 , n12606 );
nand ( n12608 , n12604 , n12607 );
buf ( n12609 , n5249 );
buf ( n12610 , n12609 );
and ( n12611 , n12608 , n12610 );
not ( n12612 , n12608 );
not ( n12613 , n12609 );
and ( n12614 , n12612 , n12613 );
nor ( n12615 , n12611 , n12614 );
buf ( n12616 , n5250 );
nand ( n12617 , n7293 , n12616 );
buf ( n12618 , n5251 );
buf ( n12619 , n12618 );
and ( n12620 , n12617 , n12619 );
not ( n12621 , n12617 );
not ( n12622 , n12618 );
and ( n12623 , n12621 , n12622 );
nor ( n12624 , n12620 , n12623 );
xor ( n12625 , n12615 , n12624 );
buf ( n12626 , n5252 );
nand ( n12627 , n11946 , n12626 );
buf ( n12628 , n5253 );
buf ( n12629 , n12628 );
and ( n12630 , n12627 , n12629 );
not ( n12631 , n12627 );
not ( n12632 , n12628 );
and ( n12633 , n12631 , n12632 );
nor ( n12634 , n12630 , n12633 );
xnor ( n12635 , n12625 , n12634 );
buf ( n12636 , n12635 );
buf ( n12637 , n12636 );
not ( n12638 , n12637 );
and ( n12639 , n12597 , n12638 );
not ( n12640 , n12597 );
and ( n12641 , n12640 , n12637 );
nor ( n12642 , n12639 , n12641 );
not ( n12643 , n12642 );
and ( n12644 , n12551 , n12643 );
and ( n12645 , n12550 , n12642 );
nor ( n12646 , n12644 , n12645 );
not ( n12647 , n12646 );
not ( n12648 , n12647 );
xor ( n12649 , n10646 , n10665 );
not ( n12650 , n10655 );
xnor ( n12651 , n12649 , n12650 );
not ( n12652 , n12651 );
buf ( n12653 , n5254 );
buf ( n12654 , n12653 );
not ( n12655 , n12654 );
and ( n12656 , n12652 , n12655 );
and ( n12657 , n12651 , n12654 );
nor ( n12658 , n12656 , n12657 );
and ( n12659 , n12658 , n10679 );
not ( n12660 , n12658 );
and ( n12661 , n12660 , n10678 );
nor ( n12662 , n12659 , n12661 );
buf ( n12663 , n5255 );
buf ( n12664 , n12663 );
not ( n12665 , n12664 );
buf ( n12666 , n5256 );
nand ( n12667 , n6770 , n12666 );
buf ( n12668 , n5257 );
buf ( n12669 , n12668 );
and ( n12670 , n12667 , n12669 );
not ( n12671 , n12667 );
not ( n12672 , n12668 );
and ( n12673 , n12671 , n12672 );
nor ( n12674 , n12670 , n12673 );
not ( n12675 , n12674 );
buf ( n12676 , n5258 );
nand ( n12677 , n7868 , n12676 );
buf ( n12678 , n5259 );
not ( n12679 , n12678 );
and ( n12680 , n12677 , n12679 );
not ( n12681 , n12677 );
buf ( n12682 , n12678 );
and ( n12683 , n12681 , n12682 );
nor ( n12684 , n12680 , n12683 );
not ( n12685 , n12684 );
or ( n12686 , n12675 , n12685 );
or ( n12687 , n12674 , n12684 );
nand ( n12688 , n12686 , n12687 );
buf ( n12689 , n5260 );
buf ( n12690 , n12689 );
not ( n12691 , n12690 );
buf ( n12692 , n5261 );
not ( n12693 , n12692 );
not ( n12694 , n12693 );
or ( n12695 , n12691 , n12694 );
not ( n12696 , n12689 );
buf ( n12697 , n12692 );
nand ( n12698 , n12696 , n12697 );
nand ( n12699 , n12695 , n12698 );
buf ( n12700 , n5262 );
buf ( n12701 , n12700 );
and ( n12702 , n12699 , n12701 );
not ( n12703 , n12699 );
not ( n12704 , n12700 );
and ( n12705 , n12703 , n12704 );
nor ( n12706 , n12702 , n12705 );
xnor ( n12707 , n12688 , n12706 );
not ( n12708 , n12707 );
or ( n12709 , n12665 , n12708 );
not ( n12710 , n12664 );
xor ( n12711 , n12706 , n12674 );
buf ( n12712 , n12684 );
xnor ( n12713 , n12711 , n12712 );
nand ( n12714 , n12710 , n12713 );
nand ( n12715 , n12709 , n12714 );
not ( n12716 , n12715 );
buf ( n12717 , n5263 );
buf ( n12718 , n12717 );
not ( n12719 , n12718 );
buf ( n12720 , n5264 );
not ( n12721 , n12720 );
not ( n12722 , n12721 );
or ( n12723 , n12719 , n12722 );
not ( n12724 , n12717 );
buf ( n12725 , n12720 );
nand ( n12726 , n12724 , n12725 );
nand ( n12727 , n12723 , n12726 );
buf ( n12728 , n5265 );
not ( n12729 , n12728 );
and ( n12730 , n12727 , n12729 );
not ( n12731 , n12727 );
buf ( n12732 , n12728 );
and ( n12733 , n12731 , n12732 );
nor ( n12734 , n12730 , n12733 );
buf ( n12735 , n5266 );
nand ( n12736 , n7977 , n12735 );
buf ( n12737 , n5267 );
buf ( n12738 , n12737 );
and ( n12739 , n12736 , n12738 );
not ( n12740 , n12736 );
not ( n12741 , n12737 );
and ( n12742 , n12740 , n12741 );
nor ( n12743 , n12739 , n12742 );
xor ( n12744 , n12734 , n12743 );
buf ( n12745 , n5268 );
nand ( n12746 , n11946 , n12745 );
buf ( n12747 , n5269 );
not ( n12748 , n12747 );
and ( n12749 , n12746 , n12748 );
not ( n12750 , n12746 );
buf ( n12751 , n12747 );
and ( n12752 , n12750 , n12751 );
nor ( n12753 , n12749 , n12752 );
xnor ( n12754 , n12744 , n12753 );
buf ( n12755 , n12754 );
buf ( n12756 , n12755 );
not ( n12757 , n12756 );
and ( n12758 , n12716 , n12757 );
and ( n12759 , n12715 , n12755 );
nor ( n12760 , n12758 , n12759 );
nand ( n12761 , n12662 , n12760 );
not ( n12762 , n12761 );
buf ( n12763 , n5270 );
nand ( n12764 , n11337 , n12763 );
buf ( n12765 , n5271 );
not ( n12766 , n12765 );
and ( n12767 , n12764 , n12766 );
not ( n12768 , n12764 );
buf ( n12769 , n12765 );
and ( n12770 , n12768 , n12769 );
nor ( n12771 , n12767 , n12770 );
buf ( n12772 , n5272 );
buf ( n12773 , n12772 );
not ( n12774 , n12773 );
buf ( n12775 , n5273 );
not ( n12776 , n12775 );
not ( n12777 , n12776 );
or ( n12778 , n12774 , n12777 );
not ( n12779 , n12772 );
buf ( n12780 , n12775 );
nand ( n12781 , n12779 , n12780 );
nand ( n12782 , n12778 , n12781 );
buf ( n12783 , n5274 );
not ( n12784 , n12783 );
and ( n12785 , n12782 , n12784 );
not ( n12786 , n12782 );
buf ( n12787 , n12783 );
and ( n12788 , n12786 , n12787 );
nor ( n12789 , n12785 , n12788 );
buf ( n12790 , n5275 );
nand ( n12791 , n8954 , n12790 );
buf ( n12792 , n5276 );
buf ( n12793 , n12792 );
and ( n12794 , n12791 , n12793 );
not ( n12795 , n12791 );
not ( n12796 , n12792 );
and ( n12797 , n12795 , n12796 );
nor ( n12798 , n12794 , n12797 );
xor ( n12799 , n12789 , n12798 );
buf ( n12800 , n5277 );
nand ( n12801 , n6871 , n12800 );
buf ( n12802 , n5278 );
buf ( n12803 , n12802 );
and ( n12804 , n12801 , n12803 );
not ( n12805 , n12801 );
not ( n12806 , n12802 );
and ( n12807 , n12805 , n12806 );
nor ( n12808 , n12804 , n12807 );
xor ( n12809 , n12799 , n12808 );
not ( n12810 , n12809 );
buf ( n12811 , n12810 );
xor ( n12812 , n12771 , n12811 );
buf ( n12813 , n5279 );
buf ( n12814 , n12813 );
buf ( n12815 , n5280 );
buf ( n12816 , n12815 );
not ( n12817 , n12816 );
buf ( n12818 , n5281 );
not ( n12819 , n12818 );
not ( n12820 , n12819 );
or ( n12821 , n12817 , n12820 );
not ( n12822 , n12815 );
buf ( n12823 , n12818 );
nand ( n12824 , n12822 , n12823 );
nand ( n12825 , n12821 , n12824 );
xor ( n12826 , n12814 , n12825 );
buf ( n12827 , n5282 );
xor ( n12828 , n9280 , n12827 );
buf ( n12829 , n5283 );
nand ( n12830 , n10874 , n12829 );
xnor ( n12831 , n12828 , n12830 );
xnor ( n12832 , n12826 , n12831 );
buf ( n12833 , n12832 );
xnor ( n12834 , n12812 , n12833 );
not ( n12835 , n12834 );
or ( n12836 , n12762 , n12835 );
or ( n12837 , n12834 , n12761 );
nand ( n12838 , n12836 , n12837 );
not ( n12839 , n12838 );
not ( n12840 , n12839 );
or ( n12841 , n12648 , n12840 );
nand ( n12842 , n12838 , n12646 );
nand ( n12843 , n12841 , n12842 );
buf ( n12844 , n5284 );
buf ( n12845 , n5285 );
buf ( n12846 , n12845 );
not ( n12847 , n12846 );
buf ( n12848 , n5286 );
not ( n12849 , n12848 );
not ( n12850 , n12849 );
or ( n12851 , n12847 , n12850 );
not ( n12852 , n12845 );
buf ( n12853 , n12848 );
nand ( n12854 , n12852 , n12853 );
nand ( n12855 , n12851 , n12854 );
xor ( n12856 , n12844 , n12855 );
buf ( n12857 , n5287 );
buf ( n12858 , n5288 );
not ( n12859 , n12858 );
xor ( n12860 , n12857 , n12859 );
buf ( n12861 , n5289 );
nand ( n12862 , n8260 , n12861 );
xnor ( n12863 , n12860 , n12862 );
xnor ( n12864 , n12856 , n12863 );
buf ( n12865 , n12864 );
not ( n12866 , n12865 );
buf ( n12867 , n5290 );
buf ( n12868 , n12867 );
not ( n12869 , n12868 );
buf ( n12870 , n5291 );
not ( n12871 , n12870 );
not ( n12872 , n12871 );
or ( n12873 , n12869 , n12872 );
not ( n12874 , n12867 );
buf ( n12875 , n12870 );
nand ( n12876 , n12874 , n12875 );
nand ( n12877 , n12873 , n12876 );
and ( n12878 , n12877 , n6943 );
not ( n12879 , n12877 );
and ( n12880 , n12879 , n6896 );
nor ( n12881 , n12878 , n12880 );
buf ( n12882 , n5292 );
nand ( n12883 , n8322 , n12882 );
buf ( n12884 , n5293 );
buf ( n12885 , n12884 );
and ( n12886 , n12883 , n12885 );
not ( n12887 , n12883 );
not ( n12888 , n12884 );
and ( n12889 , n12887 , n12888 );
nor ( n12890 , n12886 , n12889 );
xor ( n12891 , n12881 , n12890 );
buf ( n12892 , n5294 );
nand ( n12893 , n8454 , n12892 );
buf ( n12894 , n5295 );
not ( n12895 , n12894 );
xor ( n12896 , n12893 , n12895 );
xnor ( n12897 , n12891 , n12896 );
buf ( n12898 , n5296 );
buf ( n12899 , n12898 );
nand ( n12900 , n12897 , n12899 );
not ( n12901 , n12900 );
nor ( n12902 , n12897 , n12899 );
nor ( n12903 , n12901 , n12902 );
not ( n12904 , n12903 );
or ( n12905 , n12866 , n12904 );
not ( n12906 , n12864 );
not ( n12907 , n12906 );
or ( n12908 , n12907 , n12903 );
nand ( n12909 , n12905 , n12908 );
not ( n12910 , n7477 );
buf ( n12911 , n5297 );
not ( n12912 , n12911 );
nand ( n12913 , n7489 , n12912 );
not ( n12914 , n12913 );
nor ( n12915 , n7489 , n12912 );
nor ( n12916 , n12914 , n12915 );
not ( n12917 , n12916 );
and ( n12918 , n12910 , n12917 );
and ( n12919 , n7477 , n12916 );
nor ( n12920 , n12918 , n12919 );
not ( n12921 , n12920 );
not ( n12922 , n10916 );
and ( n12923 , n12921 , n12922 );
and ( n12924 , n12920 , n10916 );
nor ( n12925 , n12923 , n12924 );
nand ( n12926 , n12909 , n12925 );
not ( n12927 , n9044 );
not ( n12928 , n10226 );
or ( n12929 , n12927 , n12928 );
not ( n12930 , n9044 );
buf ( n12931 , n10189 );
xor ( n12932 , n10221 , n12931 );
xnor ( n12933 , n12932 , n10199 );
nand ( n12934 , n12930 , n12933 );
nand ( n12935 , n12929 , n12934 );
not ( n12936 , n6734 );
and ( n12937 , n12935 , n12936 );
not ( n12938 , n12935 );
not ( n12939 , n6731 );
and ( n12940 , n12938 , n12939 );
nor ( n12941 , n12937 , n12940 );
and ( n12942 , n12926 , n12941 );
not ( n12943 , n12926 );
not ( n12944 , n12941 );
and ( n12945 , n12943 , n12944 );
nor ( n12946 , n12942 , n12945 );
not ( n12947 , n12946 );
not ( n12948 , n12947 );
not ( n12949 , n10957 );
buf ( n12950 , n5298 );
buf ( n12951 , n12950 );
not ( n12952 , n12951 );
and ( n12953 , n12949 , n12952 );
and ( n12954 , n10957 , n12951 );
nor ( n12955 , n12953 , n12954 );
buf ( n12956 , n5299 );
buf ( n12957 , n12956 );
not ( n12958 , n12957 );
buf ( n12959 , n5300 );
not ( n12960 , n12959 );
not ( n12961 , n12960 );
or ( n12962 , n12958 , n12961 );
not ( n12963 , n12956 );
buf ( n12964 , n12959 );
nand ( n12965 , n12963 , n12964 );
nand ( n12966 , n12962 , n12965 );
buf ( n12967 , n5301 );
not ( n12968 , n12967 );
and ( n12969 , n12966 , n12968 );
not ( n12970 , n12966 );
buf ( n12971 , n12967 );
and ( n12972 , n12970 , n12971 );
nor ( n12973 , n12969 , n12972 );
buf ( n12974 , n5302 );
nand ( n12975 , n6646 , n12974 );
buf ( n12976 , n5303 );
buf ( n12977 , n12976 );
and ( n12978 , n12975 , n12977 );
not ( n12979 , n12975 );
not ( n12980 , n12976 );
and ( n12981 , n12979 , n12980 );
nor ( n12982 , n12978 , n12981 );
xor ( n12983 , n12973 , n12982 );
buf ( n12984 , n5304 );
nand ( n12985 , n6927 , n12984 );
buf ( n12986 , n5305 );
not ( n12987 , n12986 );
and ( n12988 , n12985 , n12987 );
not ( n12989 , n12985 );
buf ( n12990 , n12986 );
and ( n12991 , n12989 , n12990 );
nor ( n12992 , n12988 , n12991 );
xnor ( n12993 , n12983 , n12992 );
buf ( n12994 , n12993 );
and ( n12995 , n12955 , n12994 );
not ( n12996 , n12955 );
not ( n12997 , n12982 );
not ( n12998 , n12992 );
or ( n12999 , n12997 , n12998 );
or ( n13000 , n12982 , n12992 );
nand ( n13001 , n12999 , n13000 );
not ( n13002 , n12973 );
and ( n13003 , n13001 , n13002 );
not ( n13004 , n13001 );
and ( n13005 , n13004 , n12973 );
nor ( n13006 , n13003 , n13005 );
buf ( n13007 , n13006 );
and ( n13008 , n12996 , n13007 );
nor ( n13009 , n12995 , n13008 );
buf ( n13010 , n5306 );
not ( n13011 , n13010 );
not ( n13012 , n13011 );
buf ( n13013 , n5307 );
buf ( n13014 , n13013 );
not ( n13015 , n13014 );
buf ( n13016 , n5308 );
not ( n13017 , n13016 );
not ( n13018 , n13017 );
or ( n13019 , n13015 , n13018 );
not ( n13020 , n13013 );
buf ( n13021 , n13016 );
nand ( n13022 , n13020 , n13021 );
nand ( n13023 , n13019 , n13022 );
not ( n13024 , n13023 );
or ( n13025 , n13012 , n13024 );
or ( n13026 , n13023 , n13011 );
nand ( n13027 , n13025 , n13026 );
not ( n13028 , n13027 );
buf ( n13029 , n5309 );
buf ( n13030 , n5310 );
not ( n13031 , n13030 );
xor ( n13032 , n13029 , n13031 );
buf ( n13033 , n5311 );
not ( n13034 , n13033 );
buf ( n13035 , n5312 );
nand ( n13036 , n6577 , n13035 );
not ( n13037 , n13036 );
or ( n13038 , n13034 , n13037 );
nand ( n13039 , n8070 , n13035 );
or ( n13040 , n13039 , n13033 );
nand ( n13041 , n13038 , n13040 );
xnor ( n13042 , n13032 , n13041 );
not ( n13043 , n13042 );
not ( n13044 , n13043 );
or ( n13045 , n13028 , n13044 );
or ( n13046 , n13043 , n13027 );
nand ( n13047 , n13045 , n13046 );
not ( n13048 , n13047 );
buf ( n13049 , n5313 );
buf ( n13050 , n13049 );
not ( n13051 , n13050 );
buf ( n13052 , n5314 );
not ( n13053 , n13052 );
not ( n13054 , n13053 );
or ( n13055 , n13051 , n13054 );
not ( n13056 , n13049 );
buf ( n13057 , n13052 );
nand ( n13058 , n13056 , n13057 );
nand ( n13059 , n13055 , n13058 );
buf ( n13060 , n5315 );
not ( n13061 , n13060 );
and ( n13062 , n13059 , n13061 );
not ( n13063 , n13059 );
buf ( n13064 , n13060 );
and ( n13065 , n13063 , n13064 );
nor ( n13066 , n13062 , n13065 );
buf ( n13067 , n5316 );
nand ( n13068 , n7344 , n13067 );
buf ( n13069 , n5317 );
buf ( n13070 , n13069 );
and ( n13071 , n13068 , n13070 );
not ( n13072 , n13068 );
not ( n13073 , n13069 );
and ( n13074 , n13072 , n13073 );
nor ( n13075 , n13071 , n13074 );
xor ( n13076 , n13066 , n13075 );
buf ( n13077 , n5318 );
nand ( n13078 , n8954 , n13077 );
buf ( n13079 , n5319 );
buf ( n13080 , n13079 );
and ( n13081 , n13078 , n13080 );
not ( n13082 , n13078 );
not ( n13083 , n13079 );
and ( n13084 , n13082 , n13083 );
nor ( n13085 , n13081 , n13084 );
not ( n13086 , n13085 );
xnor ( n13087 , n13076 , n13086 );
buf ( n13088 , n13087 );
not ( n13089 , n13088 );
and ( n13090 , n13048 , n13089 );
and ( n13091 , n13088 , n13047 );
nor ( n13092 , n13090 , n13091 );
nand ( n13093 , n13009 , n13092 );
not ( n13094 , n13093 );
buf ( n13095 , n5320 );
buf ( n13096 , n13095 );
not ( n13097 , n13096 );
buf ( n13098 , n5321 );
not ( n13099 , n13098 );
not ( n13100 , n13099 );
or ( n13101 , n13097 , n13100 );
not ( n13102 , n13095 );
buf ( n13103 , n13098 );
nand ( n13104 , n13102 , n13103 );
nand ( n13105 , n13101 , n13104 );
buf ( n13106 , n5322 );
buf ( n13107 , n13106 );
and ( n13108 , n13105 , n13107 );
not ( n13109 , n13105 );
not ( n13110 , n13106 );
and ( n13111 , n13109 , n13110 );
nor ( n13112 , n13108 , n13111 );
buf ( n13113 , n5323 );
nand ( n13114 , n7563 , n13113 );
buf ( n13115 , n5324 );
buf ( n13116 , n13115 );
and ( n13117 , n13114 , n13116 );
not ( n13118 , n13114 );
not ( n13119 , n13115 );
and ( n13120 , n13118 , n13119 );
nor ( n13121 , n13117 , n13120 );
xor ( n13122 , n13112 , n13121 );
buf ( n13123 , n5325 );
nand ( n13124 , n8454 , n13123 );
buf ( n13125 , n5326 );
buf ( n13126 , n13125 );
and ( n13127 , n13124 , n13126 );
not ( n13128 , n13124 );
not ( n13129 , n13125 );
and ( n13130 , n13128 , n13129 );
nor ( n13131 , n13127 , n13130 );
xnor ( n13132 , n13122 , n13131 );
buf ( n13133 , n13132 );
not ( n13134 , n13133 );
not ( n13135 , n11076 );
buf ( n13136 , n5327 );
buf ( n13137 , n13136 );
not ( n13138 , n13137 );
buf ( n13139 , n5328 );
not ( n13140 , n13139 );
not ( n13141 , n13140 );
or ( n13142 , n13138 , n13141 );
not ( n13143 , n13136 );
buf ( n13144 , n13139 );
nand ( n13145 , n13143 , n13144 );
nand ( n13146 , n13142 , n13145 );
not ( n13147 , n13146 );
not ( n13148 , n13147 );
or ( n13149 , n13135 , n13148 );
or ( n13150 , n13147 , n11076 );
nand ( n13151 , n13149 , n13150 );
not ( n13152 , n13151 );
buf ( n13153 , n5329 );
nand ( n13154 , n8454 , n13153 );
not ( n13155 , n13154 );
buf ( n13156 , n5330 );
not ( n13157 , n13156 );
and ( n13158 , n13155 , n13157 );
nand ( n13159 , n6557 , n13153 );
and ( n13160 , n13159 , n13156 );
nor ( n13161 , n13158 , n13160 );
not ( n13162 , n13161 );
buf ( n13163 , n5331 );
nand ( n13164 , n6577 , n13163 );
buf ( n13165 , n5332 );
not ( n13166 , n13165 );
and ( n13167 , n13164 , n13166 );
not ( n13168 , n13164 );
buf ( n13169 , n13165 );
and ( n13170 , n13168 , n13169 );
nor ( n13171 , n13167 , n13170 );
not ( n13172 , n13171 );
or ( n13173 , n13162 , n13172 );
not ( n13174 , n13171 );
not ( n13175 , n13161 );
nand ( n13176 , n13174 , n13175 );
nand ( n13177 , n13173 , n13176 );
buf ( n13178 , n5333 );
not ( n13179 , n13178 );
and ( n13180 , n13177 , n13179 );
not ( n13181 , n13177 );
buf ( n13182 , n13178 );
and ( n13183 , n13181 , n13182 );
nor ( n13184 , n13180 , n13183 );
not ( n13185 , n13184 );
or ( n13186 , n13152 , n13185 );
or ( n13187 , n13184 , n13151 );
nand ( n13188 , n13186 , n13187 );
not ( n13189 , n13188 );
and ( n13190 , n13134 , n13189 );
and ( n13191 , n13133 , n13188 );
nor ( n13192 , n13190 , n13191 );
not ( n13193 , n13192 );
not ( n13194 , n13193 );
and ( n13195 , n13094 , n13194 );
and ( n13196 , n13093 , n13193 );
nor ( n13197 , n13195 , n13196 );
not ( n13198 , n13197 );
not ( n13199 , n13198 );
or ( n13200 , n12948 , n13199 );
nand ( n13201 , n12946 , n13197 );
nand ( n13202 , n13200 , n13201 );
buf ( n13203 , n5334 );
buf ( n13204 , n13203 );
not ( n13205 , n13204 );
not ( n13206 , n8385 );
or ( n13207 , n13205 , n13206 );
not ( n13208 , n13204 );
nand ( n13209 , n13208 , n8398 );
nand ( n13210 , n13207 , n13209 );
and ( n13211 , n13210 , n8439 );
not ( n13212 , n13210 );
and ( n13213 , n13212 , n8440 );
nor ( n13214 , n13211 , n13213 );
buf ( n13215 , n5335 );
not ( n13216 , n13215 );
buf ( n13217 , n5336 );
nand ( n13218 , n8069 , n13217 );
buf ( n13219 , n5337 );
buf ( n13220 , n13219 );
and ( n13221 , n13218 , n13220 );
not ( n13222 , n13218 );
not ( n13223 , n13219 );
and ( n13224 , n13222 , n13223 );
nor ( n13225 , n13221 , n13224 );
xor ( n13226 , n13216 , n13225 );
buf ( n13227 , n5338 );
nand ( n13228 , n7344 , n13227 );
buf ( n13229 , n5339 );
buf ( n13230 , n13229 );
and ( n13231 , n13228 , n13230 );
not ( n13232 , n13228 );
not ( n13233 , n13229 );
and ( n13234 , n13232 , n13233 );
nor ( n13235 , n13231 , n13234 );
xnor ( n13236 , n13226 , n13235 );
not ( n13237 , n13236 );
buf ( n13238 , n5340 );
buf ( n13239 , n13238 );
not ( n13240 , n13239 );
buf ( n13241 , n5341 );
not ( n13242 , n13241 );
not ( n13243 , n13242 );
or ( n13244 , n13240 , n13243 );
not ( n13245 , n13238 );
buf ( n13246 , n13241 );
nand ( n13247 , n13245 , n13246 );
nand ( n13248 , n13244 , n13247 );
not ( n13249 , n13248 );
not ( n13250 , n13249 );
and ( n13251 , n13237 , n13250 );
and ( n13252 , n13236 , n13249 );
nor ( n13253 , n13251 , n13252 );
buf ( n13254 , n13253 );
not ( n13255 , n13254 );
buf ( n13256 , n5342 );
buf ( n13257 , n13256 );
not ( n13258 , n13257 );
buf ( n13259 , n5343 );
buf ( n13260 , n5344 );
buf ( n13261 , n13260 );
not ( n13262 , n13261 );
buf ( n13263 , n5345 );
not ( n13264 , n13263 );
not ( n13265 , n13264 );
or ( n13266 , n13262 , n13265 );
not ( n13267 , n13260 );
buf ( n13268 , n13263 );
nand ( n13269 , n13267 , n13268 );
nand ( n13270 , n13266 , n13269 );
xor ( n13271 , n13259 , n13270 );
buf ( n13272 , n5346 );
buf ( n13273 , n5347 );
not ( n13274 , n13273 );
xor ( n13275 , n13272 , n13274 );
buf ( n13276 , n5348 );
nand ( n13277 , n7293 , n13276 );
xnor ( n13278 , n13275 , n13277 );
xnor ( n13279 , n13271 , n13278 );
not ( n13280 , n13279 );
not ( n13281 , n13280 );
or ( n13282 , n13258 , n13281 );
or ( n13283 , n13280 , n13257 );
nand ( n13284 , n13282 , n13283 );
not ( n13285 , n13284 );
and ( n13286 , n13255 , n13285 );
and ( n13287 , n13254 , n13284 );
nor ( n13288 , n13286 , n13287 );
not ( n13289 , n13288 );
nand ( n13290 , n13214 , n13289 );
not ( n13291 , n13290 );
xor ( n13292 , n12320 , n12339 );
not ( n13293 , n12329 );
xor ( n13294 , n13292 , n13293 );
buf ( n13295 , n5349 );
nand ( n13296 , n7258 , n13295 );
buf ( n13297 , n5350 );
buf ( n13298 , n13297 );
and ( n13299 , n13296 , n13298 );
not ( n13300 , n13296 );
not ( n13301 , n13297 );
and ( n13302 , n13300 , n13301 );
nor ( n13303 , n13299 , n13302 );
nor ( n13304 , n13294 , n13303 );
not ( n13305 , n13304 );
nand ( n13306 , n13303 , n13294 );
nand ( n13307 , n13305 , n13306 );
not ( n13308 , n12376 );
and ( n13309 , n13307 , n13308 );
not ( n13310 , n13307 );
and ( n13311 , n13310 , n12379 );
nor ( n13312 , n13309 , n13311 );
not ( n13313 , n13312 );
and ( n13314 , n13291 , n13313 );
and ( n13315 , n13290 , n13312 );
nor ( n13316 , n13314 , n13315 );
and ( n13317 , n13202 , n13316 );
not ( n13318 , n13202 );
not ( n13319 , n13316 );
and ( n13320 , n13318 , n13319 );
nor ( n13321 , n13317 , n13320 );
xor ( n13322 , n12843 , n13321 );
buf ( n13323 , n13322 );
and ( n13324 , n12405 , n13323 );
not ( n13325 , n12405 );
not ( n13326 , n13321 );
not ( n13327 , n13326 );
not ( n13328 , n12843 );
not ( n13329 , n13328 );
or ( n13330 , n13327 , n13329 );
nand ( n13331 , n13321 , n12843 );
nand ( n13332 , n13330 , n13331 );
buf ( n13333 , n13332 );
and ( n13334 , n13325 , n13333 );
nor ( n13335 , n13324 , n13334 );
not ( n13336 , n13335 );
nand ( n13337 , n11304 , n13336 );
buf ( n13338 , n11337 );
buf ( n13339 , n6496 );
nor ( n13340 , n13338 , n13339 );
buf ( n13341 , n5351 );
not ( n13342 , n13341 );
not ( n13343 , n13342 );
or ( n13344 , n13340 , n13343 );
buf ( n13345 , n13344 );
buf ( n13346 , n13345 );
not ( n13347 , n13346 );
nand ( n13348 , n9095 , n13337 , n13347 );
buf ( n13349 , n13345 );
nor ( n13350 , n13335 , n13349 );
nand ( n13351 , n9094 , n13350 , n11304 );
and ( n13352 , n13340 , n13342 );
buf ( n13353 , n13352 );
buf ( n13354 , n5352 );
buf ( n13355 , n13354 );
nand ( n13356 , n13353 , n13355 );
nand ( n13357 , n13348 , n13351 , n13356 );
buf ( n13358 , n13357 );
buf ( n13359 , n13358 );
buf ( n13360 , n5353 );
buf ( n13361 , n13360 );
not ( n13362 , n13361 );
buf ( n13363 , n5354 );
not ( n13364 , n13363 );
not ( n13365 , n13364 );
or ( n13366 , n13362 , n13365 );
not ( n13367 , n13360 );
buf ( n13368 , n13363 );
nand ( n13369 , n13367 , n13368 );
nand ( n13370 , n13366 , n13369 );
buf ( n13371 , n5355 );
buf ( n13372 , n13371 );
and ( n13373 , n13370 , n13372 );
not ( n13374 , n13370 );
not ( n13375 , n13371 );
and ( n13376 , n13374 , n13375 );
nor ( n13377 , n13373 , n13376 );
buf ( n13378 , n5356 );
nand ( n13379 , n8454 , n13378 );
buf ( n13380 , n5357 );
buf ( n13381 , n13380 );
and ( n13382 , n13379 , n13381 );
not ( n13383 , n13379 );
not ( n13384 , n13380 );
and ( n13385 , n13383 , n13384 );
nor ( n13386 , n13382 , n13385 );
not ( n13387 , n13386 );
xor ( n13388 , n13377 , n13387 );
buf ( n13389 , n5358 );
nand ( n13390 , n11946 , n13389 );
buf ( n13391 , n5359 );
not ( n13392 , n13391 );
and ( n13393 , n13390 , n13392 );
not ( n13394 , n13390 );
buf ( n13395 , n13391 );
and ( n13396 , n13394 , n13395 );
nor ( n13397 , n13393 , n13396 );
xnor ( n13398 , n13388 , n13397 );
buf ( n13399 , n13398 );
not ( n13400 , n13399 );
buf ( n13401 , n5360 );
buf ( n13402 , n13401 );
not ( n13403 , n13402 );
buf ( n13404 , n5361 );
nand ( n13405 , n8454 , n13404 );
buf ( n13406 , n5362 );
buf ( n13407 , n13406 );
and ( n13408 , n13405 , n13407 );
not ( n13409 , n13405 );
not ( n13410 , n13406 );
and ( n13411 , n13409 , n13410 );
nor ( n13412 , n13408 , n13411 );
not ( n13413 , n13412 );
buf ( n13414 , n5363 );
nand ( n13415 , n6577 , n13414 );
buf ( n13416 , n5364 );
not ( n13417 , n13416 );
and ( n13418 , n13415 , n13417 );
not ( n13419 , n13415 );
buf ( n13420 , n13416 );
and ( n13421 , n13419 , n13420 );
nor ( n13422 , n13418 , n13421 );
not ( n13423 , n13422 );
or ( n13424 , n13413 , n13423 );
or ( n13425 , n13412 , n13422 );
nand ( n13426 , n13424 , n13425 );
buf ( n13427 , n5365 );
buf ( n13428 , n13427 );
not ( n13429 , n13428 );
buf ( n13430 , n5366 );
not ( n13431 , n13430 );
not ( n13432 , n13431 );
or ( n13433 , n13429 , n13432 );
not ( n13434 , n13427 );
buf ( n13435 , n13430 );
nand ( n13436 , n13434 , n13435 );
nand ( n13437 , n13433 , n13436 );
buf ( n13438 , n5367 );
not ( n13439 , n13438 );
and ( n13440 , n13437 , n13439 );
not ( n13441 , n13437 );
buf ( n13442 , n13438 );
and ( n13443 , n13441 , n13442 );
nor ( n13444 , n13440 , n13443 );
xor ( n13445 , n13426 , n13444 );
buf ( n13446 , n13445 );
not ( n13447 , n13446 );
or ( n13448 , n13403 , n13447 );
or ( n13449 , n13446 , n13402 );
nand ( n13450 , n13448 , n13449 );
not ( n13451 , n13450 );
or ( n13452 , n13400 , n13451 );
or ( n13453 , n13450 , n13399 );
nand ( n13454 , n13452 , n13453 );
not ( n13455 , n13454 );
xor ( n13456 , n9968 , n9978 );
xnor ( n13457 , n13456 , n9988 );
buf ( n13458 , n13457 );
xor ( n13459 , n10557 , n13458 );
xnor ( n13460 , n13459 , n10011 );
not ( n13461 , n13460 );
nand ( n13462 , n13455 , n13461 );
not ( n13463 , n13462 );
buf ( n13464 , n5368 );
buf ( n13465 , n13464 );
not ( n13466 , n13465 );
buf ( n13467 , n5369 );
not ( n13468 , n13467 );
not ( n13469 , n13468 );
or ( n13470 , n13466 , n13469 );
not ( n13471 , n13464 );
buf ( n13472 , n13467 );
nand ( n13473 , n13471 , n13472 );
nand ( n13474 , n13470 , n13473 );
buf ( n13475 , n5370 );
not ( n13476 , n13475 );
and ( n13477 , n13474 , n13476 );
not ( n13478 , n13474 );
buf ( n13479 , n13475 );
and ( n13480 , n13478 , n13479 );
nor ( n13481 , n13477 , n13480 );
buf ( n13482 , n5371 );
nand ( n13483 , n7698 , n13482 );
buf ( n13484 , n5372 );
buf ( n13485 , n13484 );
and ( n13486 , n13483 , n13485 );
not ( n13487 , n13483 );
not ( n13488 , n13484 );
and ( n13489 , n13487 , n13488 );
nor ( n13490 , n13486 , n13489 );
xor ( n13491 , n13481 , n13490 );
buf ( n13492 , n5373 );
nand ( n13493 , n10165 , n13492 );
buf ( n13494 , n5374 );
not ( n13495 , n13494 );
and ( n13496 , n13493 , n13495 );
not ( n13497 , n13493 );
buf ( n13498 , n13494 );
and ( n13499 , n13497 , n13498 );
nor ( n13500 , n13496 , n13499 );
buf ( n13501 , n13500 );
xnor ( n13502 , n13491 , n13501 );
buf ( n13503 , n5375 );
buf ( n13504 , n13503 );
nand ( n13505 , n13502 , n13504 );
not ( n13506 , n13505 );
nor ( n13507 , n13502 , n13504 );
nor ( n13508 , n13506 , n13507 );
not ( n13509 , n13508 );
not ( n13510 , n7219 );
not ( n13511 , n13510 );
not ( n13512 , n7206 );
or ( n13513 , n13511 , n13512 );
or ( n13514 , n7206 , n13510 );
nand ( n13515 , n13513 , n13514 );
buf ( n13516 , n13515 );
not ( n13517 , n13516 );
or ( n13518 , n13509 , n13517 );
or ( n13519 , n13516 , n13508 );
nand ( n13520 , n13518 , n13519 );
not ( n13521 , n13520 );
not ( n13522 , n13521 );
not ( n13523 , n13522 );
and ( n13524 , n13463 , n13523 );
not ( n13525 , n13454 );
nand ( n13526 , n13525 , n13461 );
and ( n13527 , n13526 , n13522 );
nor ( n13528 , n13524 , n13527 );
buf ( n13529 , n13528 );
not ( n13530 , n13529 );
not ( n13531 , n11789 );
not ( n13532 , n13531 );
not ( n13533 , n11818 );
not ( n13534 , n13533 );
or ( n13535 , n13532 , n13534 );
nand ( n13536 , n11818 , n11789 );
nand ( n13537 , n13535 , n13536 );
not ( n13538 , n13537 );
not ( n13539 , n13538 );
not ( n13540 , n10342 );
not ( n13541 , n11154 );
or ( n13542 , n13540 , n13541 );
or ( n13543 , n11154 , n10342 );
nand ( n13544 , n13542 , n13543 );
not ( n13545 , n13544 );
and ( n13546 , n13539 , n13545 );
buf ( n13547 , n13538 );
and ( n13548 , n13547 , n13544 );
nor ( n13549 , n13546 , n13548 );
not ( n13550 , n8786 );
not ( n13551 , n13550 );
buf ( n13552 , n5376 );
buf ( n13553 , n13552 );
not ( n13554 , n13553 );
not ( n13555 , n11187 );
buf ( n13556 , n5377 );
not ( n13557 , n13556 );
not ( n13558 , n13557 );
or ( n13559 , n13555 , n13558 );
not ( n13560 , n11186 );
buf ( n13561 , n13556 );
nand ( n13562 , n13560 , n13561 );
nand ( n13563 , n13559 , n13562 );
and ( n13564 , n13563 , n11863 );
not ( n13565 , n13563 );
not ( n13566 , n11862 );
and ( n13567 , n13565 , n13566 );
nor ( n13568 , n13564 , n13567 );
not ( n13569 , n13568 );
buf ( n13570 , n5378 );
nand ( n13571 , n8375 , n13570 );
buf ( n13572 , n5379 );
buf ( n13573 , n13572 );
and ( n13574 , n13571 , n13573 );
not ( n13575 , n13571 );
not ( n13576 , n13572 );
and ( n13577 , n13575 , n13576 );
nor ( n13578 , n13574 , n13577 );
buf ( n13579 , n13578 );
xor ( n13580 , n13569 , n13579 );
buf ( n13581 , n6577 );
buf ( n13582 , n5380 );
nand ( n13583 , n13581 , n13582 );
buf ( n13584 , n5381 );
not ( n13585 , n13584 );
and ( n13586 , n13583 , n13585 );
not ( n13587 , n13583 );
buf ( n13588 , n13584 );
and ( n13589 , n13587 , n13588 );
nor ( n13590 , n13586 , n13589 );
xnor ( n13591 , n13580 , n13590 );
not ( n13592 , n13591 );
or ( n13593 , n13554 , n13592 );
xor ( n13594 , n13568 , n13578 );
xnor ( n13595 , n13594 , n13590 );
not ( n13596 , n13552 );
nand ( n13597 , n13595 , n13596 );
nand ( n13598 , n13593 , n13597 );
not ( n13599 , n13598 );
and ( n13600 , n13551 , n13599 );
and ( n13601 , n13550 , n13598 );
nor ( n13602 , n13600 , n13601 );
not ( n13603 , n13602 );
nand ( n13604 , n13549 , n13603 );
buf ( n13605 , n5382 );
buf ( n13606 , n13605 );
buf ( n13607 , n5383 );
buf ( n13608 , n13607 );
not ( n13609 , n13608 );
buf ( n13610 , n5384 );
not ( n13611 , n13610 );
not ( n13612 , n13611 );
or ( n13613 , n13609 , n13612 );
not ( n13614 , n13607 );
buf ( n13615 , n13610 );
nand ( n13616 , n13614 , n13615 );
nand ( n13617 , n13613 , n13616 );
xor ( n13618 , n13606 , n13617 );
buf ( n13619 , n5385 );
nand ( n13620 , n6633 , n13619 );
buf ( n13621 , n5386 );
buf ( n13622 , n13621 );
and ( n13623 , n13620 , n13622 );
not ( n13624 , n13620 );
not ( n13625 , n13621 );
and ( n13626 , n13624 , n13625 );
nor ( n13627 , n13623 , n13626 );
not ( n13628 , n13627 );
buf ( n13629 , n5387 );
nand ( n13630 , n6815 , n13629 );
buf ( n13631 , n5388 );
not ( n13632 , n13631 );
and ( n13633 , n13630 , n13632 );
not ( n13634 , n13630 );
buf ( n13635 , n13631 );
and ( n13636 , n13634 , n13635 );
nor ( n13637 , n13633 , n13636 );
not ( n13638 , n13637 );
or ( n13639 , n13628 , n13638 );
or ( n13640 , n13627 , n13637 );
nand ( n13641 , n13639 , n13640 );
xnor ( n13642 , n13618 , n13641 );
not ( n13643 , n13642 );
buf ( n13644 , n5389 );
buf ( n13645 , n13644 );
not ( n13646 , n13645 );
buf ( n13647 , n5390 );
not ( n13648 , n13647 );
not ( n13649 , n13648 );
or ( n13650 , n13646 , n13649 );
not ( n13651 , n13644 );
buf ( n13652 , n13647 );
nand ( n13653 , n13651 , n13652 );
nand ( n13654 , n13650 , n13653 );
buf ( n13655 , n5391 );
buf ( n13656 , n13655 );
and ( n13657 , n13654 , n13656 );
not ( n13658 , n13654 );
not ( n13659 , n13655 );
and ( n13660 , n13658 , n13659 );
nor ( n13661 , n13657 , n13660 );
buf ( n13662 , n5392 );
nand ( n13663 , n6815 , n13662 );
buf ( n13664 , n5393 );
xor ( n13665 , n13663 , n13664 );
xor ( n13666 , n13661 , n13665 );
buf ( n13667 , n5394 );
nand ( n13668 , n8260 , n13667 );
buf ( n13669 , n5395 );
not ( n13670 , n13669 );
and ( n13671 , n13668 , n13670 );
not ( n13672 , n13668 );
buf ( n13673 , n13669 );
and ( n13674 , n13672 , n13673 );
nor ( n13675 , n13671 , n13674 );
xnor ( n13676 , n13666 , n13675 );
not ( n13677 , n13676 );
buf ( n13678 , n5396 );
nand ( n13679 , n7698 , n13678 );
buf ( n13680 , n5397 );
buf ( n13681 , n13680 );
and ( n13682 , n13679 , n13681 );
not ( n13683 , n13679 );
not ( n13684 , n13680 );
and ( n13685 , n13683 , n13684 );
nor ( n13686 , n13682 , n13685 );
buf ( n13687 , n13686 );
not ( n13688 , n13687 );
and ( n13689 , n13677 , n13688 );
not ( n13690 , n13676 );
not ( n13691 , n13690 );
and ( n13692 , n13691 , n13687 );
nor ( n13693 , n13689 , n13692 );
not ( n13694 , n13693 );
and ( n13695 , n13643 , n13694 );
not ( n13696 , n13643 );
and ( n13697 , n13696 , n13693 );
nor ( n13698 , n13695 , n13697 );
not ( n13699 , n13698 );
and ( n13700 , n13604 , n13699 );
not ( n13701 , n13604 );
and ( n13702 , n13701 , n13698 );
nor ( n13703 , n13700 , n13702 );
not ( n13704 , n13703 );
not ( n13705 , n13704 );
buf ( n13706 , n5398 );
buf ( n13707 , n13706 );
not ( n13708 , n13707 );
not ( n13709 , n7450 );
or ( n13710 , n13708 , n13709 );
buf ( n13711 , n7449 );
not ( n13712 , n13711 );
or ( n13713 , n13712 , n13707 );
nand ( n13714 , n13710 , n13713 );
not ( n13715 , n13714 );
not ( n13716 , n7495 );
and ( n13717 , n13715 , n13716 );
buf ( n13718 , n7494 );
and ( n13719 , n13714 , n13718 );
nor ( n13720 , n13717 , n13719 );
buf ( n13721 , n5399 );
buf ( n13722 , n13721 );
not ( n13723 , n13722 );
buf ( n13724 , n11857 );
not ( n13725 , n13724 );
or ( n13726 , n13723 , n13725 );
not ( n13727 , n13722 );
nand ( n13728 , n13727 , n11858 );
nand ( n13729 , n13726 , n13728 );
not ( n13730 , n12897 );
not ( n13731 , n13730 );
and ( n13732 , n13729 , n13731 );
not ( n13733 , n13729 );
not ( n13734 , n12881 );
not ( n13735 , n12890 );
not ( n13736 , n12896 );
or ( n13737 , n13735 , n13736 );
or ( n13738 , n12890 , n12896 );
nand ( n13739 , n13737 , n13738 );
not ( n13740 , n13739 );
or ( n13741 , n13734 , n13740 );
or ( n13742 , n13739 , n12881 );
nand ( n13743 , n13741 , n13742 );
buf ( n13744 , n13743 );
and ( n13745 , n13733 , n13744 );
nor ( n13746 , n13732 , n13745 );
not ( n13747 , n13746 );
nand ( n13748 , n13720 , n13747 );
not ( n13749 , n13748 );
buf ( n13750 , n5400 );
buf ( n13751 , n13750 );
not ( n13752 , n13751 );
buf ( n13753 , n5401 );
not ( n13754 , n13753 );
not ( n13755 , n13754 );
or ( n13756 , n13752 , n13755 );
not ( n13757 , n13750 );
buf ( n13758 , n13753 );
nand ( n13759 , n13757 , n13758 );
nand ( n13760 , n13756 , n13759 );
buf ( n13761 , n5402 );
not ( n13762 , n13761 );
and ( n13763 , n13760 , n13762 );
not ( n13764 , n13760 );
buf ( n13765 , n13761 );
and ( n13766 , n13764 , n13765 );
nor ( n13767 , n13763 , n13766 );
buf ( n13768 , n5403 );
nand ( n13769 , n6502 , n13768 );
buf ( n13770 , n5404 );
buf ( n13771 , n13770 );
and ( n13772 , n13769 , n13771 );
not ( n13773 , n13769 );
not ( n13774 , n13770 );
and ( n13775 , n13773 , n13774 );
nor ( n13776 , n13772 , n13775 );
xor ( n13777 , n13767 , n13776 );
buf ( n13778 , n5405 );
nand ( n13779 , n7912 , n13778 );
not ( n13780 , n13354 );
and ( n13781 , n13779 , n13780 );
not ( n13782 , n13779 );
and ( n13783 , n13782 , n13355 );
nor ( n13784 , n13781 , n13783 );
xor ( n13785 , n13777 , n13784 );
not ( n13786 , n13785 );
not ( n13787 , n13786 );
buf ( n13788 , n5406 );
buf ( n13789 , n13788 );
not ( n13790 , n13789 );
buf ( n13791 , n5407 );
nand ( n13792 , n8966 , n13791 );
buf ( n13793 , n5408 );
buf ( n13794 , n13793 );
and ( n13795 , n13792 , n13794 );
not ( n13796 , n13792 );
not ( n13797 , n13793 );
and ( n13798 , n13796 , n13797 );
nor ( n13799 , n13795 , n13798 );
not ( n13800 , n13799 );
buf ( n13801 , n5409 );
nand ( n13802 , n8954 , n13801 );
buf ( n13803 , n5410 );
not ( n13804 , n13803 );
and ( n13805 , n13802 , n13804 );
not ( n13806 , n13802 );
buf ( n13807 , n13803 );
and ( n13808 , n13806 , n13807 );
nor ( n13809 , n13805 , n13808 );
not ( n13810 , n13809 );
or ( n13811 , n13800 , n13810 );
or ( n13812 , n13799 , n13809 );
nand ( n13813 , n13811 , n13812 );
buf ( n13814 , n5411 );
buf ( n13815 , n13814 );
not ( n13816 , n13815 );
buf ( n13817 , n5412 );
not ( n13818 , n13817 );
not ( n13819 , n13818 );
or ( n13820 , n13816 , n13819 );
not ( n13821 , n13814 );
buf ( n13822 , n13817 );
nand ( n13823 , n13821 , n13822 );
nand ( n13824 , n13820 , n13823 );
buf ( n13825 , n5413 );
not ( n13826 , n13825 );
and ( n13827 , n13824 , n13826 );
not ( n13828 , n13824 );
buf ( n13829 , n13825 );
and ( n13830 , n13828 , n13829 );
nor ( n13831 , n13827 , n13830 );
xor ( n13832 , n13813 , n13831 );
not ( n13833 , n13832 );
or ( n13834 , n13790 , n13833 );
not ( n13835 , n13809 );
xor ( n13836 , n13831 , n13835 );
buf ( n13837 , n13799 );
xnor ( n13838 , n13836 , n13837 );
not ( n13839 , n13788 );
nand ( n13840 , n13838 , n13839 );
nand ( n13841 , n13834 , n13840 );
not ( n13842 , n13841 );
or ( n13843 , n13787 , n13842 );
or ( n13844 , n13841 , n13786 );
nand ( n13845 , n13843 , n13844 );
buf ( n13846 , n13845 );
not ( n13847 , n13846 );
and ( n13848 , n13749 , n13847 );
and ( n13849 , n13748 , n13846 );
nor ( n13850 , n13848 , n13849 );
not ( n13851 , n13850 );
not ( n13852 , n13851 );
or ( n13853 , n13705 , n13852 );
nand ( n13854 , n13850 , n13703 );
nand ( n13855 , n13853 , n13854 );
buf ( n13856 , n5414 );
buf ( n13857 , n13856 );
not ( n13858 , n9643 );
xor ( n13859 , n13857 , n13858 );
xnor ( n13860 , n13859 , n9598 );
buf ( n13861 , n5415 );
buf ( n13862 , n13861 );
not ( n13863 , n13862 );
not ( n13864 , n9181 );
or ( n13865 , n13863 , n13864 );
or ( n13866 , n9181 , n13862 );
nand ( n13867 , n13865 , n13866 );
buf ( n13868 , n5416 );
buf ( n13869 , n13868 );
not ( n13870 , n13869 );
buf ( n13871 , n5417 );
not ( n13872 , n13871 );
not ( n13873 , n13872 );
or ( n13874 , n13870 , n13873 );
not ( n13875 , n13868 );
buf ( n13876 , n13871 );
nand ( n13877 , n13875 , n13876 );
nand ( n13878 , n13874 , n13877 );
buf ( n13879 , n5418 );
buf ( n13880 , n13879 );
and ( n13881 , n13878 , n13880 );
not ( n13882 , n13878 );
not ( n13883 , n13879 );
and ( n13884 , n13882 , n13883 );
nor ( n13885 , n13881 , n13884 );
buf ( n13886 , n5419 );
nand ( n13887 , n8124 , n13886 );
buf ( n13888 , n5420 );
buf ( n13889 , n13888 );
and ( n13890 , n13887 , n13889 );
not ( n13891 , n13887 );
not ( n13892 , n13888 );
and ( n13893 , n13891 , n13892 );
nor ( n13894 , n13890 , n13893 );
xor ( n13895 , n13885 , n13894 );
buf ( n13896 , n5421 );
nand ( n13897 , n8125 , n13896 );
buf ( n13898 , n5422 );
not ( n13899 , n13898 );
and ( n13900 , n13897 , n13899 );
not ( n13901 , n13897 );
buf ( n13902 , n13898 );
and ( n13903 , n13901 , n13902 );
nor ( n13904 , n13900 , n13903 );
xnor ( n13905 , n13895 , n13904 );
not ( n13906 , n13905 );
not ( n13907 , n13906 );
and ( n13908 , n13867 , n13907 );
not ( n13909 , n13867 );
and ( n13910 , n13909 , n13906 );
nor ( n13911 , n13908 , n13910 );
not ( n13912 , n13911 );
nand ( n13913 , n13860 , n13912 );
not ( n13914 , n13913 );
buf ( n13915 , n5423 );
buf ( n13916 , n13915 );
buf ( n13917 , n5424 );
buf ( n13918 , n13917 );
not ( n13919 , n13918 );
buf ( n13920 , n5425 );
not ( n13921 , n13920 );
not ( n13922 , n13921 );
or ( n13923 , n13919 , n13922 );
not ( n13924 , n13917 );
buf ( n13925 , n13920 );
nand ( n13926 , n13924 , n13925 );
nand ( n13927 , n13923 , n13926 );
xor ( n13928 , n13916 , n13927 );
buf ( n13929 , n5426 );
buf ( n13930 , n5427 );
xor ( n13931 , n13929 , n13930 );
buf ( n13932 , n5428 );
nand ( n13933 , n11847 , n13932 );
xnor ( n13934 , n13931 , n13933 );
xnor ( n13935 , n13928 , n13934 );
buf ( n13936 , n13935 );
not ( n13937 , n13936 );
not ( n13938 , n9511 );
buf ( n13939 , n5429 );
nand ( n13940 , n7344 , n13939 );
buf ( n13941 , n5430 );
buf ( n13942 , n13941 );
and ( n13943 , n13940 , n13942 );
not ( n13944 , n13940 );
not ( n13945 , n13941 );
and ( n13946 , n13944 , n13945 );
nor ( n13947 , n13943 , n13946 );
not ( n13948 , n13947 );
buf ( n13949 , n5431 );
nand ( n13950 , n6871 , n13949 );
buf ( n13951 , n5432 );
not ( n13952 , n13951 );
and ( n13953 , n13950 , n13952 );
not ( n13954 , n13950 );
buf ( n13955 , n13951 );
and ( n13956 , n13954 , n13955 );
nor ( n13957 , n13953 , n13956 );
not ( n13958 , n13957 );
or ( n13959 , n13948 , n13958 );
or ( n13960 , n13947 , n13957 );
nand ( n13961 , n13959 , n13960 );
buf ( n13962 , n5433 );
buf ( n13963 , n13962 );
not ( n13964 , n13963 );
buf ( n13965 , n5434 );
not ( n13966 , n13965 );
not ( n13967 , n13966 );
or ( n13968 , n13964 , n13967 );
not ( n13969 , n13962 );
buf ( n13970 , n13965 );
nand ( n13971 , n13969 , n13970 );
nand ( n13972 , n13968 , n13971 );
buf ( n13973 , n5435 );
not ( n13974 , n13973 );
and ( n13975 , n13972 , n13974 );
not ( n13976 , n13972 );
buf ( n13977 , n13973 );
and ( n13978 , n13976 , n13977 );
nor ( n13979 , n13975 , n13978 );
and ( n13980 , n13961 , n13979 );
not ( n13981 , n13961 );
not ( n13982 , n13979 );
and ( n13983 , n13981 , n13982 );
nor ( n13984 , n13980 , n13983 );
not ( n13985 , n13984 );
or ( n13986 , n13938 , n13985 );
not ( n13987 , n9511 );
not ( n13988 , n13957 );
xor ( n13989 , n13979 , n13988 );
buf ( n13990 , n13947 );
xnor ( n13991 , n13989 , n13990 );
nand ( n13992 , n13987 , n13991 );
nand ( n13993 , n13986 , n13992 );
not ( n13994 , n13993 );
and ( n13995 , n13937 , n13994 );
and ( n13996 , n13936 , n13993 );
nor ( n13997 , n13995 , n13996 );
not ( n13998 , n13997 );
not ( n13999 , n13998 );
and ( n14000 , n13914 , n13999 );
and ( n14001 , n13913 , n13998 );
nor ( n14002 , n14000 , n14001 );
not ( n14003 , n14002 );
and ( n14004 , n13855 , n14003 );
not ( n14005 , n13855 );
and ( n14006 , n14005 , n14002 );
nor ( n14007 , n14004 , n14006 );
nand ( n14008 , n13454 , n13521 );
not ( n14009 , n14008 );
buf ( n14010 , n6716 );
not ( n14011 , n14010 );
not ( n14012 , n12951 );
buf ( n14013 , n5436 );
not ( n14014 , n14013 );
not ( n14015 , n14014 );
or ( n14016 , n14012 , n14015 );
not ( n14017 , n12950 );
buf ( n14018 , n14013 );
nand ( n14019 , n14017 , n14018 );
nand ( n14020 , n14016 , n14019 );
buf ( n14021 , n5437 );
not ( n14022 , n14021 );
and ( n14023 , n14020 , n14022 );
not ( n14024 , n14020 );
buf ( n14025 , n14021 );
and ( n14026 , n14024 , n14025 );
nor ( n14027 , n14023 , n14026 );
buf ( n14028 , n5438 );
nand ( n14029 , n6927 , n14028 );
buf ( n14030 , n5439 );
buf ( n14031 , n14030 );
and ( n14032 , n14029 , n14031 );
not ( n14033 , n14029 );
not ( n14034 , n14030 );
and ( n14035 , n14033 , n14034 );
nor ( n14036 , n14032 , n14035 );
xor ( n14037 , n14027 , n14036 );
buf ( n14038 , n5440 );
nand ( n14039 , n8455 , n14038 );
buf ( n14040 , n5441 );
not ( n14041 , n14040 );
and ( n14042 , n14039 , n14041 );
not ( n14043 , n14039 );
buf ( n14044 , n14040 );
and ( n14045 , n14043 , n14044 );
nor ( n14046 , n14042 , n14045 );
xnor ( n14047 , n14037 , n14046 );
not ( n14048 , n14047 );
not ( n14049 , n14048 );
or ( n14050 , n14011 , n14049 );
buf ( n14051 , n14047 );
not ( n14052 , n14051 );
or ( n14053 , n14052 , n14010 );
nand ( n14054 , n14050 , n14053 );
buf ( n14055 , n5442 );
buf ( n14056 , n14055 );
not ( n14057 , n14056 );
buf ( n14058 , n5443 );
not ( n14059 , n14058 );
not ( n14060 , n14059 );
or ( n14061 , n14057 , n14060 );
not ( n14062 , n14055 );
buf ( n14063 , n14058 );
nand ( n14064 , n14062 , n14063 );
nand ( n14065 , n14061 , n14064 );
buf ( n14066 , n5444 );
not ( n14067 , n14066 );
and ( n14068 , n14065 , n14067 );
not ( n14069 , n14065 );
buf ( n14070 , n14066 );
and ( n14071 , n14069 , n14070 );
nor ( n14072 , n14068 , n14071 );
buf ( n14073 , n5445 );
nand ( n14074 , n6577 , n14073 );
buf ( n14075 , n5446 );
buf ( n14076 , n14075 );
and ( n14077 , n14074 , n14076 );
not ( n14078 , n14074 );
not ( n14079 , n14075 );
and ( n14080 , n14078 , n14079 );
nor ( n14081 , n14077 , n14080 );
xor ( n14082 , n14072 , n14081 );
buf ( n14083 , n5447 );
nand ( n14084 , n10383 , n14083 );
buf ( n14085 , n5448 );
buf ( n14086 , n14085 );
and ( n14087 , n14084 , n14086 );
not ( n14088 , n14084 );
not ( n14089 , n14085 );
and ( n14090 , n14088 , n14089 );
nor ( n14091 , n14087 , n14090 );
xnor ( n14092 , n14082 , n14091 );
not ( n14093 , n14092 );
not ( n14094 , n14093 );
not ( n14095 , n14094 );
xor ( n14096 , n14054 , n14095 );
not ( n14097 , n14096 );
not ( n14098 , n14097 );
and ( n14099 , n14009 , n14098 );
and ( n14100 , n14008 , n14097 );
nor ( n14101 , n14099 , n14100 );
not ( n14102 , n14101 );
buf ( n14103 , n5449 );
nand ( n14104 , n6577 , n14103 );
buf ( n14105 , n5450 );
buf ( n14106 , n14105 );
and ( n14107 , n14104 , n14106 );
not ( n14108 , n14104 );
not ( n14109 , n14105 );
and ( n14110 , n14108 , n14109 );
nor ( n14111 , n14107 , n14110 );
buf ( n14112 , n14111 );
buf ( n14113 , n5451 );
buf ( n14114 , n14113 );
not ( n14115 , n14114 );
buf ( n14116 , n5452 );
not ( n14117 , n14116 );
not ( n14118 , n14117 );
or ( n14119 , n14115 , n14118 );
not ( n14120 , n14113 );
buf ( n14121 , n14116 );
nand ( n14122 , n14120 , n14121 );
nand ( n14123 , n14119 , n14122 );
buf ( n14124 , n5453 );
buf ( n14125 , n14124 );
and ( n14126 , n14123 , n14125 );
not ( n14127 , n14123 );
not ( n14128 , n14124 );
and ( n14129 , n14127 , n14128 );
nor ( n14130 , n14126 , n14129 );
buf ( n14131 , n5454 );
nand ( n14132 , n6647 , n14131 );
buf ( n14133 , n5455 );
buf ( n14134 , n14133 );
and ( n14135 , n14132 , n14134 );
not ( n14136 , n14132 );
not ( n14137 , n14133 );
and ( n14138 , n14136 , n14137 );
nor ( n14139 , n14135 , n14138 );
xor ( n14140 , n14130 , n14139 );
buf ( n14141 , n5456 );
nand ( n14142 , n7014 , n14141 );
buf ( n14143 , n5457 );
buf ( n14144 , n14143 );
and ( n14145 , n14142 , n14144 );
not ( n14146 , n14142 );
not ( n14147 , n14143 );
and ( n14148 , n14146 , n14147 );
nor ( n14149 , n14145 , n14148 );
not ( n14150 , n14149 );
xnor ( n14151 , n14140 , n14150 );
buf ( n14152 , n14151 );
not ( n14153 , n14152 );
xor ( n14154 , n14112 , n14153 );
buf ( n14155 , n5458 );
buf ( n14156 , n5459 );
buf ( n14157 , n14156 );
not ( n14158 , n14157 );
buf ( n14159 , n5460 );
not ( n14160 , n14159 );
not ( n14161 , n14160 );
or ( n14162 , n14158 , n14161 );
not ( n14163 , n14156 );
buf ( n14164 , n14159 );
nand ( n14165 , n14163 , n14164 );
nand ( n14166 , n14162 , n14165 );
xor ( n14167 , n14155 , n14166 );
buf ( n14168 , n5461 );
buf ( n14169 , n5462 );
xor ( n14170 , n14168 , n14169 );
buf ( n14171 , n5463 );
nand ( n14172 , n6719 , n14171 );
xnor ( n14173 , n14170 , n14172 );
xnor ( n14174 , n14167 , n14173 );
not ( n14175 , n14174 );
xnor ( n14176 , n14154 , n14175 );
not ( n14177 , n14176 );
not ( n14178 , n14177 );
buf ( n14179 , n5464 );
buf ( n14180 , n14179 );
not ( n14181 , n14180 );
buf ( n14182 , n5465 );
buf ( n14183 , n14182 );
not ( n14184 , n14183 );
buf ( n14185 , n5466 );
not ( n14186 , n14185 );
not ( n14187 , n14186 );
or ( n14188 , n14184 , n14187 );
not ( n14189 , n14182 );
buf ( n14190 , n14185 );
nand ( n14191 , n14189 , n14190 );
nand ( n14192 , n14188 , n14191 );
buf ( n14193 , n5467 );
buf ( n14194 , n14193 );
and ( n14195 , n14192 , n14194 );
not ( n14196 , n14192 );
not ( n14197 , n14193 );
and ( n14198 , n14196 , n14197 );
nor ( n14199 , n14195 , n14198 );
buf ( n14200 , n5468 );
nand ( n14201 , n7868 , n14200 );
buf ( n14202 , n5469 );
not ( n14203 , n14202 );
and ( n14204 , n14201 , n14203 );
not ( n14205 , n14201 );
buf ( n14206 , n14202 );
and ( n14207 , n14205 , n14206 );
nor ( n14208 , n14204 , n14207 );
xor ( n14209 , n14199 , n14208 );
buf ( n14210 , n5470 );
nand ( n14211 , n6973 , n14210 );
buf ( n14212 , n5471 );
not ( n14213 , n14212 );
and ( n14214 , n14211 , n14213 );
not ( n14215 , n14211 );
buf ( n14216 , n14212 );
and ( n14217 , n14215 , n14216 );
nor ( n14218 , n14214 , n14217 );
xnor ( n14219 , n14209 , n14218 );
not ( n14220 , n14219 );
not ( n14221 , n14220 );
not ( n14222 , n14221 );
or ( n14223 , n14181 , n14222 );
buf ( n14224 , n14219 );
not ( n14225 , n14224 );
not ( n14226 , n14179 );
nand ( n14227 , n14225 , n14226 );
nand ( n14228 , n14223 , n14227 );
buf ( n14229 , n5472 );
buf ( n14230 , n14229 );
not ( n14231 , n14230 );
buf ( n14232 , n5473 );
not ( n14233 , n14232 );
not ( n14234 , n14233 );
or ( n14235 , n14231 , n14234 );
not ( n14236 , n14229 );
buf ( n14237 , n14232 );
nand ( n14238 , n14236 , n14237 );
nand ( n14239 , n14235 , n14238 );
buf ( n14240 , n5474 );
not ( n14241 , n14240 );
and ( n14242 , n14239 , n14241 );
not ( n14243 , n14239 );
buf ( n14244 , n14240 );
and ( n14245 , n14243 , n14244 );
nor ( n14246 , n14242 , n14245 );
buf ( n14247 , n5475 );
nand ( n14248 , n7977 , n14247 );
buf ( n14249 , n5476 );
buf ( n14250 , n14249 );
and ( n14251 , n14248 , n14250 );
not ( n14252 , n14248 );
not ( n14253 , n14249 );
and ( n14254 , n14252 , n14253 );
nor ( n14255 , n14251 , n14254 );
xor ( n14256 , n14246 , n14255 );
buf ( n14257 , n5477 );
nand ( n14258 , n7258 , n14257 );
buf ( n14259 , n5478 );
buf ( n14260 , n14259 );
and ( n14261 , n14258 , n14260 );
not ( n14262 , n14258 );
not ( n14263 , n14259 );
and ( n14264 , n14262 , n14263 );
nor ( n14265 , n14261 , n14264 );
not ( n14266 , n14265 );
xnor ( n14267 , n14256 , n14266 );
buf ( n14268 , n14267 );
and ( n14269 , n14228 , n14268 );
not ( n14270 , n14228 );
xor ( n14271 , n14246 , n14265 );
xnor ( n14272 , n14271 , n14255 );
buf ( n14273 , n14272 );
and ( n14274 , n14270 , n14273 );
nor ( n14275 , n14269 , n14274 );
not ( n14276 , n11981 );
not ( n14277 , n10824 );
not ( n14278 , n14277 );
or ( n14279 , n14276 , n14278 );
not ( n14280 , n14277 );
nand ( n14281 , n14280 , n11977 );
nand ( n14282 , n14279 , n14281 );
buf ( n14283 , n5479 );
buf ( n14284 , n14283 );
not ( n14285 , n14284 );
buf ( n14286 , n5480 );
not ( n14287 , n14286 );
not ( n14288 , n14287 );
or ( n14289 , n14285 , n14288 );
not ( n14290 , n14283 );
buf ( n14291 , n14286 );
nand ( n14292 , n14290 , n14291 );
nand ( n14293 , n14289 , n14292 );
not ( n14294 , n12300 );
and ( n14295 , n14293 , n14294 );
not ( n14296 , n14293 );
and ( n14297 , n14296 , n12301 );
nor ( n14298 , n14295 , n14297 );
xor ( n14299 , n14298 , n13303 );
buf ( n14300 , n5481 );
nand ( n14301 , n8675 , n14300 );
buf ( n14302 , n5482 );
buf ( n14303 , n14302 );
and ( n14304 , n14301 , n14303 );
not ( n14305 , n14301 );
not ( n14306 , n14302 );
and ( n14307 , n14305 , n14306 );
nor ( n14308 , n14304 , n14307 );
xnor ( n14309 , n14299 , n14308 );
buf ( n14310 , n14309 );
not ( n14311 , n14310 );
buf ( n14312 , n14311 );
not ( n14313 , n14312 );
and ( n14314 , n14282 , n14313 );
not ( n14315 , n14282 );
and ( n14316 , n14315 , n14312 );
nor ( n14317 , n14314 , n14316 );
nand ( n14318 , n14275 , n14317 );
not ( n14319 , n14318 );
or ( n14320 , n14178 , n14319 );
nand ( n14321 , n14275 , n14317 );
or ( n14322 , n14321 , n14177 );
nand ( n14323 , n14320 , n14322 );
not ( n14324 , n14323 );
or ( n14325 , n14102 , n14324 );
or ( n14326 , n14323 , n14101 );
nand ( n14327 , n14325 , n14326 );
buf ( n14328 , n14327 );
xnor ( n14329 , n14007 , n14328 );
not ( n14330 , n14329 );
not ( n14331 , n14330 );
or ( n14332 , n13530 , n14331 );
xor ( n14333 , n14002 , n13855 );
xor ( n14334 , n14333 , n14327 );
not ( n14335 , n14334 );
or ( n14336 , n14335 , n13529 );
nand ( n14337 , n14332 , n14336 );
not ( n14338 , n14337 );
buf ( n14339 , n5483 );
buf ( n14340 , n5484 );
nand ( n14341 , n6827 , n14340 );
buf ( n14342 , n5485 );
buf ( n14343 , n14342 );
and ( n14344 , n14341 , n14343 );
not ( n14345 , n14341 );
not ( n14346 , n14342 );
and ( n14347 , n14345 , n14346 );
nor ( n14348 , n14344 , n14347 );
xor ( n14349 , n14339 , n14348 );
buf ( n14350 , n5486 );
nand ( n14351 , n6557 , n14350 );
buf ( n14352 , n5487 );
not ( n14353 , n14352 );
and ( n14354 , n14351 , n14353 );
not ( n14355 , n14351 );
buf ( n14356 , n14352 );
and ( n14357 , n14355 , n14356 );
nor ( n14358 , n14354 , n14357 );
xnor ( n14359 , n14349 , n14358 );
not ( n14360 , n14359 );
buf ( n14361 , n5488 );
not ( n14362 , n14361 );
buf ( n14363 , n5489 );
buf ( n14364 , n14363 );
and ( n14365 , n14362 , n14364 );
not ( n14366 , n14362 );
not ( n14367 , n14363 );
and ( n14368 , n14366 , n14367 );
nor ( n14369 , n14365 , n14368 );
not ( n14370 , n14369 );
and ( n14371 , n14360 , n14370 );
and ( n14372 , n14359 , n14369 );
nor ( n14373 , n14371 , n14372 );
not ( n14374 , n14373 );
xor ( n14375 , n7076 , n14374 );
buf ( n14376 , n5490 );
buf ( n14377 , n5491 );
not ( n14378 , n14377 );
buf ( n14379 , n5492 );
buf ( n14380 , n14379 );
nand ( n14381 , n14378 , n14380 );
not ( n14382 , n14379 );
buf ( n14383 , n14377 );
nand ( n14384 , n14382 , n14383 );
and ( n14385 , n14381 , n14384 );
xor ( n14386 , n14376 , n14385 );
buf ( n14387 , n5493 );
buf ( n14388 , n5494 );
xor ( n14389 , n14387 , n14388 );
buf ( n14390 , n5495 );
nand ( n14391 , n8223 , n14390 );
xnor ( n14392 , n14389 , n14391 );
xnor ( n14393 , n14386 , n14392 );
xor ( n14394 , n14375 , n14393 );
not ( n14395 , n9669 );
xor ( n14396 , n12789 , n12808 );
xor ( n14397 , n14396 , n12798 );
not ( n14398 , n14397 );
or ( n14399 , n14395 , n14398 );
or ( n14400 , n14397 , n9669 );
nand ( n14401 , n14399 , n14400 );
not ( n14402 , n6526 );
and ( n14403 , n14401 , n14402 );
not ( n14404 , n14401 );
buf ( n14405 , n6525 );
not ( n14406 , n14405 );
and ( n14407 , n14404 , n14406 );
nor ( n14408 , n14403 , n14407 );
nand ( n14409 , n14394 , n14408 );
not ( n14410 , n14409 );
buf ( n14411 , n5496 );
buf ( n14412 , n14411 );
not ( n14413 , n14412 );
buf ( n14414 , n5497 );
not ( n14415 , n14414 );
not ( n14416 , n14415 );
or ( n14417 , n14413 , n14416 );
not ( n14418 , n14411 );
buf ( n14419 , n14414 );
nand ( n14420 , n14418 , n14419 );
nand ( n14421 , n14417 , n14420 );
and ( n14422 , n14421 , n8146 );
not ( n14423 , n14421 );
not ( n14424 , n8145 );
and ( n14425 , n14423 , n14424 );
nor ( n14426 , n14422 , n14425 );
buf ( n14427 , n5498 );
nand ( n14428 , n6770 , n14427 );
buf ( n14429 , n5499 );
buf ( n14430 , n14429 );
and ( n14431 , n14428 , n14430 );
not ( n14432 , n14428 );
not ( n14433 , n14429 );
and ( n14434 , n14432 , n14433 );
nor ( n14435 , n14431 , n14434 );
xor ( n14436 , n14426 , n14435 );
buf ( n14437 , n5500 );
nand ( n14438 , n8032 , n14437 );
buf ( n14439 , n5501 );
not ( n14440 , n14439 );
and ( n14441 , n14438 , n14440 );
not ( n14442 , n14438 );
buf ( n14443 , n14439 );
and ( n14444 , n14442 , n14443 );
nor ( n14445 , n14441 , n14444 );
xnor ( n14446 , n14436 , n14445 );
not ( n14447 , n14446 );
not ( n14448 , n14447 );
not ( n14449 , n14448 );
not ( n14450 , n14449 );
not ( n14451 , n6899 );
not ( n14452 , n13132 );
or ( n14453 , n14451 , n14452 );
or ( n14454 , n13132 , n6899 );
nand ( n14455 , n14453 , n14454 );
not ( n14456 , n14455 );
or ( n14457 , n14450 , n14456 );
not ( n14458 , n14448 );
or ( n14459 , n14455 , n14458 );
nand ( n14460 , n14457 , n14459 );
not ( n14461 , n14460 );
and ( n14462 , n14410 , n14461 );
not ( n14463 , n14408 );
not ( n14464 , n14463 );
nand ( n14465 , n14464 , n14394 );
and ( n14466 , n14465 , n14460 );
nor ( n14467 , n14462 , n14466 );
not ( n14468 , n14467 );
buf ( n14469 , n5502 );
buf ( n14470 , n14469 );
not ( n14471 , n14470 );
buf ( n14472 , n5503 );
not ( n14473 , n14472 );
not ( n14474 , n14473 );
or ( n14475 , n14471 , n14474 );
not ( n14476 , n14469 );
buf ( n14477 , n14472 );
nand ( n14478 , n14476 , n14477 );
nand ( n14479 , n14475 , n14478 );
buf ( n14480 , n5504 );
buf ( n14481 , n14480 );
and ( n14482 , n14479 , n14481 );
not ( n14483 , n14479 );
not ( n14484 , n14480 );
and ( n14485 , n14483 , n14484 );
nor ( n14486 , n14482 , n14485 );
buf ( n14487 , n5505 );
nand ( n14488 , n7563 , n14487 );
buf ( n14489 , n5506 );
not ( n14490 , n14489 );
and ( n14491 , n14488 , n14490 );
not ( n14492 , n14488 );
buf ( n14493 , n14489 );
and ( n14494 , n14492 , n14493 );
nor ( n14495 , n14491 , n14494 );
xor ( n14496 , n14486 , n14495 );
buf ( n14497 , n5507 );
nand ( n14498 , n10383 , n14497 );
buf ( n14499 , n5508 );
not ( n14500 , n14499 );
and ( n14501 , n14498 , n14500 );
not ( n14502 , n14498 );
buf ( n14503 , n14499 );
and ( n14504 , n14502 , n14503 );
nor ( n14505 , n14501 , n14504 );
xnor ( n14506 , n14496 , n14505 );
not ( n14507 , n14506 );
buf ( n14508 , n14507 );
not ( n14509 , n14508 );
not ( n14510 , n14509 );
not ( n14511 , n7961 );
buf ( n14512 , n5509 );
buf ( n14513 , n14512 );
not ( n14514 , n14513 );
buf ( n14515 , n5510 );
not ( n14516 , n14515 );
not ( n14517 , n14516 );
or ( n14518 , n14514 , n14517 );
not ( n14519 , n14512 );
buf ( n14520 , n14515 );
nand ( n14521 , n14519 , n14520 );
nand ( n14522 , n14518 , n14521 );
buf ( n14523 , n5511 );
not ( n14524 , n14523 );
and ( n14525 , n14522 , n14524 );
not ( n14526 , n14522 );
buf ( n14527 , n14523 );
and ( n14528 , n14526 , n14527 );
nor ( n14529 , n14525 , n14528 );
xor ( n14530 , n14529 , n11969 );
buf ( n14531 , n5512 );
nand ( n14532 , n9310 , n14531 );
buf ( n14533 , n5513 );
buf ( n14534 , n14533 );
and ( n14535 , n14532 , n14534 );
not ( n14536 , n14532 );
not ( n14537 , n14533 );
and ( n14538 , n14536 , n14537 );
nor ( n14539 , n14535 , n14538 );
xnor ( n14540 , n14530 , n14539 );
buf ( n14541 , n14540 );
not ( n14542 , n14541 );
or ( n14543 , n14511 , n14542 );
not ( n14544 , n14540 );
buf ( n14545 , n7960 );
nand ( n14546 , n14544 , n14545 );
nand ( n14547 , n14543 , n14546 );
not ( n14548 , n14547 );
or ( n14549 , n14510 , n14548 );
or ( n14550 , n14547 , n14509 );
nand ( n14551 , n14549 , n14550 );
not ( n14552 , n14551 );
not ( n14553 , n8427 );
not ( n14554 , n14553 );
buf ( n14555 , n5514 );
not ( n14556 , n14555 );
buf ( n14557 , n5515 );
buf ( n14558 , n14557 );
not ( n14559 , n14558 );
buf ( n14560 , n5516 );
not ( n14561 , n14560 );
not ( n14562 , n14561 );
or ( n14563 , n14559 , n14562 );
not ( n14564 , n14557 );
buf ( n14565 , n14560 );
nand ( n14566 , n14564 , n14565 );
nand ( n14567 , n14563 , n14566 );
not ( n14568 , n14567 );
xor ( n14569 , n14556 , n14568 );
buf ( n14570 , n5517 );
buf ( n14571 , n5518 );
xor ( n14572 , n14570 , n14571 );
buf ( n14573 , n7293 );
buf ( n14574 , n5519 );
nand ( n14575 , n14573 , n14574 );
xnor ( n14576 , n14572 , n14575 );
xnor ( n14577 , n14569 , n14576 );
not ( n14578 , n14577 );
or ( n14579 , n14554 , n14578 );
not ( n14580 , n14553 );
not ( n14581 , n14577 );
nand ( n14582 , n14580 , n14581 );
nand ( n14583 , n14579 , n14582 );
buf ( n14584 , n5520 );
buf ( n14585 , n14584 );
not ( n14586 , n14585 );
buf ( n14587 , n5521 );
not ( n14588 , n14587 );
not ( n14589 , n14588 );
or ( n14590 , n14586 , n14589 );
not ( n14591 , n14584 );
buf ( n14592 , n14587 );
nand ( n14593 , n14591 , n14592 );
nand ( n14594 , n14590 , n14593 );
not ( n14595 , n14594 );
buf ( n14596 , n5522 );
not ( n14597 , n14596 );
buf ( n14598 , n5523 );
nand ( n14599 , n6633 , n14598 );
buf ( n14600 , n5524 );
buf ( n14601 , n14600 );
and ( n14602 , n14599 , n14601 );
not ( n14603 , n14599 );
not ( n14604 , n14600 );
and ( n14605 , n14603 , n14604 );
nor ( n14606 , n14602 , n14605 );
xor ( n14607 , n14597 , n14606 );
buf ( n14608 , n5525 );
nand ( n14609 , n7868 , n14608 );
buf ( n14610 , n5526 );
buf ( n14611 , n14610 );
and ( n14612 , n14609 , n14611 );
not ( n14613 , n14609 );
not ( n14614 , n14610 );
and ( n14615 , n14613 , n14614 );
nor ( n14616 , n14612 , n14615 );
xnor ( n14617 , n14607 , n14616 );
not ( n14618 , n14617 );
not ( n14619 , n14618 );
or ( n14620 , n14595 , n14619 );
not ( n14621 , n14594 );
nand ( n14622 , n14617 , n14621 );
nand ( n14623 , n14620 , n14622 );
buf ( n14624 , n14623 );
and ( n14625 , n14583 , n14624 );
not ( n14626 , n14583 );
not ( n14627 , n14624 );
and ( n14628 , n14626 , n14627 );
nor ( n14629 , n14625 , n14628 );
nand ( n14630 , n14552 , n14629 );
buf ( n14631 , n5527 );
buf ( n14632 , n5528 );
buf ( n14633 , n14632 );
not ( n14634 , n14633 );
buf ( n14635 , n5529 );
not ( n14636 , n14635 );
not ( n14637 , n14636 );
or ( n14638 , n14634 , n14637 );
not ( n14639 , n14632 );
buf ( n14640 , n14635 );
nand ( n14641 , n14639 , n14640 );
nand ( n14642 , n14638 , n14641 );
xor ( n14643 , n14631 , n14642 );
buf ( n14644 , n5530 );
buf ( n14645 , n5531 );
not ( n14646 , n14645 );
xor ( n14647 , n14644 , n14646 );
buf ( n14648 , n5532 );
nand ( n14649 , n8223 , n14648 );
xnor ( n14650 , n14647 , n14649 );
xnor ( n14651 , n14643 , n14650 );
not ( n14652 , n14651 );
not ( n14653 , n14652 );
not ( n14654 , n11242 );
buf ( n14655 , n5533 );
buf ( n14656 , n14655 );
not ( n14657 , n14656 );
buf ( n14658 , n5534 );
not ( n14659 , n14658 );
not ( n14660 , n14659 );
or ( n14661 , n14657 , n14660 );
not ( n14662 , n14655 );
buf ( n14663 , n14658 );
nand ( n14664 , n14662 , n14663 );
nand ( n14665 , n14661 , n14664 );
buf ( n14666 , n5535 );
buf ( n14667 , n14666 );
and ( n14668 , n14665 , n14667 );
not ( n14669 , n14665 );
not ( n14670 , n14666 );
and ( n14671 , n14669 , n14670 );
nor ( n14672 , n14668 , n14671 );
xor ( n14673 , n14672 , n11888 );
buf ( n14674 , n5536 );
nand ( n14675 , n11688 , n14674 );
buf ( n14676 , n5537 );
not ( n14677 , n14676 );
and ( n14678 , n14675 , n14677 );
not ( n14679 , n14675 );
buf ( n14680 , n14676 );
and ( n14681 , n14679 , n14680 );
nor ( n14682 , n14678 , n14681 );
xnor ( n14683 , n14673 , n14682 );
not ( n14684 , n14683 );
not ( n14685 , n14684 );
or ( n14686 , n14654 , n14685 );
nand ( n14687 , n14683 , n11238 );
nand ( n14688 , n14686 , n14687 );
not ( n14689 , n14688 );
and ( n14690 , n14653 , n14689 );
buf ( n14691 , n14651 );
not ( n14692 , n14691 );
and ( n14693 , n14692 , n14688 );
nor ( n14694 , n14690 , n14693 );
buf ( n14695 , n14694 );
and ( n14696 , n14630 , n14695 );
not ( n14697 , n14630 );
not ( n14698 , n14695 );
and ( n14699 , n14697 , n14698 );
nor ( n14700 , n14696 , n14699 );
not ( n14701 , n14700 );
or ( n14702 , n14468 , n14701 );
or ( n14703 , n14700 , n14467 );
nand ( n14704 , n14702 , n14703 );
buf ( n14705 , n5538 );
nand ( n14706 , n6502 , n14705 );
buf ( n14707 , n5539 );
not ( n14708 , n14707 );
and ( n14709 , n14706 , n14708 );
not ( n14710 , n14706 );
buf ( n14711 , n14707 );
and ( n14712 , n14710 , n14711 );
nor ( n14713 , n14709 , n14712 );
buf ( n14714 , n8398 );
xor ( n14715 , n14713 , n14714 );
buf ( n14716 , n5540 );
buf ( n14717 , n14716 );
not ( n14718 , n14717 );
buf ( n14719 , n5541 );
not ( n14720 , n14719 );
not ( n14721 , n14720 );
or ( n14722 , n14718 , n14721 );
not ( n14723 , n14716 );
buf ( n14724 , n14719 );
nand ( n14725 , n14723 , n14724 );
nand ( n14726 , n14722 , n14725 );
not ( n14727 , n14726 );
buf ( n14728 , n5542 );
buf ( n14729 , n14728 );
buf ( n14730 , n5543 );
nand ( n14731 , n8454 , n14730 );
buf ( n14732 , n5544 );
buf ( n14733 , n14732 );
and ( n14734 , n14731 , n14733 );
not ( n14735 , n14731 );
not ( n14736 , n14732 );
and ( n14737 , n14735 , n14736 );
nor ( n14738 , n14734 , n14737 );
xor ( n14739 , n14729 , n14738 );
buf ( n14740 , n5545 );
nand ( n14741 , n8032 , n14740 );
buf ( n14742 , n5546 );
not ( n14743 , n14742 );
and ( n14744 , n14741 , n14743 );
not ( n14745 , n14741 );
buf ( n14746 , n14742 );
and ( n14747 , n14745 , n14746 );
nor ( n14748 , n14744 , n14747 );
xnor ( n14749 , n14739 , n14748 );
and ( n14750 , n14727 , n14749 );
not ( n14751 , n14727 );
not ( n14752 , n14749 );
and ( n14753 , n14751 , n14752 );
nor ( n14754 , n14750 , n14753 );
buf ( n14755 , n14754 );
xnor ( n14756 , n14715 , n14755 );
buf ( n14757 , n13215 );
not ( n14758 , n14757 );
not ( n14759 , n13707 );
buf ( n14760 , n5547 );
not ( n14761 , n14760 );
not ( n14762 , n14761 );
or ( n14763 , n14759 , n14762 );
not ( n14764 , n13706 );
buf ( n14765 , n14760 );
nand ( n14766 , n14764 , n14765 );
nand ( n14767 , n14763 , n14766 );
not ( n14768 , n7426 );
and ( n14769 , n14767 , n14768 );
not ( n14770 , n14767 );
and ( n14771 , n14770 , n7427 );
nor ( n14772 , n14769 , n14771 );
buf ( n14773 , n5548 );
nand ( n14774 , n7202 , n14773 );
buf ( n14775 , n5549 );
buf ( n14776 , n14775 );
and ( n14777 , n14774 , n14776 );
not ( n14778 , n14774 );
not ( n14779 , n14775 );
and ( n14780 , n14778 , n14779 );
nor ( n14781 , n14777 , n14780 );
xor ( n14782 , n14772 , n14781 );
buf ( n14783 , n5550 );
nand ( n14784 , n9310 , n14783 );
buf ( n14785 , n5551 );
buf ( n14786 , n14785 );
and ( n14787 , n14784 , n14786 );
not ( n14788 , n14784 );
not ( n14789 , n14785 );
and ( n14790 , n14788 , n14789 );
nor ( n14791 , n14787 , n14790 );
xnor ( n14792 , n14782 , n14791 );
buf ( n14793 , n14792 );
not ( n14794 , n14793 );
not ( n14795 , n14794 );
or ( n14796 , n14758 , n14795 );
not ( n14797 , n14792 );
buf ( n14798 , n14797 );
not ( n14799 , n14798 );
not ( n14800 , n14799 );
or ( n14801 , n14800 , n14757 );
nand ( n14802 , n14796 , n14801 );
buf ( n14803 , n5552 );
buf ( n14804 , n14803 );
not ( n14805 , n14804 );
not ( n14806 , n12912 );
or ( n14807 , n14805 , n14806 );
not ( n14808 , n14803 );
buf ( n14809 , n12911 );
nand ( n14810 , n14808 , n14809 );
nand ( n14811 , n14807 , n14810 );
buf ( n14812 , n5553 );
buf ( n14813 , n14812 );
and ( n14814 , n14811 , n14813 );
not ( n14815 , n14811 );
not ( n14816 , n14812 );
and ( n14817 , n14815 , n14816 );
nor ( n14818 , n14814 , n14817 );
buf ( n14819 , n5554 );
nand ( n14820 , n6770 , n14819 );
buf ( n14821 , n5555 );
buf ( n14822 , n14821 );
and ( n14823 , n14820 , n14822 );
not ( n14824 , n14820 );
not ( n14825 , n14821 );
and ( n14826 , n14824 , n14825 );
nor ( n14827 , n14823 , n14826 );
xor ( n14828 , n14818 , n14827 );
buf ( n14829 , n5556 );
nand ( n14830 , n8608 , n14829 );
buf ( n14831 , n5557 );
not ( n14832 , n14831 );
and ( n14833 , n14830 , n14832 );
not ( n14834 , n14830 );
buf ( n14835 , n14831 );
and ( n14836 , n14834 , n14835 );
nor ( n14837 , n14833 , n14836 );
xnor ( n14838 , n14828 , n14837 );
not ( n14839 , n14838 );
not ( n14840 , n14839 );
and ( n14841 , n14802 , n14840 );
not ( n14842 , n14802 );
not ( n14843 , n14827 );
xor ( n14844 , n14818 , n14843 );
xnor ( n14845 , n14844 , n14837 );
not ( n14846 , n14845 );
not ( n14847 , n14846 );
and ( n14848 , n14842 , n14847 );
nor ( n14849 , n14841 , n14848 );
not ( n14850 , n14849 );
nand ( n14851 , n14756 , n14850 );
xor ( n14852 , n10355 , n11155 );
xnor ( n14853 , n14852 , n7833 );
and ( n14854 , n14851 , n14853 );
not ( n14855 , n14851 );
not ( n14856 , n14853 );
and ( n14857 , n14855 , n14856 );
nor ( n14858 , n14854 , n14857 );
not ( n14859 , n14858 );
and ( n14860 , n14704 , n14859 );
not ( n14861 , n14704 );
and ( n14862 , n14861 , n14858 );
nor ( n14863 , n14860 , n14862 );
not ( n14864 , n7513 );
buf ( n14865 , n5558 );
nand ( n14866 , n6646 , n14865 );
buf ( n14867 , n5559 );
buf ( n14868 , n14867 );
and ( n14869 , n14866 , n14868 );
not ( n14870 , n14866 );
not ( n14871 , n14867 );
and ( n14872 , n14870 , n14871 );
nor ( n14873 , n14869 , n14872 );
not ( n14874 , n14873 );
buf ( n14875 , n5560 );
nand ( n14876 , n6927 , n14875 );
buf ( n14877 , n5561 );
not ( n14878 , n14877 );
and ( n14879 , n14876 , n14878 );
not ( n14880 , n14876 );
buf ( n14881 , n14877 );
and ( n14882 , n14880 , n14881 );
nor ( n14883 , n14879 , n14882 );
not ( n14884 , n14883 );
or ( n14885 , n14874 , n14884 );
or ( n14886 , n14873 , n14883 );
nand ( n14887 , n14885 , n14886 );
buf ( n14888 , n5562 );
buf ( n14889 , n14888 );
not ( n14890 , n14889 );
buf ( n14891 , n5563 );
not ( n14892 , n14891 );
not ( n14893 , n14892 );
or ( n14894 , n14890 , n14893 );
not ( n14895 , n14888 );
buf ( n14896 , n14891 );
nand ( n14897 , n14895 , n14896 );
nand ( n14898 , n14894 , n14897 );
buf ( n14899 , n5564 );
not ( n14900 , n14899 );
and ( n14901 , n14898 , n14900 );
not ( n14902 , n14898 );
buf ( n14903 , n14899 );
and ( n14904 , n14902 , n14903 );
nor ( n14905 , n14901 , n14904 );
buf ( n14906 , n14905 );
and ( n14907 , n14887 , n14906 );
not ( n14908 , n14887 );
not ( n14909 , n14906 );
and ( n14910 , n14908 , n14909 );
nor ( n14911 , n14907 , n14910 );
not ( n14912 , n14911 );
not ( n14913 , n14912 );
not ( n14914 , n14913 );
or ( n14915 , n14864 , n14914 );
xor ( n14916 , n14905 , n14873 );
not ( n14917 , n14883 );
xnor ( n14918 , n14916 , n14917 );
not ( n14919 , n14918 );
not ( n14920 , n14919 );
nand ( n14921 , n14920 , n7516 );
nand ( n14922 , n14915 , n14921 );
buf ( n14923 , n5565 );
not ( n14924 , n14923 );
buf ( n14925 , n5566 );
not ( n14926 , n14925 );
buf ( n14927 , n5567 );
buf ( n14928 , n14927 );
nand ( n14929 , n14926 , n14928 );
not ( n14930 , n14927 );
buf ( n14931 , n14925 );
nand ( n14932 , n14930 , n14931 );
and ( n14933 , n14929 , n14932 );
xor ( n14934 , n14924 , n14933 );
buf ( n14935 , n5568 );
buf ( n14936 , n5569 );
not ( n14937 , n14936 );
xor ( n14938 , n14935 , n14937 );
buf ( n14939 , n5570 );
nand ( n14940 , n9310 , n14939 );
xnor ( n14941 , n14938 , n14940 );
xnor ( n14942 , n14934 , n14941 );
buf ( n14943 , n14942 );
and ( n14944 , n14922 , n14943 );
not ( n14945 , n14922 );
buf ( n14946 , n14923 );
xor ( n14947 , n14946 , n14933 );
xnor ( n14948 , n14947 , n14941 );
buf ( n14949 , n14948 );
and ( n14950 , n14945 , n14949 );
nor ( n14951 , n14944 , n14950 );
not ( n14952 , n14951 );
buf ( n14953 , n13041 );
not ( n14954 , n14953 );
buf ( n14955 , n5571 );
buf ( n14956 , n14955 );
not ( n14957 , n14956 );
buf ( n14958 , n5572 );
not ( n14959 , n14958 );
not ( n14960 , n14959 );
or ( n14961 , n14957 , n14960 );
not ( n14962 , n14955 );
buf ( n14963 , n14958 );
nand ( n14964 , n14962 , n14963 );
nand ( n14965 , n14961 , n14964 );
buf ( n14966 , n5573 );
buf ( n14967 , n14966 );
and ( n14968 , n14965 , n14967 );
not ( n14969 , n14965 );
not ( n14970 , n14966 );
and ( n14971 , n14969 , n14970 );
nor ( n14972 , n14968 , n14971 );
buf ( n14973 , n5574 );
nand ( n14974 , n8176 , n14973 );
buf ( n14975 , n5575 );
buf ( n14976 , n14975 );
and ( n14977 , n14974 , n14976 );
not ( n14978 , n14974 );
not ( n14979 , n14975 );
and ( n14980 , n14978 , n14979 );
nor ( n14981 , n14977 , n14980 );
xor ( n14982 , n14972 , n14981 );
buf ( n14983 , n5576 );
nand ( n14984 , n6816 , n14983 );
buf ( n14985 , n5577 );
not ( n14986 , n14985 );
and ( n14987 , n14984 , n14986 );
not ( n14988 , n14984 );
buf ( n14989 , n14985 );
and ( n14990 , n14988 , n14989 );
nor ( n14991 , n14987 , n14990 );
xnor ( n14992 , n14982 , n14991 );
not ( n14993 , n14992 );
not ( n14994 , n14993 );
or ( n14995 , n14954 , n14994 );
not ( n14996 , n14953 );
not ( n14997 , n14993 );
nand ( n14998 , n14996 , n14997 );
nand ( n14999 , n14995 , n14998 );
buf ( n15000 , n5578 );
nand ( n15001 , n7977 , n15000 );
buf ( n15002 , n5579 );
buf ( n15003 , n15002 );
and ( n15004 , n15001 , n15003 );
not ( n15005 , n15001 );
not ( n15006 , n15002 );
and ( n15007 , n15005 , n15006 );
nor ( n15008 , n15004 , n15007 );
not ( n15009 , n15008 );
buf ( n15010 , n5580 );
nand ( n15011 , n7868 , n15010 );
buf ( n15012 , n5581 );
not ( n15013 , n15012 );
and ( n15014 , n15011 , n15013 );
not ( n15015 , n15011 );
buf ( n15016 , n15012 );
and ( n15017 , n15015 , n15016 );
nor ( n15018 , n15014 , n15017 );
not ( n15019 , n15018 );
or ( n15020 , n15009 , n15019 );
or ( n15021 , n15008 , n15018 );
nand ( n15022 , n15020 , n15021 );
buf ( n15023 , n5582 );
buf ( n15024 , n15023 );
not ( n15025 , n15024 );
buf ( n15026 , n5583 );
not ( n15027 , n15026 );
not ( n15028 , n15027 );
or ( n15029 , n15025 , n15028 );
not ( n15030 , n15023 );
buf ( n15031 , n15026 );
nand ( n15032 , n15030 , n15031 );
nand ( n15033 , n15029 , n15032 );
buf ( n15034 , n5584 );
not ( n15035 , n15034 );
and ( n15036 , n15033 , n15035 );
not ( n15037 , n15033 );
buf ( n15038 , n15034 );
and ( n15039 , n15037 , n15038 );
nor ( n15040 , n15036 , n15039 );
and ( n15041 , n15022 , n15040 );
not ( n15042 , n15022 );
not ( n15043 , n15040 );
and ( n15044 , n15042 , n15043 );
nor ( n15045 , n15041 , n15044 );
buf ( n15046 , n15045 );
buf ( n15047 , n15046 );
and ( n15048 , n14999 , n15047 );
not ( n15049 , n14999 );
not ( n15050 , n15008 );
xor ( n15051 , n15040 , n15050 );
xnor ( n15052 , n15051 , n15018 );
buf ( n15053 , n15052 );
not ( n15054 , n15053 );
not ( n15055 , n15054 );
and ( n15056 , n15049 , n15055 );
nor ( n15057 , n15048 , n15056 );
not ( n15058 , n15057 );
nand ( n15059 , n14952 , n15058 );
not ( n15060 , n12304 );
buf ( n15061 , n5585 );
buf ( n15062 , n15061 );
not ( n15063 , n15062 );
buf ( n15064 , n5586 );
not ( n15065 , n15064 );
not ( n15066 , n15065 );
or ( n15067 , n15063 , n15066 );
not ( n15068 , n15061 );
buf ( n15069 , n15064 );
nand ( n15070 , n15068 , n15069 );
nand ( n15071 , n15067 , n15070 );
buf ( n15072 , n5587 );
buf ( n15073 , n15072 );
and ( n15074 , n15071 , n15073 );
not ( n15075 , n15071 );
not ( n15076 , n15072 );
and ( n15077 , n15075 , n15076 );
nor ( n15078 , n15074 , n15077 );
buf ( n15079 , n5588 );
nand ( n15080 , n7014 , n15079 );
buf ( n15081 , n5589 );
buf ( n15082 , n15081 );
and ( n15083 , n15080 , n15082 );
not ( n15084 , n15080 );
not ( n15085 , n15081 );
and ( n15086 , n15084 , n15085 );
nor ( n15087 , n15083 , n15086 );
xor ( n15088 , n15078 , n15087 );
buf ( n15089 , n5590 );
nand ( n15090 , n10874 , n15089 );
buf ( n15091 , n5591 );
buf ( n15092 , n15091 );
and ( n15093 , n15090 , n15092 );
not ( n15094 , n15090 );
not ( n15095 , n15091 );
and ( n15096 , n15094 , n15095 );
nor ( n15097 , n15093 , n15096 );
xnor ( n15098 , n15088 , n15097 );
buf ( n15099 , n15098 );
buf ( n15100 , n15099 );
not ( n15101 , n15100 );
or ( n15102 , n15060 , n15101 );
or ( n15103 , n15100 , n12304 );
nand ( n15104 , n15102 , n15103 );
not ( n15105 , n10535 );
not ( n15106 , n15105 );
and ( n15107 , n15104 , n15106 );
not ( n15108 , n15104 );
and ( n15109 , n15108 , n15105 );
nor ( n15110 , n15107 , n15109 );
buf ( n15111 , n15110 );
xor ( n15112 , n15059 , n15111 );
not ( n15113 , n15112 );
buf ( n15114 , n5592 );
not ( n15115 , n15114 );
not ( n15116 , n15115 );
buf ( n15117 , n5593 );
buf ( n15118 , n5594 );
not ( n15119 , n15118 );
buf ( n15120 , n5595 );
buf ( n15121 , n15120 );
and ( n15122 , n15119 , n15121 );
not ( n15123 , n15119 );
not ( n15124 , n15120 );
and ( n15125 , n15123 , n15124 );
nor ( n15126 , n15122 , n15125 );
xor ( n15127 , n15117 , n15126 );
buf ( n15128 , n5596 );
nand ( n15129 , n6770 , n15128 );
not ( n15130 , n15129 );
buf ( n15131 , n5597 );
not ( n15132 , n15131 );
and ( n15133 , n15130 , n15132 );
nand ( n15134 , n6515 , n15128 );
and ( n15135 , n15134 , n15131 );
nor ( n15136 , n15133 , n15135 );
not ( n15137 , n15136 );
buf ( n15138 , n5598 );
not ( n15139 , n15138 );
and ( n15140 , n15137 , n15139 );
and ( n15141 , n15136 , n15138 );
nor ( n15142 , n15140 , n15141 );
xnor ( n15143 , n15127 , n15142 );
buf ( n15144 , n15143 );
not ( n15145 , n15144 );
not ( n15146 , n15145 );
or ( n15147 , n15116 , n15146 );
not ( n15148 , n15144 );
or ( n15149 , n15148 , n15115 );
nand ( n15150 , n15147 , n15149 );
buf ( n15151 , n5599 );
not ( n15152 , n15151 );
not ( n15153 , n15152 );
buf ( n15154 , n5600 );
not ( n15155 , n15154 );
and ( n15156 , n15153 , n15155 );
and ( n15157 , n15154 , n15152 );
nor ( n15158 , n15156 , n15157 );
not ( n15159 , n15158 );
not ( n15160 , n15159 );
buf ( n15161 , n5601 );
not ( n15162 , n15161 );
buf ( n15163 , n5602 );
nand ( n15164 , n6502 , n15163 );
buf ( n15165 , n5603 );
buf ( n15166 , n15165 );
and ( n15167 , n15164 , n15166 );
not ( n15168 , n15164 );
not ( n15169 , n15165 );
and ( n15170 , n15168 , n15169 );
nor ( n15171 , n15167 , n15170 );
xor ( n15172 , n15162 , n15171 );
buf ( n15173 , n5604 );
nand ( n15174 , n8966 , n15173 );
buf ( n15175 , n5605 );
buf ( n15176 , n15175 );
and ( n15177 , n15174 , n15176 );
not ( n15178 , n15174 );
not ( n15179 , n15175 );
and ( n15180 , n15178 , n15179 );
nor ( n15181 , n15177 , n15180 );
xnor ( n15182 , n15172 , n15181 );
not ( n15183 , n15182 );
not ( n15184 , n15183 );
or ( n15185 , n15160 , n15184 );
nand ( n15186 , n15182 , n15158 );
nand ( n15187 , n15185 , n15186 );
and ( n15188 , n15150 , n15187 );
not ( n15189 , n15150 );
not ( n15190 , n15187 );
and ( n15191 , n15189 , n15190 );
nor ( n15192 , n15188 , n15191 );
not ( n15193 , n15192 );
buf ( n15194 , n14616 );
not ( n15195 , n15194 );
not ( n15196 , n15195 );
not ( n15197 , n13257 );
buf ( n15198 , n5606 );
not ( n15199 , n15198 );
not ( n15200 , n15199 );
or ( n15201 , n15197 , n15200 );
not ( n15202 , n13256 );
buf ( n15203 , n15198 );
nand ( n15204 , n15202 , n15203 );
nand ( n15205 , n15201 , n15204 );
buf ( n15206 , n5607 );
buf ( n15207 , n15206 );
and ( n15208 , n15205 , n15207 );
not ( n15209 , n15205 );
not ( n15210 , n15206 );
and ( n15211 , n15209 , n15210 );
nor ( n15212 , n15208 , n15211 );
buf ( n15213 , n5608 );
nand ( n15214 , n6770 , n15213 );
buf ( n15215 , n5609 );
buf ( n15216 , n15215 );
and ( n15217 , n15214 , n15216 );
not ( n15218 , n15214 );
not ( n15219 , n15215 );
and ( n15220 , n15218 , n15219 );
nor ( n15221 , n15217 , n15220 );
xor ( n15222 , n15212 , n15221 );
buf ( n15223 , n5610 );
nand ( n15224 , n6634 , n15223 );
buf ( n15225 , n5611 );
not ( n15226 , n15225 );
and ( n15227 , n15224 , n15226 );
not ( n15228 , n15224 );
buf ( n15229 , n15225 );
and ( n15230 , n15228 , n15229 );
nor ( n15231 , n15227 , n15230 );
xnor ( n15232 , n15222 , n15231 );
not ( n15233 , n15232 );
buf ( n15234 , n15233 );
not ( n15235 , n15234 );
or ( n15236 , n15196 , n15235 );
buf ( n15237 , n15232 );
nand ( n15238 , n15237 , n15194 );
nand ( n15239 , n15236 , n15238 );
not ( n15240 , n10749 );
not ( n15241 , n15240 );
buf ( n15242 , n15241 );
and ( n15243 , n15239 , n15242 );
not ( n15244 , n15239 );
buf ( n15245 , n10744 );
and ( n15246 , n15244 , n15245 );
nor ( n15247 , n15243 , n15246 );
nand ( n15248 , n15193 , n15247 );
not ( n15249 , n15248 );
buf ( n15250 , n5612 );
buf ( n15251 , n15250 );
not ( n15252 , n15251 );
buf ( n15253 , n5613 );
buf ( n15254 , n15253 );
not ( n15255 , n15254 );
buf ( n15256 , n5614 );
not ( n15257 , n15256 );
not ( n15258 , n15257 );
or ( n15259 , n15255 , n15258 );
not ( n15260 , n15253 );
buf ( n15261 , n15256 );
nand ( n15262 , n15260 , n15261 );
nand ( n15263 , n15259 , n15262 );
buf ( n15264 , n5615 );
buf ( n15265 , n15264 );
and ( n15266 , n15263 , n15265 );
not ( n15267 , n15263 );
not ( n15268 , n15264 );
and ( n15269 , n15267 , n15268 );
nor ( n15270 , n15266 , n15269 );
buf ( n15271 , n5616 );
nand ( n15272 , n6557 , n15271 );
buf ( n15273 , n5617 );
not ( n15274 , n15273 );
and ( n15275 , n15272 , n15274 );
not ( n15276 , n15272 );
buf ( n15277 , n15273 );
and ( n15278 , n15276 , n15277 );
nor ( n15279 , n15275 , n15278 );
xor ( n15280 , n15270 , n15279 );
buf ( n15281 , n5618 );
nand ( n15282 , n8223 , n15281 );
buf ( n15283 , n5619 );
not ( n15284 , n15283 );
and ( n15285 , n15282 , n15284 );
not ( n15286 , n15282 );
buf ( n15287 , n15283 );
and ( n15288 , n15286 , n15287 );
nor ( n15289 , n15285 , n15288 );
xnor ( n15290 , n15280 , n15289 );
buf ( n15291 , n15290 );
not ( n15292 , n15291 );
or ( n15293 , n15252 , n15292 );
or ( n15294 , n15291 , n15251 );
nand ( n15295 , n15293 , n15294 );
not ( n15296 , n15295 );
not ( n15297 , n14224 );
not ( n15298 , n15297 );
not ( n15299 , n15298 );
and ( n15300 , n15296 , n15299 );
and ( n15301 , n15295 , n14221 );
nor ( n15302 , n15300 , n15301 );
not ( n15303 , n15302 );
not ( n15304 , n15303 );
and ( n15305 , n15249 , n15304 );
and ( n15306 , n15248 , n15303 );
nor ( n15307 , n15305 , n15306 );
not ( n15308 , n15307 );
or ( n15309 , n15113 , n15308 );
not ( n15310 , n15112 );
not ( n15311 , n15307 );
nand ( n15312 , n15310 , n15311 );
nand ( n15313 , n15309 , n15312 );
and ( n15314 , n14863 , n15313 );
not ( n15315 , n14863 );
not ( n15316 , n15313 );
and ( n15317 , n15315 , n15316 );
nor ( n15318 , n15314 , n15317 );
buf ( n15319 , n15318 );
not ( n15320 , n15319 );
and ( n15321 , n14338 , n15320 );
and ( n15322 , n14337 , n15319 );
nor ( n15323 , n15321 , n15322 );
buf ( n15324 , n13344 );
buf ( n15325 , n15324 );
buf ( n15326 , n15325 );
not ( n15327 , n15326 );
nand ( n15328 , n15323 , n15327 );
buf ( n15329 , n5620 );
buf ( n15330 , n15329 );
not ( n15331 , n15330 );
buf ( n15332 , n5621 );
not ( n15333 , n15332 );
not ( n15334 , n15333 );
or ( n15335 , n15331 , n15334 );
not ( n15336 , n15329 );
buf ( n15337 , n15332 );
nand ( n15338 , n15336 , n15337 );
nand ( n15339 , n15335 , n15338 );
buf ( n15340 , n15339 );
not ( n15341 , n15340 );
buf ( n15342 , n5622 );
buf ( n15343 , n5623 );
not ( n15344 , n15343 );
xor ( n15345 , n15342 , n15344 );
buf ( n15346 , n5624 );
nand ( n15347 , n7247 , n15346 );
buf ( n15348 , n5625 );
not ( n15349 , n15348 );
and ( n15350 , n15347 , n15349 );
not ( n15351 , n15347 );
buf ( n15352 , n15348 );
and ( n15353 , n15351 , n15352 );
nor ( n15354 , n15350 , n15353 );
xnor ( n15355 , n15345 , n15354 );
not ( n15356 , n15355 );
not ( n15357 , n15356 );
or ( n15358 , n15341 , n15357 );
not ( n15359 , n15340 );
nand ( n15360 , n15359 , n15355 );
nand ( n15361 , n15358 , n15360 );
not ( n15362 , n15361 );
not ( n15363 , n11500 );
buf ( n15364 , n5626 );
nand ( n15365 , n6557 , n15364 );
buf ( n15366 , n5627 );
buf ( n15367 , n15366 );
and ( n15368 , n15365 , n15367 );
not ( n15369 , n15365 );
not ( n15370 , n15366 );
and ( n15371 , n15369 , n15370 );
nor ( n15372 , n15368 , n15371 );
buf ( n15373 , n15372 );
not ( n15374 , n15373 );
and ( n15375 , n15363 , n15374 );
not ( n15376 , n11501 );
and ( n15377 , n15376 , n15373 );
nor ( n15378 , n15375 , n15377 );
not ( n15379 , n15378 );
and ( n15380 , n15362 , n15379 );
buf ( n15381 , n15361 );
and ( n15382 , n15381 , n15378 );
nor ( n15383 , n15380 , n15382 );
not ( n15384 , n15383 );
not ( n15385 , n10087 );
buf ( n15386 , n5628 );
buf ( n15387 , n15386 );
not ( n15388 , n15387 );
buf ( n15389 , n5629 );
not ( n15390 , n15389 );
not ( n15391 , n15390 );
or ( n15392 , n15388 , n15391 );
not ( n15393 , n15386 );
buf ( n15394 , n15389 );
nand ( n15395 , n15393 , n15394 );
nand ( n15396 , n15392 , n15395 );
buf ( n15397 , n5630 );
not ( n15398 , n15397 );
and ( n15399 , n15396 , n15398 );
not ( n15400 , n15396 );
buf ( n15401 , n15397 );
and ( n15402 , n15400 , n15401 );
nor ( n15403 , n15399 , n15402 );
buf ( n15404 , n5631 );
nand ( n15405 , n6502 , n15404 );
buf ( n15406 , n5632 );
buf ( n15407 , n15406 );
and ( n15408 , n15405 , n15407 );
not ( n15409 , n15405 );
not ( n15410 , n15406 );
and ( n15411 , n15409 , n15410 );
nor ( n15412 , n15408 , n15411 );
xor ( n15413 , n15403 , n15412 );
buf ( n15414 , n5633 );
nand ( n15415 , n6647 , n15414 );
buf ( n15416 , n5634 );
not ( n15417 , n15416 );
and ( n15418 , n15415 , n15417 );
not ( n15419 , n15415 );
buf ( n15420 , n15416 );
and ( n15421 , n15419 , n15420 );
nor ( n15422 , n15418 , n15421 );
xor ( n15423 , n15413 , n15422 );
not ( n15424 , n15423 );
not ( n15425 , n15424 );
or ( n15426 , n15385 , n15425 );
not ( n15427 , n10087 );
not ( n15428 , n15423 );
not ( n15429 , n15428 );
nand ( n15430 , n15427 , n15429 );
nand ( n15431 , n15426 , n15430 );
buf ( n15432 , n5635 );
buf ( n15433 , n15432 );
not ( n15434 , n15433 );
buf ( n15435 , n5636 );
not ( n15436 , n15435 );
not ( n15437 , n15436 );
or ( n15438 , n15434 , n15437 );
not ( n15439 , n15432 );
buf ( n15440 , n15435 );
nand ( n15441 , n15439 , n15440 );
nand ( n15442 , n15438 , n15441 );
buf ( n15443 , n5637 );
buf ( n15444 , n15443 );
and ( n15445 , n15442 , n15444 );
not ( n15446 , n15442 );
not ( n15447 , n15443 );
and ( n15448 , n15446 , n15447 );
nor ( n15449 , n15445 , n15448 );
buf ( n15450 , n5638 );
nand ( n15451 , n9812 , n15450 );
buf ( n15452 , n5639 );
buf ( n15453 , n15452 );
and ( n15454 , n15451 , n15453 );
not ( n15455 , n15451 );
not ( n15456 , n15452 );
and ( n15457 , n15455 , n15456 );
nor ( n15458 , n15454 , n15457 );
xor ( n15459 , n15449 , n15458 );
buf ( n15460 , n5640 );
nand ( n15461 , n10947 , n15460 );
buf ( n15462 , n5641 );
not ( n15463 , n15462 );
and ( n15464 , n15461 , n15463 );
not ( n15465 , n15461 );
buf ( n15466 , n15462 );
and ( n15467 , n15465 , n15466 );
nor ( n15468 , n15464 , n15467 );
xor ( n15469 , n15459 , n15468 );
buf ( n15470 , n15469 );
not ( n15471 , n15470 );
and ( n15472 , n15431 , n15471 );
not ( n15473 , n15431 );
not ( n15474 , n15469 );
not ( n15475 , n15474 );
and ( n15476 , n15473 , n15475 );
nor ( n15477 , n15472 , n15476 );
not ( n15478 , n15477 );
nand ( n15479 , n15384 , n15478 );
buf ( n15480 , n5642 );
buf ( n15481 , n15480 );
not ( n15482 , n15481 );
buf ( n15483 , n5643 );
not ( n15484 , n15483 );
not ( n15485 , n15484 );
or ( n15486 , n15482 , n15485 );
not ( n15487 , n15480 );
buf ( n15488 , n15483 );
nand ( n15489 , n15487 , n15488 );
nand ( n15490 , n15486 , n15489 );
buf ( n15491 , n5644 );
not ( n15492 , n15491 );
and ( n15493 , n15490 , n15492 );
not ( n15494 , n15490 );
buf ( n15495 , n15491 );
and ( n15496 , n15494 , n15495 );
nor ( n15497 , n15493 , n15496 );
buf ( n15498 , n5645 );
nand ( n15499 , n8124 , n15498 );
buf ( n15500 , n5646 );
buf ( n15501 , n15500 );
and ( n15502 , n15499 , n15501 );
not ( n15503 , n15499 );
not ( n15504 , n15500 );
and ( n15505 , n15503 , n15504 );
nor ( n15506 , n15502 , n15505 );
xor ( n15507 , n15497 , n15506 );
buf ( n15508 , n5647 );
nand ( n15509 , n6816 , n15508 );
buf ( n15510 , n5648 );
buf ( n15511 , n15510 );
and ( n15512 , n15509 , n15511 );
not ( n15513 , n15509 );
not ( n15514 , n15510 );
and ( n15515 , n15513 , n15514 );
nor ( n15516 , n15512 , n15515 );
xnor ( n15517 , n15507 , n15516 );
not ( n15518 , n15517 );
nor ( n15519 , n15518 , n14125 );
not ( n15520 , n15519 );
buf ( n15521 , n15517 );
not ( n15522 , n15521 );
nand ( n15523 , n15522 , n14125 );
nand ( n15524 , n15520 , n15523 );
buf ( n15525 , n5649 );
buf ( n15526 , n15525 );
not ( n15527 , n15526 );
buf ( n15528 , n5650 );
not ( n15529 , n15528 );
not ( n15530 , n15529 );
or ( n15531 , n15527 , n15530 );
not ( n15532 , n15525 );
buf ( n15533 , n15528 );
nand ( n15534 , n15532 , n15533 );
nand ( n15535 , n15531 , n15534 );
not ( n15536 , n9096 );
and ( n15537 , n15535 , n15536 );
not ( n15538 , n15535 );
and ( n15539 , n15538 , n9097 );
nor ( n15540 , n15537 , n15539 );
buf ( n15541 , n5651 );
nand ( n15542 , n7698 , n15541 );
buf ( n15543 , n5652 );
not ( n15544 , n15543 );
and ( n15545 , n15542 , n15544 );
not ( n15546 , n15542 );
buf ( n15547 , n15543 );
and ( n15548 , n15546 , n15547 );
nor ( n15549 , n15545 , n15548 );
not ( n15550 , n15549 );
xor ( n15551 , n15540 , n15550 );
buf ( n15552 , n5653 );
nand ( n15553 , n6557 , n15552 );
buf ( n15554 , n5654 );
buf ( n15555 , n15554 );
and ( n15556 , n15553 , n15555 );
not ( n15557 , n15553 );
not ( n15558 , n15554 );
and ( n15559 , n15557 , n15558 );
nor ( n15560 , n15556 , n15559 );
buf ( n15561 , n15560 );
xnor ( n15562 , n15551 , n15561 );
buf ( n15563 , n15562 );
and ( n15564 , n15524 , n15563 );
not ( n15565 , n15524 );
not ( n15566 , n15560 );
not ( n15567 , n15549 );
or ( n15568 , n15566 , n15567 );
or ( n15569 , n15560 , n15549 );
nand ( n15570 , n15568 , n15569 );
and ( n15571 , n15570 , n15540 );
not ( n15572 , n15570 );
not ( n15573 , n15540 );
and ( n15574 , n15572 , n15573 );
nor ( n15575 , n15571 , n15574 );
buf ( n15576 , n15575 );
and ( n15577 , n15565 , n15576 );
nor ( n15578 , n15564 , n15577 );
not ( n15579 , n15578 );
and ( n15580 , n15479 , n15579 );
not ( n15581 , n15479 );
and ( n15582 , n15581 , n15578 );
nor ( n15583 , n15580 , n15582 );
not ( n15584 , n15583 );
buf ( n15585 , n5655 );
buf ( n15586 , n15585 );
not ( n15587 , n15586 );
not ( n15588 , n13203 );
not ( n15589 , n15588 );
or ( n15590 , n15587 , n15589 );
not ( n15591 , n15585 );
nand ( n15592 , n15591 , n13204 );
nand ( n15593 , n15590 , n15592 );
xor ( n15594 , n8344 , n15593 );
buf ( n15595 , n5656 );
buf ( n15596 , n5657 );
not ( n15597 , n15596 );
xor ( n15598 , n15595 , n15597 );
buf ( n15599 , n5658 );
nand ( n15600 , n8675 , n15599 );
xnor ( n15601 , n15598 , n15600 );
xnor ( n15602 , n15594 , n15601 );
not ( n15603 , n15602 );
not ( n15604 , n15603 );
buf ( n15605 , n5659 );
buf ( n15606 , n15605 );
not ( n15607 , n15606 );
buf ( n15608 , n5660 );
not ( n15609 , n15608 );
not ( n15610 , n15609 );
or ( n15611 , n15607 , n15610 );
not ( n15612 , n15605 );
buf ( n15613 , n15608 );
nand ( n15614 , n15612 , n15613 );
nand ( n15615 , n15611 , n15614 );
buf ( n15616 , n5661 );
buf ( n15617 , n15616 );
and ( n15618 , n15615 , n15617 );
not ( n15619 , n15615 );
not ( n15620 , n15616 );
and ( n15621 , n15619 , n15620 );
nor ( n15622 , n15618 , n15621 );
xor ( n15623 , n15622 , n14713 );
buf ( n15624 , n5662 );
nand ( n15625 , n14573 , n15624 );
buf ( n15626 , n5663 );
not ( n15627 , n15626 );
and ( n15628 , n15625 , n15627 );
not ( n15629 , n15625 );
buf ( n15630 , n15626 );
and ( n15631 , n15629 , n15630 );
nor ( n15632 , n15628 , n15631 );
xnor ( n15633 , n15623 , n15632 );
not ( n15634 , n15633 );
not ( n15635 , n15634 );
buf ( n15636 , n6524 );
not ( n15637 , n15636 );
and ( n15638 , n15635 , n15637 );
not ( n15639 , n15633 );
and ( n15640 , n15639 , n15636 );
nor ( n15641 , n15638 , n15640 );
xor ( n15642 , n15604 , n15641 );
not ( n15643 , n15642 );
buf ( n15644 , n5664 );
buf ( n15645 , n15644 );
not ( n15646 , n15645 );
buf ( n15647 , n5665 );
buf ( n15648 , n15647 );
not ( n15649 , n15648 );
buf ( n15650 , n5666 );
not ( n15651 , n15650 );
not ( n15652 , n15651 );
or ( n15653 , n15649 , n15652 );
not ( n15654 , n15647 );
buf ( n15655 , n15650 );
nand ( n15656 , n15654 , n15655 );
nand ( n15657 , n15653 , n15656 );
buf ( n15658 , n5667 );
not ( n15659 , n15658 );
and ( n15660 , n15657 , n15659 );
not ( n15661 , n15657 );
buf ( n15662 , n15658 );
and ( n15663 , n15661 , n15662 );
nor ( n15664 , n15660 , n15663 );
buf ( n15665 , n5668 );
nand ( n15666 , n10165 , n15665 );
buf ( n15667 , n5669 );
buf ( n15668 , n15667 );
and ( n15669 , n15666 , n15668 );
not ( n15670 , n15666 );
not ( n15671 , n15667 );
and ( n15672 , n15670 , n15671 );
nor ( n15673 , n15669 , n15672 );
xor ( n15674 , n15664 , n15673 );
buf ( n15675 , n5670 );
nand ( n15676 , n8323 , n15675 );
buf ( n15677 , n5671 );
buf ( n15678 , n15677 );
and ( n15679 , n15676 , n15678 );
not ( n15680 , n15676 );
not ( n15681 , n15677 );
and ( n15682 , n15680 , n15681 );
nor ( n15683 , n15679 , n15682 );
not ( n15684 , n15683 );
xnor ( n15685 , n15674 , n15684 );
not ( n15686 , n15685 );
or ( n15687 , n15646 , n15686 );
not ( n15688 , n15645 );
not ( n15689 , n15685 );
nand ( n15690 , n15688 , n15689 );
nand ( n15691 , n15687 , n15690 );
not ( n15692 , n12498 );
and ( n15693 , n15691 , n15692 );
not ( n15694 , n15691 );
and ( n15695 , n15694 , n12498 );
nor ( n15696 , n15693 , n15695 );
not ( n15697 , n15696 );
nand ( n15698 , n15643 , n15697 );
not ( n15699 , n15698 );
not ( n15700 , n15062 );
buf ( n15701 , n14506 );
not ( n15702 , n15701 );
or ( n15703 , n15700 , n15702 );
not ( n15704 , n14507 );
or ( n15705 , n15704 , n15062 );
nand ( n15706 , n15703 , n15705 );
buf ( n15707 , n5672 );
buf ( n15708 , n15707 );
not ( n15709 , n15708 );
buf ( n15710 , n5673 );
not ( n15711 , n15710 );
not ( n15712 , n15711 );
or ( n15713 , n15709 , n15712 );
not ( n15714 , n15707 );
buf ( n15715 , n15710 );
nand ( n15716 , n15714 , n15715 );
nand ( n15717 , n15713 , n15716 );
buf ( n15718 , n5674 );
not ( n15719 , n15718 );
and ( n15720 , n15717 , n15719 );
not ( n15721 , n15717 );
buf ( n15722 , n15718 );
and ( n15723 , n15721 , n15722 );
nor ( n15724 , n15720 , n15723 );
buf ( n15725 , n5675 );
nand ( n15726 , n6604 , n15725 );
buf ( n15727 , n5676 );
not ( n15728 , n15727 );
and ( n15729 , n15726 , n15728 );
not ( n15730 , n15726 );
buf ( n15731 , n15727 );
and ( n15732 , n15730 , n15731 );
nor ( n15733 , n15729 , n15732 );
xor ( n15734 , n15724 , n15733 );
buf ( n15735 , n5677 );
nand ( n15736 , n7258 , n15735 );
buf ( n15737 , n5678 );
buf ( n15738 , n15737 );
and ( n15739 , n15736 , n15738 );
not ( n15740 , n15736 );
not ( n15741 , n15737 );
and ( n15742 , n15740 , n15741 );
nor ( n15743 , n15739 , n15742 );
xor ( n15744 , n15734 , n15743 );
not ( n15745 , n15744 );
and ( n15746 , n15706 , n15745 );
not ( n15747 , n15706 );
not ( n15748 , n15744 );
not ( n15749 , n15748 );
not ( n15750 , n15749 );
not ( n15751 , n15750 );
and ( n15752 , n15747 , n15751 );
nor ( n15753 , n15746 , n15752 );
not ( n15754 , n15753 );
not ( n15755 , n15754 );
and ( n15756 , n15699 , n15755 );
and ( n15757 , n15698 , n15754 );
nor ( n15758 , n15756 , n15757 );
not ( n15759 , n15758 );
buf ( n15760 , n12712 );
not ( n15761 , n15760 );
buf ( n15762 , n5679 );
not ( n15763 , n15762 );
buf ( n15764 , n5680 );
buf ( n15765 , n15764 );
not ( n15766 , n15765 );
buf ( n15767 , n5681 );
not ( n15768 , n15767 );
not ( n15769 , n15768 );
or ( n15770 , n15766 , n15769 );
not ( n15771 , n15764 );
buf ( n15772 , n15767 );
nand ( n15773 , n15771 , n15772 );
nand ( n15774 , n15770 , n15773 );
xor ( n15775 , n15763 , n15774 );
buf ( n15776 , n5682 );
nand ( n15777 , n7606 , n15776 );
buf ( n15778 , n5683 );
buf ( n15779 , n15778 );
and ( n15780 , n15777 , n15779 );
not ( n15781 , n15777 );
not ( n15782 , n15778 );
and ( n15783 , n15781 , n15782 );
nor ( n15784 , n15780 , n15783 );
not ( n15785 , n15784 );
buf ( n15786 , n5684 );
not ( n15787 , n15786 );
and ( n15788 , n15785 , n15787 );
and ( n15789 , n15784 , n15786 );
nor ( n15790 , n15788 , n15789 );
xnor ( n15791 , n15775 , n15790 );
not ( n15792 , n15791 );
or ( n15793 , n15761 , n15792 );
or ( n15794 , n15791 , n15760 );
nand ( n15795 , n15793 , n15794 );
buf ( n15796 , n5685 );
buf ( n15797 , n15796 );
not ( n15798 , n15797 );
buf ( n15799 , n5686 );
not ( n15800 , n15799 );
not ( n15801 , n15800 );
or ( n15802 , n15798 , n15801 );
not ( n15803 , n15796 );
buf ( n15804 , n15799 );
nand ( n15805 , n15803 , n15804 );
nand ( n15806 , n15802 , n15805 );
buf ( n15807 , n5687 );
buf ( n15808 , n15807 );
and ( n15809 , n15806 , n15808 );
not ( n15810 , n15806 );
not ( n15811 , n15807 );
and ( n15812 , n15810 , n15811 );
nor ( n15813 , n15809 , n15812 );
buf ( n15814 , n5688 );
nand ( n15815 , n6927 , n15814 );
buf ( n15816 , n5689 );
buf ( n15817 , n15816 );
and ( n15818 , n15815 , n15817 );
not ( n15819 , n15815 );
not ( n15820 , n15816 );
and ( n15821 , n15819 , n15820 );
nor ( n15822 , n15818 , n15821 );
xor ( n15823 , n15813 , n15822 );
buf ( n15824 , n5690 );
nand ( n15825 , n14573 , n15824 );
buf ( n15826 , n5691 );
not ( n15827 , n15826 );
and ( n15828 , n15825 , n15827 );
not ( n15829 , n15825 );
buf ( n15830 , n15826 );
and ( n15831 , n15829 , n15830 );
nor ( n15832 , n15828 , n15831 );
xor ( n15833 , n15823 , n15832 );
not ( n15834 , n15833 );
not ( n15835 , n15834 );
and ( n15836 , n15795 , n15835 );
not ( n15837 , n15795 );
xor ( n15838 , n15813 , n15822 );
xnor ( n15839 , n15838 , n15832 );
buf ( n15840 , n15839 );
and ( n15841 , n15837 , n15840 );
nor ( n15842 , n15836 , n15841 );
not ( n15843 , n15842 );
not ( n15844 , n8547 );
not ( n15845 , n6589 );
and ( n15846 , n15844 , n15845 );
and ( n15847 , n8547 , n6589 );
nor ( n15848 , n15846 , n15847 );
not ( n15849 , n10443 );
and ( n15850 , n15848 , n15849 );
not ( n15851 , n15848 );
and ( n15852 , n15851 , n10443 );
nor ( n15853 , n15850 , n15852 );
not ( n15854 , n15853 );
nand ( n15855 , n15843 , n15854 );
buf ( n15856 , n5692 );
not ( n15857 , n7499 );
buf ( n15858 , n5693 );
not ( n15859 , n15858 );
not ( n15860 , n15859 );
or ( n15861 , n15857 , n15860 );
not ( n15862 , n7498 );
buf ( n15863 , n15858 );
nand ( n15864 , n15862 , n15863 );
nand ( n15865 , n15861 , n15864 );
xor ( n15866 , n15856 , n15865 );
buf ( n15867 , n5694 );
buf ( n15868 , n5695 );
buf ( n15869 , n15868 );
xor ( n15870 , n15867 , n15869 );
buf ( n15871 , n5696 );
nand ( n15872 , n6973 , n15871 );
xnor ( n15873 , n15870 , n15872 );
xnor ( n15874 , n15866 , n15873 );
not ( n15875 , n15874 );
buf ( n15876 , n5697 );
buf ( n15877 , n15876 );
not ( n15878 , n15877 );
not ( n15879 , n10025 );
buf ( n15880 , n5698 );
not ( n15881 , n15880 );
not ( n15882 , n15881 );
or ( n15883 , n15879 , n15882 );
not ( n15884 , n10024 );
buf ( n15885 , n15880 );
nand ( n15886 , n15884 , n15885 );
nand ( n15887 , n15883 , n15886 );
buf ( n15888 , n5699 );
buf ( n15889 , n15888 );
and ( n15890 , n15887 , n15889 );
not ( n15891 , n15887 );
not ( n15892 , n15888 );
and ( n15893 , n15891 , n15892 );
nor ( n15894 , n15890 , n15893 );
xor ( n15895 , n15894 , n8933 );
buf ( n15896 , n5700 );
nand ( n15897 , n6515 , n15896 );
buf ( n15898 , n5701 );
not ( n15899 , n15898 );
and ( n15900 , n15897 , n15899 );
not ( n15901 , n15897 );
buf ( n15902 , n15898 );
and ( n15903 , n15901 , n15902 );
nor ( n15904 , n15900 , n15903 );
xnor ( n15905 , n15895 , n15904 );
not ( n15906 , n15905 );
not ( n15907 , n15906 );
or ( n15908 , n15878 , n15907 );
or ( n15909 , n15906 , n15877 );
nand ( n15910 , n15908 , n15909 );
and ( n15911 , n15875 , n15910 );
not ( n15912 , n15875 );
not ( n15913 , n15910 );
and ( n15914 , n15912 , n15913 );
nor ( n15915 , n15911 , n15914 );
not ( n15916 , n15915 );
and ( n15917 , n15855 , n15916 );
not ( n15918 , n15855 );
and ( n15919 , n15918 , n15915 );
nor ( n15920 , n15917 , n15919 );
not ( n15921 , n15920 );
or ( n15922 , n15759 , n15921 );
or ( n15923 , n15920 , n15758 );
nand ( n15924 , n15922 , n15923 );
nand ( n15925 , n15579 , n15477 );
not ( n15926 , n15925 );
buf ( n15927 , n5702 );
buf ( n15928 , n15927 );
buf ( n15929 , n5703 );
nand ( n15930 , n6557 , n15929 );
buf ( n15931 , n5704 );
buf ( n15932 , n15931 );
and ( n15933 , n15930 , n15932 );
not ( n15934 , n15930 );
not ( n15935 , n15931 );
and ( n15936 , n15934 , n15935 );
nor ( n15937 , n15933 , n15936 );
not ( n15938 , n15937 );
buf ( n15939 , n5705 );
nand ( n15940 , n7197 , n15939 );
buf ( n15941 , n5706 );
not ( n15942 , n15941 );
and ( n15943 , n15940 , n15942 );
not ( n15944 , n15940 );
buf ( n15945 , n15941 );
and ( n15946 , n15944 , n15945 );
nor ( n15947 , n15943 , n15946 );
not ( n15948 , n15947 );
or ( n15949 , n15938 , n15948 );
or ( n15950 , n15937 , n15947 );
nand ( n15951 , n15949 , n15950 );
buf ( n15952 , n5707 );
buf ( n15953 , n15952 );
not ( n15954 , n15953 );
buf ( n15955 , n5708 );
not ( n15956 , n15955 );
not ( n15957 , n15956 );
or ( n15958 , n15954 , n15957 );
not ( n15959 , n15952 );
buf ( n15960 , n15955 );
nand ( n15961 , n15959 , n15960 );
nand ( n15962 , n15958 , n15961 );
buf ( n15963 , n5709 );
not ( n15964 , n15963 );
and ( n15965 , n15962 , n15964 );
not ( n15966 , n15962 );
buf ( n15967 , n15963 );
and ( n15968 , n15966 , n15967 );
nor ( n15969 , n15965 , n15968 );
and ( n15970 , n15951 , n15969 );
not ( n15971 , n15951 );
not ( n15972 , n15969 );
and ( n15973 , n15971 , n15972 );
nor ( n15974 , n15970 , n15973 );
not ( n15975 , n15974 );
not ( n15976 , n15975 );
xor ( n15977 , n15928 , n15976 );
buf ( n15978 , n5710 );
buf ( n15979 , n15978 );
not ( n15980 , n15979 );
buf ( n15981 , n5711 );
not ( n15982 , n15981 );
not ( n15983 , n15982 );
or ( n15984 , n15980 , n15983 );
not ( n15985 , n15978 );
buf ( n15986 , n15981 );
nand ( n15987 , n15985 , n15986 );
nand ( n15988 , n15984 , n15987 );
not ( n15989 , n15988 );
not ( n15990 , n15989 );
buf ( n15991 , n5712 );
buf ( n15992 , n5713 );
not ( n15993 , n15992 );
xor ( n15994 , n15991 , n15993 );
buf ( n15995 , n5714 );
not ( n15996 , n15995 );
buf ( n15997 , n5715 );
nand ( n15998 , n6646 , n15997 );
not ( n15999 , n15998 );
or ( n16000 , n15996 , n15999 );
nand ( n16001 , n6604 , n15997 );
or ( n16002 , n16001 , n15995 );
nand ( n16003 , n16000 , n16002 );
xnor ( n16004 , n15994 , n16003 );
not ( n16005 , n16004 );
or ( n16006 , n15990 , n16005 );
or ( n16007 , n16004 , n15989 );
nand ( n16008 , n16006 , n16007 );
buf ( n16009 , n16008 );
not ( n16010 , n16009 );
xnor ( n16011 , n15977 , n16010 );
not ( n16012 , n16011 );
not ( n16013 , n16012 );
and ( n16014 , n15926 , n16013 );
and ( n16015 , n15925 , n16012 );
nor ( n16016 , n16014 , n16015 );
and ( n16017 , n15924 , n16016 );
not ( n16018 , n15924 );
not ( n16019 , n16016 );
and ( n16020 , n16018 , n16019 );
nor ( n16021 , n16017 , n16020 );
not ( n16022 , n16021 );
not ( n16023 , n16022 );
not ( n16024 , n16023 );
buf ( n16025 , n15822 );
not ( n16026 , n16025 );
not ( n16027 , n16026 );
buf ( n16028 , n5716 );
buf ( n16029 , n16028 );
not ( n16030 , n16029 );
buf ( n16031 , n5717 );
not ( n16032 , n16031 );
not ( n16033 , n16032 );
or ( n16034 , n16030 , n16033 );
not ( n16035 , n16028 );
buf ( n16036 , n16031 );
nand ( n16037 , n16035 , n16036 );
nand ( n16038 , n16034 , n16037 );
buf ( n16039 , n5718 );
not ( n16040 , n16039 );
and ( n16041 , n16038 , n16040 );
not ( n16042 , n16038 );
buf ( n16043 , n16039 );
and ( n16044 , n16042 , n16043 );
nor ( n16045 , n16041 , n16044 );
xor ( n16046 , n16045 , n14111 );
buf ( n16047 , n5719 );
nand ( n16048 , n6647 , n16047 );
buf ( n16049 , n5720 );
buf ( n16050 , n16049 );
and ( n16051 , n16048 , n16050 );
not ( n16052 , n16048 );
not ( n16053 , n16049 );
and ( n16054 , n16052 , n16053 );
nor ( n16055 , n16051 , n16054 );
xnor ( n16056 , n16046 , n16055 );
buf ( n16057 , n16056 );
not ( n16058 , n16057 );
not ( n16059 , n16058 );
or ( n16060 , n16027 , n16059 );
buf ( n16061 , n16057 );
nand ( n16062 , n16061 , n16025 );
nand ( n16063 , n16060 , n16062 );
buf ( n16064 , n5721 );
buf ( n16065 , n5722 );
not ( n16066 , n16065 );
buf ( n16067 , n5723 );
buf ( n16068 , n16067 );
nand ( n16069 , n16066 , n16068 );
not ( n16070 , n16067 );
buf ( n16071 , n16065 );
nand ( n16072 , n16070 , n16071 );
and ( n16073 , n16069 , n16072 );
xor ( n16074 , n16064 , n16073 );
buf ( n16075 , n5724 );
nand ( n16076 , n6633 , n16075 );
buf ( n16077 , n5725 );
buf ( n16078 , n16077 );
and ( n16079 , n16076 , n16078 );
not ( n16080 , n16076 );
not ( n16081 , n16077 );
and ( n16082 , n16080 , n16081 );
nor ( n16083 , n16079 , n16082 );
not ( n16084 , n16083 );
buf ( n16085 , n5726 );
nand ( n16086 , n6815 , n16085 );
buf ( n16087 , n5727 );
not ( n16088 , n16087 );
and ( n16089 , n16086 , n16088 );
not ( n16090 , n16086 );
buf ( n16091 , n16087 );
and ( n16092 , n16090 , n16091 );
nor ( n16093 , n16089 , n16092 );
not ( n16094 , n16093 );
or ( n16095 , n16084 , n16094 );
or ( n16096 , n16083 , n16093 );
nand ( n16097 , n16095 , n16096 );
xnor ( n16098 , n16074 , n16097 );
buf ( n16099 , n16098 );
not ( n16100 , n16099 );
and ( n16101 , n16063 , n16100 );
not ( n16102 , n16063 );
not ( n16103 , n16098 );
not ( n16104 , n16103 );
and ( n16105 , n16102 , n16104 );
nor ( n16106 , n16101 , n16105 );
not ( n16107 , n16106 );
buf ( n16108 , n5728 );
buf ( n16109 , n16108 );
buf ( n16110 , n5729 );
buf ( n16111 , n16110 );
not ( n16112 , n16111 );
buf ( n16113 , n5730 );
not ( n16114 , n16113 );
not ( n16115 , n16114 );
or ( n16116 , n16112 , n16115 );
not ( n16117 , n16110 );
buf ( n16118 , n16113 );
nand ( n16119 , n16117 , n16118 );
nand ( n16120 , n16116 , n16119 );
buf ( n16121 , n5731 );
not ( n16122 , n16121 );
and ( n16123 , n16120 , n16122 );
not ( n16124 , n16120 );
buf ( n16125 , n16121 );
and ( n16126 , n16124 , n16125 );
nor ( n16127 , n16123 , n16126 );
buf ( n16128 , n5732 );
nand ( n16129 , n8537 , n16128 );
buf ( n16130 , n5733 );
buf ( n16131 , n16130 );
and ( n16132 , n16129 , n16131 );
not ( n16133 , n16129 );
not ( n16134 , n16130 );
and ( n16135 , n16133 , n16134 );
nor ( n16136 , n16132 , n16135 );
xor ( n16137 , n16127 , n16136 );
buf ( n16138 , n5734 );
nand ( n16139 , n7014 , n16138 );
buf ( n16140 , n5735 );
not ( n16141 , n16140 );
and ( n16142 , n16139 , n16141 );
not ( n16143 , n16139 );
buf ( n16144 , n16140 );
and ( n16145 , n16143 , n16144 );
nor ( n16146 , n16142 , n16145 );
xnor ( n16147 , n16137 , n16146 );
not ( n16148 , n16147 );
not ( n16149 , n16148 );
xor ( n16150 , n16109 , n16149 );
not ( n16151 , n11775 );
xnor ( n16152 , n16150 , n16151 );
nand ( n16153 , n16107 , n16152 );
not ( n16154 , n16153 );
buf ( n16155 , n8896 );
xor ( n16156 , n16155 , n13690 );
buf ( n16157 , n5736 );
buf ( n16158 , n16157 );
not ( n16159 , n16158 );
buf ( n16160 , n5737 );
not ( n16161 , n16160 );
not ( n16162 , n16161 );
or ( n16163 , n16159 , n16162 );
not ( n16164 , n16157 );
buf ( n16165 , n16160 );
nand ( n16166 , n16164 , n16165 );
nand ( n16167 , n16163 , n16166 );
not ( n16168 , n16167 );
buf ( n16169 , n5738 );
buf ( n16170 , n5739 );
nand ( n16171 , n8454 , n16170 );
buf ( n16172 , n5740 );
buf ( n16173 , n16172 );
and ( n16174 , n16171 , n16173 );
not ( n16175 , n16171 );
not ( n16176 , n16172 );
and ( n16177 , n16175 , n16176 );
nor ( n16178 , n16174 , n16177 );
xor ( n16179 , n16169 , n16178 );
buf ( n16180 , n5741 );
nand ( n16181 , n6647 , n16180 );
buf ( n16182 , n5742 );
not ( n16183 , n16182 );
and ( n16184 , n16181 , n16183 );
not ( n16185 , n16181 );
buf ( n16186 , n16182 );
and ( n16187 , n16185 , n16186 );
nor ( n16188 , n16184 , n16187 );
xnor ( n16189 , n16179 , n16188 );
not ( n16190 , n16189 );
not ( n16191 , n16190 );
or ( n16192 , n16168 , n16191 );
not ( n16193 , n16167 );
nand ( n16194 , n16189 , n16193 );
nand ( n16195 , n16192 , n16194 );
buf ( n16196 , n16195 );
not ( n16197 , n16196 );
xnor ( n16198 , n16156 , n16197 );
not ( n16199 , n16198 );
not ( n16200 , n16199 );
and ( n16201 , n16154 , n16200 );
and ( n16202 , n16153 , n16199 );
nor ( n16203 , n16201 , n16202 );
not ( n16204 , n16203 );
not ( n16205 , n12410 );
not ( n16206 , n6659 );
or ( n16207 , n16205 , n16206 );
or ( n16208 , n6659 , n12410 );
nand ( n16209 , n16207 , n16208 );
and ( n16210 , n16209 , n12287 );
not ( n16211 , n16209 );
not ( n16212 , n12287 );
and ( n16213 , n16211 , n16212 );
nor ( n16214 , n16210 , n16213 );
not ( n16215 , n16214 );
not ( n16216 , n16215 );
buf ( n16217 , n5743 );
not ( n16218 , n16217 );
not ( n16219 , n12128 );
or ( n16220 , n16218 , n16219 );
or ( n16221 , n12128 , n16217 );
nand ( n16222 , n16220 , n16221 );
not ( n16223 , n13023 );
not ( n16224 , n13043 );
or ( n16225 , n16223 , n16224 );
not ( n16226 , n13023 );
nand ( n16227 , n13042 , n16226 );
nand ( n16228 , n16225 , n16227 );
buf ( n16229 , n16228 );
buf ( n16230 , n16229 );
and ( n16231 , n16222 , n16230 );
not ( n16232 , n16222 );
not ( n16233 , n16229 );
and ( n16234 , n16232 , n16233 );
nor ( n16235 , n16231 , n16234 );
not ( n16236 , n16235 );
buf ( n16237 , n5744 );
nand ( n16238 , n10947 , n16237 );
buf ( n16239 , n16238 );
buf ( n16240 , n5745 );
buf ( n16241 , n16240 );
and ( n16242 , n16239 , n16241 );
not ( n16243 , n16239 );
not ( n16244 , n16240 );
and ( n16245 , n16243 , n16244 );
nor ( n16246 , n16242 , n16245 );
not ( n16247 , n16246 );
not ( n16248 , n16247 );
xor ( n16249 , n10994 , n11013 );
xnor ( n16250 , n16249 , n11003 );
buf ( n16251 , n16250 );
not ( n16252 , n16251 );
or ( n16253 , n16248 , n16252 );
buf ( n16254 , n11015 );
nand ( n16255 , n16254 , n16246 );
nand ( n16256 , n16253 , n16255 );
buf ( n16257 , n11054 );
not ( n16258 , n16257 );
buf ( n16259 , n16258 );
and ( n16260 , n16256 , n16259 );
not ( n16261 , n16256 );
not ( n16262 , n16259 );
and ( n16263 , n16261 , n16262 );
nor ( n16264 , n16260 , n16263 );
nand ( n16265 , n16236 , n16264 );
not ( n16266 , n16265 );
or ( n16267 , n16216 , n16266 );
or ( n16268 , n16265 , n16215 );
nand ( n16269 , n16267 , n16268 );
not ( n16270 , n16269 );
and ( n16271 , n16204 , n16270 );
and ( n16272 , n16203 , n16269 );
nor ( n16273 , n16271 , n16272 );
not ( n16274 , n16273 );
not ( n16275 , n16274 );
and ( n16276 , n16024 , n16275 );
and ( n16277 , n16023 , n16274 );
nor ( n16278 , n16276 , n16277 );
not ( n16279 , n16278 );
or ( n16280 , n15584 , n16279 );
not ( n16281 , n15583 );
not ( n16282 , n16273 );
not ( n16283 , n16282 );
not ( n16284 , n16021 );
or ( n16285 , n16283 , n16284 );
nand ( n16286 , n16022 , n16273 );
nand ( n16287 , n16285 , n16286 );
nand ( n16288 , n16281 , n16287 );
nand ( n16289 , n16280 , n16288 );
buf ( n16290 , n5746 );
nand ( n16291 , n7107 , n16290 );
buf ( n16292 , n5747 );
buf ( n16293 , n16292 );
and ( n16294 , n16291 , n16293 );
not ( n16295 , n16291 );
not ( n16296 , n16292 );
and ( n16297 , n16295 , n16296 );
nor ( n16298 , n16294 , n16297 );
not ( n16299 , n16298 );
not ( n16300 , n16299 );
buf ( n16301 , n5748 );
buf ( n16302 , n16301 );
not ( n16303 , n16302 );
buf ( n16304 , n5749 );
not ( n16305 , n16304 );
not ( n16306 , n16305 );
or ( n16307 , n16303 , n16306 );
not ( n16308 , n16301 );
buf ( n16309 , n16304 );
nand ( n16310 , n16308 , n16309 );
nand ( n16311 , n16307 , n16310 );
buf ( n16312 , n5750 );
not ( n16313 , n16312 );
and ( n16314 , n16311 , n16313 );
not ( n16315 , n16311 );
buf ( n16316 , n16312 );
and ( n16317 , n16315 , n16316 );
nor ( n16318 , n16314 , n16317 );
buf ( n16319 , n5751 );
nand ( n16320 , n7013 , n16319 );
buf ( n16321 , n5752 );
buf ( n16322 , n16321 );
and ( n16323 , n16320 , n16322 );
not ( n16324 , n16320 );
not ( n16325 , n16321 );
and ( n16326 , n16324 , n16325 );
nor ( n16327 , n16323 , n16326 );
xor ( n16328 , n16318 , n16327 );
buf ( n16329 , n5753 );
nand ( n16330 , n8176 , n16329 );
buf ( n16331 , n5754 );
not ( n16332 , n16331 );
and ( n16333 , n16330 , n16332 );
not ( n16334 , n16330 );
buf ( n16335 , n16331 );
and ( n16336 , n16334 , n16335 );
nor ( n16337 , n16333 , n16336 );
xnor ( n16338 , n16328 , n16337 );
not ( n16339 , n16338 );
xor ( n16340 , n16300 , n16339 );
buf ( n16341 , n5755 );
buf ( n16342 , n16341 );
not ( n16343 , n13401 );
buf ( n16344 , n5756 );
buf ( n16345 , n16344 );
and ( n16346 , n16343 , n16345 );
not ( n16347 , n16343 );
not ( n16348 , n16344 );
and ( n16349 , n16347 , n16348 );
nor ( n16350 , n16346 , n16349 );
xor ( n16351 , n16342 , n16350 );
buf ( n16352 , n5757 );
buf ( n16353 , n5758 );
xor ( n16354 , n16352 , n16353 );
buf ( n16355 , n5759 );
nand ( n16356 , n8223 , n16355 );
xnor ( n16357 , n16354 , n16356 );
xnor ( n16358 , n16351 , n16357 );
buf ( n16359 , n16358 );
xnor ( n16360 , n16340 , n16359 );
not ( n16361 , n16360 );
not ( n16362 , n6906 );
not ( n16363 , n13133 );
or ( n16364 , n16362 , n16363 );
or ( n16365 , n13133 , n6906 );
nand ( n16366 , n16364 , n16365 );
not ( n16367 , n16366 );
not ( n16368 , n14458 );
and ( n16369 , n16367 , n16368 );
and ( n16370 , n16366 , n14458 );
nor ( n16371 , n16369 , n16370 );
not ( n16372 , n16371 );
nand ( n16373 , n16361 , n16372 );
not ( n16374 , n16373 );
buf ( n16375 , n9725 );
not ( n16376 , n16375 );
not ( n16377 , n6526 );
or ( n16378 , n16376 , n16377 );
or ( n16379 , n6526 , n16375 );
nand ( n16380 , n16378 , n16379 );
not ( n16381 , n6572 );
and ( n16382 , n16380 , n16381 );
not ( n16383 , n16380 );
and ( n16384 , n16383 , n6572 );
nor ( n16385 , n16382 , n16384 );
not ( n16386 , n16385 );
and ( n16387 , n16374 , n16386 );
and ( n16388 , n16373 , n16385 );
nor ( n16389 , n16387 , n16388 );
not ( n16390 , n16389 );
not ( n16391 , n16390 );
not ( n16392 , n16229 );
buf ( n16393 , n5760 );
nand ( n16394 , n8781 , n16393 );
buf ( n16395 , n5761 );
buf ( n16396 , n16395 );
and ( n16397 , n16394 , n16396 );
not ( n16398 , n16394 );
not ( n16399 , n16395 );
and ( n16400 , n16398 , n16399 );
nor ( n16401 , n16397 , n16400 );
buf ( n16402 , n16401 );
not ( n16403 , n12127 );
and ( n16404 , n16402 , n16403 );
not ( n16405 , n16402 );
xor ( n16406 , n12107 , n12116 );
not ( n16407 , n12126 );
xnor ( n16408 , n16406 , n16407 );
and ( n16409 , n16405 , n16408 );
nor ( n16410 , n16404 , n16409 );
not ( n16411 , n16410 );
and ( n16412 , n16392 , n16411 );
and ( n16413 , n16229 , n16410 );
nor ( n16414 , n16412 , n16413 );
buf ( n16415 , n5762 );
buf ( n16416 , n16415 );
not ( n16417 , n16416 );
buf ( n16418 , n5763 );
not ( n16419 , n16418 );
not ( n16420 , n16419 );
or ( n16421 , n16417 , n16420 );
not ( n16422 , n16415 );
buf ( n16423 , n16418 );
nand ( n16424 , n16422 , n16423 );
nand ( n16425 , n16421 , n16424 );
buf ( n16426 , n5764 );
buf ( n16427 , n16426 );
and ( n16428 , n16425 , n16427 );
not ( n16429 , n16425 );
not ( n16430 , n16426 );
and ( n16431 , n16429 , n16430 );
nor ( n16432 , n16428 , n16431 );
buf ( n16433 , n5765 );
nand ( n16434 , n9160 , n16433 );
buf ( n16435 , n5766 );
not ( n16436 , n16435 );
and ( n16437 , n16434 , n16436 );
not ( n16438 , n16434 );
buf ( n16439 , n16435 );
and ( n16440 , n16438 , n16439 );
nor ( n16441 , n16437 , n16440 );
xor ( n16442 , n16432 , n16441 );
buf ( n16443 , n5767 );
nand ( n16444 , n6647 , n16443 );
buf ( n16445 , n5768 );
not ( n16446 , n16445 );
and ( n16447 , n16444 , n16446 );
not ( n16448 , n16444 );
buf ( n16449 , n16445 );
and ( n16450 , n16448 , n16449 );
nor ( n16451 , n16447 , n16450 );
xnor ( n16452 , n16442 , n16451 );
not ( n16453 , n16452 );
not ( n16454 , n16453 );
not ( n16455 , n16454 );
not ( n16456 , n7643 );
and ( n16457 , n16455 , n16456 );
buf ( n16458 , n16452 );
and ( n16459 , n16458 , n7643 );
nor ( n16460 , n16457 , n16459 );
not ( n16461 , n15928 );
buf ( n16462 , n5769 );
not ( n16463 , n16462 );
not ( n16464 , n16463 );
or ( n16465 , n16461 , n16464 );
not ( n16466 , n15927 );
buf ( n16467 , n16462 );
nand ( n16468 , n16466 , n16467 );
nand ( n16469 , n16465 , n16468 );
buf ( n16470 , n5770 );
not ( n16471 , n16470 );
and ( n16472 , n16469 , n16471 );
not ( n16473 , n16469 );
buf ( n16474 , n16470 );
and ( n16475 , n16473 , n16474 );
nor ( n16476 , n16472 , n16475 );
buf ( n16477 , n5771 );
nand ( n16478 , n7698 , n16477 );
buf ( n16479 , n5772 );
xor ( n16480 , n16478 , n16479 );
xor ( n16481 , n16476 , n16480 );
buf ( n16482 , n5773 );
nand ( n16483 , n13581 , n16482 );
buf ( n16484 , n5774 );
not ( n16485 , n16484 );
and ( n16486 , n16483 , n16485 );
not ( n16487 , n16483 );
buf ( n16488 , n16484 );
and ( n16489 , n16487 , n16488 );
nor ( n16490 , n16486 , n16489 );
xnor ( n16491 , n16481 , n16490 );
not ( n16492 , n16491 );
not ( n16493 , n16492 );
and ( n16494 , n16460 , n16493 );
not ( n16495 , n16460 );
buf ( n16496 , n16491 );
not ( n16497 , n16496 );
and ( n16498 , n16495 , n16497 );
nor ( n16499 , n16494 , n16498 );
nand ( n16500 , n16414 , n16499 );
not ( n16501 , n16500 );
buf ( n16502 , n5775 );
buf ( n16503 , n16502 );
not ( n16504 , n16503 );
buf ( n16505 , n5776 );
not ( n16506 , n16505 );
not ( n16507 , n16506 );
or ( n16508 , n16504 , n16507 );
not ( n16509 , n16502 );
buf ( n16510 , n16505 );
nand ( n16511 , n16509 , n16510 );
nand ( n16512 , n16508 , n16511 );
buf ( n16513 , n5777 );
not ( n16514 , n16513 );
and ( n16515 , n16512 , n16514 );
not ( n16516 , n16512 );
buf ( n16517 , n16513 );
and ( n16518 , n16516 , n16517 );
nor ( n16519 , n16515 , n16518 );
buf ( n16520 , n5778 );
nand ( n16521 , n8537 , n16520 );
buf ( n16522 , n5779 );
buf ( n16523 , n16522 );
and ( n16524 , n16521 , n16523 );
not ( n16525 , n16521 );
not ( n16526 , n16522 );
and ( n16527 , n16525 , n16526 );
nor ( n16528 , n16524 , n16527 );
xor ( n16529 , n16519 , n16528 );
buf ( n16530 , n5780 );
nand ( n16531 , n7107 , n16530 );
buf ( n16532 , n5781 );
buf ( n16533 , n16532 );
and ( n16534 , n16531 , n16533 );
not ( n16535 , n16531 );
not ( n16536 , n16532 );
and ( n16537 , n16535 , n16536 );
nor ( n16538 , n16534 , n16537 );
not ( n16539 , n16538 );
xor ( n16540 , n16529 , n16539 );
not ( n16541 , n16540 );
not ( n16542 , n16541 );
buf ( n16543 , n5782 );
nand ( n16544 , n8364 , n16543 );
buf ( n16545 , n5783 );
buf ( n16546 , n16545 );
and ( n16547 , n16544 , n16546 );
not ( n16548 , n16544 );
not ( n16549 , n16545 );
and ( n16550 , n16548 , n16549 );
nor ( n16551 , n16547 , n16550 );
buf ( n16552 , n16551 );
not ( n16553 , n16552 );
not ( n16554 , n16553 );
buf ( n16555 , n5784 );
buf ( n16556 , n16555 );
not ( n16557 , n16556 );
buf ( n16558 , n5785 );
not ( n16559 , n16558 );
not ( n16560 , n16559 );
or ( n16561 , n16557 , n16560 );
not ( n16562 , n16555 );
buf ( n16563 , n16558 );
nand ( n16564 , n16562 , n16563 );
nand ( n16565 , n16561 , n16564 );
buf ( n16566 , n5786 );
not ( n16567 , n16566 );
and ( n16568 , n16565 , n16567 );
not ( n16569 , n16565 );
buf ( n16570 , n16566 );
and ( n16571 , n16569 , n16570 );
nor ( n16572 , n16568 , n16571 );
buf ( n16573 , n5787 );
nand ( n16574 , n9160 , n16573 );
buf ( n16575 , n5788 );
not ( n16576 , n16575 );
and ( n16577 , n16574 , n16576 );
not ( n16578 , n16574 );
buf ( n16579 , n16575 );
and ( n16580 , n16578 , n16579 );
nor ( n16581 , n16577 , n16580 );
xor ( n16582 , n16572 , n16581 );
buf ( n16583 , n5789 );
nand ( n16584 , n7258 , n16583 );
buf ( n16585 , n5790 );
not ( n16586 , n16585 );
and ( n16587 , n16584 , n16586 );
not ( n16588 , n16584 );
buf ( n16589 , n16585 );
and ( n16590 , n16588 , n16589 );
nor ( n16591 , n16587 , n16590 );
xnor ( n16592 , n16582 , n16591 );
not ( n16593 , n16592 );
not ( n16594 , n16593 );
or ( n16595 , n16554 , n16594 );
not ( n16596 , n16592 );
not ( n16597 , n16596 );
nand ( n16598 , n16597 , n16552 );
nand ( n16599 , n16595 , n16598 );
not ( n16600 , n16599 );
or ( n16601 , n16542 , n16600 );
or ( n16602 , n16599 , n16541 );
nand ( n16603 , n16601 , n16602 );
not ( n16604 , n16603 );
and ( n16605 , n16501 , n16604 );
and ( n16606 , n16500 , n16603 );
nor ( n16607 , n16605 , n16606 );
not ( n16608 , n16607 );
not ( n16609 , n16195 );
not ( n16610 , n16609 );
and ( n16611 , n9642 , n8885 );
not ( n16612 , n9642 );
and ( n16613 , n16612 , n8886 );
or ( n16614 , n16611 , n16613 );
not ( n16615 , n16614 );
and ( n16616 , n16610 , n16615 );
and ( n16617 , n16609 , n16614 );
nor ( n16618 , n16616 , n16617 );
not ( n16619 , n9290 );
buf ( n16620 , n5791 );
buf ( n16621 , n16620 );
not ( n16622 , n16621 );
buf ( n16623 , n5792 );
not ( n16624 , n16623 );
not ( n16625 , n16624 );
or ( n16626 , n16622 , n16625 );
not ( n16627 , n16620 );
buf ( n16628 , n16623 );
nand ( n16629 , n16627 , n16628 );
nand ( n16630 , n16626 , n16629 );
buf ( n16631 , n5793 );
buf ( n16632 , n16631 );
and ( n16633 , n16630 , n16632 );
not ( n16634 , n16630 );
not ( n16635 , n16631 );
and ( n16636 , n16634 , n16635 );
nor ( n16637 , n16633 , n16636 );
buf ( n16638 , n5794 );
nand ( n16639 , n7868 , n16638 );
buf ( n16640 , n5795 );
buf ( n16641 , n16640 );
and ( n16642 , n16639 , n16641 );
not ( n16643 , n16639 );
not ( n16644 , n16640 );
and ( n16645 , n16643 , n16644 );
nor ( n16646 , n16642 , n16645 );
xor ( n16647 , n16637 , n16646 );
buf ( n16648 , n5796 );
nand ( n16649 , n7912 , n16648 );
buf ( n16650 , n5797 );
buf ( n16651 , n16650 );
and ( n16652 , n16649 , n16651 );
not ( n16653 , n16649 );
not ( n16654 , n16650 );
and ( n16655 , n16653 , n16654 );
nor ( n16656 , n16652 , n16655 );
xnor ( n16657 , n16647 , n16656 );
buf ( n16658 , n16657 );
not ( n16659 , n16658 );
or ( n16660 , n16619 , n16659 );
not ( n16661 , n16657 );
not ( n16662 , n16661 );
or ( n16663 , n16662 , n9290 );
nand ( n16664 , n16660 , n16663 );
buf ( n16665 , n5798 );
buf ( n16666 , n16665 );
buf ( n16667 , n5799 );
buf ( n16668 , n16667 );
not ( n16669 , n16668 );
buf ( n16670 , n5800 );
not ( n16671 , n16670 );
not ( n16672 , n16671 );
or ( n16673 , n16669 , n16672 );
not ( n16674 , n16667 );
buf ( n16675 , n16670 );
nand ( n16676 , n16674 , n16675 );
nand ( n16677 , n16673 , n16676 );
xor ( n16678 , n16666 , n16677 );
xor ( n16679 , n10978 , n16244 );
xnor ( n16680 , n16679 , n16238 );
xnor ( n16681 , n16678 , n16680 );
not ( n16682 , n16681 );
and ( n16683 , n16664 , n16682 );
not ( n16684 , n16664 );
not ( n16685 , n16682 );
and ( n16686 , n16684 , n16685 );
or ( n16687 , n16683 , n16686 );
nand ( n16688 , n16618 , n16687 );
not ( n16689 , n14150 );
not ( n16690 , n15518 );
or ( n16691 , n16689 , n16690 );
not ( n16692 , n14150 );
nand ( n16693 , n16692 , n15521 );
nand ( n16694 , n16691 , n16693 );
and ( n16695 , n16694 , n15563 );
not ( n16696 , n16694 );
and ( n16697 , n16696 , n15576 );
nor ( n16698 , n16695 , n16697 );
not ( n16699 , n16698 );
and ( n16700 , n16688 , n16699 );
not ( n16701 , n16688 );
and ( n16702 , n16701 , n16698 );
nor ( n16703 , n16700 , n16702 );
not ( n16704 , n16703 );
or ( n16705 , n16608 , n16704 );
or ( n16706 , n16703 , n16607 );
nand ( n16707 , n16705 , n16706 );
not ( n16708 , n16707 );
not ( n16709 , n16708 );
or ( n16710 , n16391 , n16709 );
nand ( n16711 , n16707 , n16389 );
nand ( n16712 , n16710 , n16711 );
buf ( n16713 , n14555 );
xor ( n16714 , n16713 , n14567 );
xnor ( n16715 , n16714 , n14576 );
buf ( n16716 , n16715 );
not ( n16717 , n16716 );
buf ( n16718 , n8373 );
not ( n16719 , n16718 );
not ( n16720 , n7679 );
buf ( n16721 , n5801 );
not ( n16722 , n16721 );
not ( n16723 , n16722 );
or ( n16724 , n16720 , n16723 );
not ( n16725 , n7678 );
buf ( n16726 , n16721 );
nand ( n16727 , n16725 , n16726 );
nand ( n16728 , n16724 , n16727 );
buf ( n16729 , n5802 );
buf ( n16730 , n16729 );
and ( n16731 , n16728 , n16730 );
not ( n16732 , n16728 );
not ( n16733 , n16729 );
and ( n16734 , n16732 , n16733 );
nor ( n16735 , n16731 , n16734 );
buf ( n16736 , n5803 );
nand ( n16737 , n8364 , n16736 );
buf ( n16738 , n5804 );
buf ( n16739 , n16738 );
and ( n16740 , n16737 , n16739 );
not ( n16741 , n16737 );
not ( n16742 , n16738 );
and ( n16743 , n16741 , n16742 );
nor ( n16744 , n16740 , n16743 );
xor ( n16745 , n16735 , n16744 );
buf ( n16746 , n5805 );
nand ( n16747 , n8608 , n16746 );
buf ( n16748 , n5806 );
buf ( n16749 , n16748 );
and ( n16750 , n16747 , n16749 );
not ( n16751 , n16747 );
not ( n16752 , n16748 );
and ( n16753 , n16751 , n16752 );
nor ( n16754 , n16750 , n16753 );
xnor ( n16755 , n16745 , n16754 );
not ( n16756 , n16755 );
not ( n16757 , n16756 );
or ( n16758 , n16719 , n16757 );
or ( n16759 , n16756 , n16718 );
nand ( n16760 , n16758 , n16759 );
not ( n16761 , n16760 );
and ( n16762 , n16717 , n16761 );
not ( n16763 , n16715 );
not ( n16764 , n16763 );
and ( n16765 , n16764 , n16760 );
nor ( n16766 , n16762 , n16765 );
not ( n16767 , n16766 );
not ( n16768 , n16767 );
not ( n16769 , n11710 );
buf ( n16770 , n5807 );
not ( n16771 , n16770 );
buf ( n16772 , n5808 );
not ( n16773 , n16772 );
nand ( n16774 , n16773 , n13862 );
not ( n16775 , n13861 );
buf ( n16776 , n16772 );
nand ( n16777 , n16775 , n16776 );
and ( n16778 , n16774 , n16777 );
xor ( n16779 , n16771 , n16778 );
buf ( n16780 , n5809 );
nand ( n16781 , n8176 , n16780 );
buf ( n16782 , n5810 );
buf ( n16783 , n16782 );
and ( n16784 , n16781 , n16783 );
not ( n16785 , n16781 );
not ( n16786 , n16782 );
and ( n16787 , n16785 , n16786 );
nor ( n16788 , n16784 , n16787 );
not ( n16789 , n16788 );
buf ( n16790 , n5811 );
not ( n16791 , n16790 );
and ( n16792 , n16789 , n16791 );
and ( n16793 , n16788 , n16790 );
nor ( n16794 , n16792 , n16793 );
xnor ( n16795 , n16779 , n16794 );
not ( n16796 , n16795 );
not ( n16797 , n16796 );
or ( n16798 , n16769 , n16797 );
or ( n16799 , n16796 , n11710 );
nand ( n16800 , n16798 , n16799 );
buf ( n16801 , n12651 );
and ( n16802 , n16800 , n16801 );
not ( n16803 , n16800 );
buf ( n16804 , n10666 );
and ( n16805 , n16803 , n16804 );
nor ( n16806 , n16802 , n16805 );
not ( n16807 , n16806 );
not ( n16808 , n15877 );
buf ( n16809 , n5812 );
not ( n16810 , n16809 );
not ( n16811 , n16810 );
or ( n16812 , n16808 , n16811 );
not ( n16813 , n15876 );
buf ( n16814 , n16809 );
nand ( n16815 , n16813 , n16814 );
nand ( n16816 , n16812 , n16815 );
buf ( n16817 , n5813 );
buf ( n16818 , n16817 );
and ( n16819 , n16816 , n16818 );
not ( n16820 , n16816 );
not ( n16821 , n16817 );
and ( n16822 , n16820 , n16821 );
nor ( n16823 , n16819 , n16822 );
buf ( n16824 , n5814 );
nand ( n16825 , n6577 , n16824 );
buf ( n16826 , n5815 );
xor ( n16827 , n16825 , n16826 );
xor ( n16828 , n16823 , n16827 );
buf ( n16829 , n5816 );
nand ( n16830 , n7569 , n16829 );
buf ( n16831 , n5817 );
buf ( n16832 , n16831 );
and ( n16833 , n16830 , n16832 );
not ( n16834 , n16830 );
not ( n16835 , n16831 );
and ( n16836 , n16834 , n16835 );
nor ( n16837 , n16833 , n16836 );
xnor ( n16838 , n16828 , n16837 );
not ( n16839 , n16838 );
not ( n16840 , n13929 );
and ( n16841 , n16839 , n16840 );
and ( n16842 , n16838 , n13929 );
nor ( n16843 , n16841 , n16842 );
buf ( n16844 , n5818 );
buf ( n16845 , n16844 );
not ( n16846 , n16845 );
buf ( n16847 , n5819 );
not ( n16848 , n16847 );
not ( n16849 , n16848 );
or ( n16850 , n16846 , n16849 );
not ( n16851 , n16844 );
buf ( n16852 , n16847 );
nand ( n16853 , n16851 , n16852 );
nand ( n16854 , n16850 , n16853 );
buf ( n16855 , n5820 );
buf ( n16856 , n16855 );
and ( n16857 , n16854 , n16856 );
not ( n16858 , n16854 );
not ( n16859 , n16855 );
and ( n16860 , n16858 , n16859 );
nor ( n16861 , n16857 , n16860 );
buf ( n16862 , n5821 );
nand ( n16863 , n8364 , n16862 );
buf ( n16864 , n5822 );
buf ( n16865 , n16864 );
and ( n16866 , n16863 , n16865 );
not ( n16867 , n16863 );
not ( n16868 , n16864 );
and ( n16869 , n16867 , n16868 );
nor ( n16870 , n16866 , n16869 );
xor ( n16871 , n16861 , n16870 );
buf ( n16872 , n5823 );
nand ( n16873 , n8125 , n16872 );
buf ( n16874 , n5824 );
not ( n16875 , n16874 );
and ( n16876 , n16873 , n16875 );
not ( n16877 , n16873 );
buf ( n16878 , n16874 );
and ( n16879 , n16877 , n16878 );
nor ( n16880 , n16876 , n16879 );
xnor ( n16881 , n16871 , n16880 );
buf ( n16882 , n16881 );
xor ( n16883 , n16843 , n16882 );
buf ( n16884 , n16883 );
nand ( n16885 , n16807 , n16884 );
not ( n16886 , n16885 );
or ( n16887 , n16768 , n16886 );
or ( n16888 , n16885 , n16767 );
nand ( n16889 , n16887 , n16888 );
not ( n16890 , n16889 );
buf ( n16891 , n15087 );
not ( n16892 , n16891 );
not ( n16893 , n14507 );
or ( n16894 , n16892 , n16893 );
not ( n16895 , n15701 );
or ( n16896 , n16895 , n16891 );
nand ( n16897 , n16894 , n16896 );
buf ( n16898 , n15748 );
and ( n16899 , n16897 , n16898 );
not ( n16900 , n16897 );
and ( n16901 , n16900 , n15751 );
nor ( n16902 , n16899 , n16901 );
not ( n16903 , n11974 );
xor ( n16904 , n10803 , n10822 );
not ( n16905 , n10812 );
xnor ( n16906 , n16904 , n16905 );
not ( n16907 , n16906 );
not ( n16908 , n16907 );
or ( n16909 , n16903 , n16908 );
not ( n16910 , n10824 );
or ( n16911 , n16910 , n11974 );
nand ( n16912 , n16909 , n16911 );
not ( n16913 , n14309 );
not ( n16914 , n16913 );
and ( n16915 , n16912 , n16914 );
not ( n16916 , n16912 );
not ( n16917 , n16914 );
and ( n16918 , n16916 , n16917 );
nor ( n16919 , n16915 , n16918 );
buf ( n16920 , n16919 );
nand ( n16921 , n16902 , n16920 );
not ( n16922 , n16921 );
not ( n16923 , n16055 );
not ( n16924 , n14175 );
or ( n16925 , n16923 , n16924 );
or ( n16926 , n14175 , n16055 );
nand ( n16927 , n16925 , n16926 );
and ( n16928 , n16927 , n14153 );
not ( n16929 , n16927 );
and ( n16930 , n16929 , n14152 );
nor ( n16931 , n16928 , n16930 );
not ( n16932 , n16931 );
not ( n16933 , n16932 );
and ( n16934 , n16922 , n16933 );
and ( n16935 , n16921 , n16932 );
nor ( n16936 , n16934 , n16935 );
not ( n16937 , n16936 );
and ( n16938 , n16890 , n16937 );
and ( n16939 , n16889 , n16936 );
nor ( n16940 , n16938 , n16939 );
and ( n16941 , n16712 , n16940 );
not ( n16942 , n16712 );
not ( n16943 , n16940 );
and ( n16944 , n16942 , n16943 );
nor ( n16945 , n16941 , n16944 );
buf ( n16946 , n16945 );
and ( n16947 , n16289 , n16946 );
not ( n16948 , n16289 );
not ( n16949 , n16946 );
and ( n16950 , n16948 , n16949 );
nor ( n16951 , n16947 , n16950 );
not ( n16952 , n16951 );
not ( n16953 , n15444 );
buf ( n16954 , n5825 );
buf ( n16955 , n16954 );
not ( n16956 , n16955 );
buf ( n16957 , n5826 );
not ( n16958 , n16957 );
not ( n16959 , n16958 );
or ( n16960 , n16956 , n16959 );
not ( n16961 , n16954 );
buf ( n16962 , n16957 );
nand ( n16963 , n16961 , n16962 );
nand ( n16964 , n16960 , n16963 );
buf ( n16965 , n5827 );
buf ( n16966 , n16965 );
and ( n16967 , n16964 , n16966 );
not ( n16968 , n16964 );
not ( n16969 , n16965 );
and ( n16970 , n16968 , n16969 );
nor ( n16971 , n16967 , n16970 );
xor ( n16972 , n16971 , n16551 );
buf ( n16973 , n5828 );
nand ( n16974 , n6605 , n16973 );
buf ( n16975 , n5829 );
not ( n16976 , n16975 );
and ( n16977 , n16974 , n16976 );
not ( n16978 , n16974 );
buf ( n16979 , n16975 );
and ( n16980 , n16978 , n16979 );
nor ( n16981 , n16977 , n16980 );
xnor ( n16982 , n16972 , n16981 );
buf ( n16983 , n16982 );
not ( n16984 , n16983 );
not ( n16985 , n16984 );
or ( n16986 , n16953 , n16985 );
or ( n16987 , n16984 , n15444 );
nand ( n16988 , n16986 , n16987 );
buf ( n16989 , n15762 );
xor ( n16990 , n16989 , n15774 );
xnor ( n16991 , n16990 , n15790 );
not ( n16992 , n16991 );
not ( n16993 , n16992 );
and ( n16994 , n16988 , n16993 );
not ( n16995 , n16988 );
and ( n16996 , n16995 , n16992 );
nor ( n16997 , n16994 , n16996 );
not ( n16998 , n16997 );
nand ( n16999 , n16998 , n10964 );
not ( n17000 , n16999 );
not ( n17001 , n14889 );
buf ( n17002 , n5830 );
buf ( n17003 , n17002 );
not ( n17004 , n17003 );
buf ( n17005 , n5831 );
not ( n17006 , n17005 );
not ( n17007 , n17006 );
or ( n17008 , n17004 , n17007 );
not ( n17009 , n17002 );
buf ( n17010 , n17005 );
nand ( n17011 , n17009 , n17010 );
nand ( n17012 , n17008 , n17011 );
buf ( n17013 , n5832 );
not ( n17014 , n17013 );
and ( n17015 , n17012 , n17014 );
not ( n17016 , n17012 );
buf ( n17017 , n17013 );
and ( n17018 , n17016 , n17017 );
nor ( n17019 , n17015 , n17018 );
buf ( n17020 , n5833 );
nand ( n17021 , n8454 , n17020 );
buf ( n17022 , n5834 );
buf ( n17023 , n17022 );
and ( n17024 , n17021 , n17023 );
not ( n17025 , n17021 );
not ( n17026 , n17022 );
and ( n17027 , n17025 , n17026 );
nor ( n17028 , n17024 , n17027 );
xor ( n17029 , n17019 , n17028 );
buf ( n17030 , n5835 );
nand ( n17031 , n6634 , n17030 );
buf ( n17032 , n5836 );
not ( n17033 , n17032 );
and ( n17034 , n17031 , n17033 );
not ( n17035 , n17031 );
buf ( n17036 , n17032 );
and ( n17037 , n17035 , n17036 );
nor ( n17038 , n17034 , n17037 );
xnor ( n17039 , n17029 , n17038 );
buf ( n17040 , n17039 );
not ( n17041 , n17040 );
or ( n17042 , n17001 , n17041 );
not ( n17043 , n17039 );
not ( n17044 , n17043 );
or ( n17045 , n17044 , n14889 );
nand ( n17046 , n17042 , n17045 );
buf ( n17047 , n5837 );
buf ( n17048 , n17047 );
not ( n17049 , n17048 );
buf ( n17050 , n5838 );
not ( n17051 , n17050 );
not ( n17052 , n17051 );
or ( n17053 , n17049 , n17052 );
not ( n17054 , n17047 );
buf ( n17055 , n17050 );
nand ( n17056 , n17054 , n17055 );
nand ( n17057 , n17053 , n17056 );
buf ( n17058 , n5839 );
not ( n17059 , n17058 );
and ( n17060 , n17057 , n17059 );
not ( n17061 , n17057 );
buf ( n17062 , n17058 );
and ( n17063 , n17061 , n17062 );
nor ( n17064 , n17060 , n17063 );
buf ( n17065 , n5840 );
nand ( n17066 , n7202 , n17065 );
buf ( n17067 , n5841 );
buf ( n17068 , n17067 );
and ( n17069 , n17066 , n17068 );
not ( n17070 , n17066 );
not ( n17071 , n17067 );
and ( n17072 , n17070 , n17071 );
nor ( n17073 , n17069 , n17072 );
xor ( n17074 , n17064 , n17073 );
buf ( n17075 , n5842 );
nand ( n17076 , n11946 , n17075 );
buf ( n17077 , n5843 );
buf ( n17078 , n17077 );
and ( n17079 , n17076 , n17078 );
not ( n17080 , n17076 );
not ( n17081 , n17077 );
and ( n17082 , n17080 , n17081 );
nor ( n17083 , n17079 , n17082 );
xnor ( n17084 , n17074 , n17083 );
not ( n17085 , n17084 );
buf ( n17086 , n17085 );
xor ( n17087 , n17046 , n17086 );
not ( n17088 , n17087 );
not ( n17089 , n17088 );
and ( n17090 , n17000 , n17089 );
and ( n17091 , n16999 , n17088 );
nor ( n17092 , n17090 , n17091 );
buf ( n17093 , n17092 );
not ( n17094 , n17093 );
buf ( n17095 , n5844 );
not ( n17096 , n17095 );
not ( n17097 , n17096 );
not ( n17098 , n15143 );
not ( n17099 , n17098 );
or ( n17100 , n17097 , n17099 );
not ( n17101 , n15144 );
or ( n17102 , n17101 , n17096 );
nand ( n17103 , n17100 , n17102 );
buf ( n17104 , n15187 );
not ( n17105 , n17104 );
and ( n17106 , n17103 , n17105 );
not ( n17107 , n17103 );
and ( n17108 , n17107 , n17104 );
nor ( n17109 , n17106 , n17108 );
buf ( n17110 , n13642 );
xor ( n17111 , n13661 , n13665 );
xnor ( n17112 , n17111 , n13675 );
not ( n17113 , n17112 );
not ( n17114 , n17113 );
buf ( n17115 , n5845 );
buf ( n17116 , n17115 );
not ( n17117 , n17116 );
and ( n17118 , n17114 , n17117 );
and ( n17119 , n13690 , n17116 );
nor ( n17120 , n17118 , n17119 );
not ( n17121 , n17120 );
xor ( n17122 , n17110 , n17121 );
not ( n17123 , n17122 );
nand ( n17124 , n17109 , n17123 );
not ( n17125 , n10589 );
and ( n17126 , n17124 , n17125 );
not ( n17127 , n17124 );
and ( n17128 , n17127 , n10589 );
nor ( n17129 , n17126 , n17128 );
not ( n17130 , n17129 );
not ( n17131 , n17130 );
not ( n17132 , n11094 );
buf ( n17133 , n5846 );
buf ( n17134 , n17133 );
not ( n17135 , n17134 );
buf ( n17136 , n9861 );
xor ( n17137 , n9893 , n17136 );
buf ( n17138 , n9871 );
xnor ( n17139 , n17137 , n17138 );
not ( n17140 , n17139 );
or ( n17141 , n17135 , n17140 );
not ( n17142 , n17134 );
nand ( n17143 , n17142 , n9898 );
nand ( n17144 , n17141 , n17143 );
not ( n17145 , n9940 );
buf ( n17146 , n17145 );
and ( n17147 , n17144 , n17146 );
not ( n17148 , n17144 );
and ( n17149 , n17148 , n9942 );
nor ( n17150 , n17147 , n17149 );
not ( n17151 , n8803 );
buf ( n17152 , n5847 );
buf ( n17153 , n17152 );
not ( n17154 , n17153 );
buf ( n17155 , n5848 );
not ( n17156 , n17155 );
not ( n17157 , n17156 );
or ( n17158 , n17154 , n17157 );
not ( n17159 , n17152 );
buf ( n17160 , n17155 );
nand ( n17161 , n17159 , n17160 );
nand ( n17162 , n17158 , n17161 );
buf ( n17163 , n5849 );
buf ( n17164 , n17163 );
and ( n17165 , n17162 , n17164 );
not ( n17166 , n17162 );
not ( n17167 , n17163 );
and ( n17168 , n17166 , n17167 );
nor ( n17169 , n17165 , n17168 );
buf ( n17170 , n5850 );
nand ( n17171 , n6634 , n17170 );
buf ( n17172 , n5851 );
buf ( n17173 , n17172 );
and ( n17174 , n17171 , n17173 );
not ( n17175 , n17171 );
not ( n17176 , n17172 );
and ( n17177 , n17175 , n17176 );
nor ( n17178 , n17174 , n17177 );
xor ( n17179 , n17169 , n17178 );
buf ( n17180 , n5852 );
nand ( n17181 , n8323 , n17180 );
buf ( n17182 , n5853 );
buf ( n17183 , n17182 );
and ( n17184 , n17181 , n17183 );
not ( n17185 , n17181 );
not ( n17186 , n17182 );
and ( n17187 , n17185 , n17186 );
nor ( n17188 , n17184 , n17187 );
buf ( n17189 , n17188 );
xnor ( n17190 , n17179 , n17189 );
not ( n17191 , n17190 );
or ( n17192 , n17151 , n17191 );
or ( n17193 , n17190 , n8803 );
nand ( n17194 , n17192 , n17193 );
buf ( n17195 , n5854 );
buf ( n17196 , n17195 );
not ( n17197 , n17196 );
buf ( n17198 , n5855 );
not ( n17199 , n17198 );
not ( n17200 , n17199 );
or ( n17201 , n17197 , n17200 );
not ( n17202 , n17195 );
buf ( n17203 , n17198 );
nand ( n17204 , n17202 , n17203 );
nand ( n17205 , n17201 , n17204 );
buf ( n17206 , n5856 );
buf ( n17207 , n17206 );
and ( n17208 , n17205 , n17207 );
not ( n17209 , n17205 );
not ( n17210 , n17206 );
and ( n17211 , n17209 , n17210 );
nor ( n17212 , n17208 , n17211 );
buf ( n17213 , n5857 );
nand ( n17214 , n7977 , n17213 );
buf ( n17215 , n5858 );
buf ( n17216 , n17215 );
and ( n17217 , n17214 , n17216 );
not ( n17218 , n17214 );
not ( n17219 , n17215 );
and ( n17220 , n17218 , n17219 );
nor ( n17221 , n17217 , n17220 );
xor ( n17222 , n17212 , n17221 );
buf ( n17223 , n5859 );
nand ( n17224 , n7355 , n17223 );
buf ( n17225 , n5860 );
buf ( n17226 , n17225 );
and ( n17227 , n17224 , n17226 );
not ( n17228 , n17224 );
not ( n17229 , n17225 );
and ( n17230 , n17228 , n17229 );
nor ( n17231 , n17227 , n17230 );
not ( n17232 , n17231 );
xor ( n17233 , n17222 , n17232 );
not ( n17234 , n17233 );
not ( n17235 , n17234 );
and ( n17236 , n17194 , n17235 );
not ( n17237 , n17194 );
buf ( n17238 , n17233 );
not ( n17239 , n17238 );
and ( n17240 , n17237 , n17239 );
nor ( n17241 , n17236 , n17240 );
nand ( n17242 , n17150 , n17241 );
not ( n17243 , n17242 );
or ( n17244 , n17132 , n17243 );
or ( n17245 , n17242 , n11094 );
nand ( n17246 , n17244 , n17245 );
not ( n17247 , n15603 );
not ( n17248 , n15633 );
not ( n17249 , n6479 );
and ( n17250 , n17248 , n17249 );
and ( n17251 , n15633 , n6479 );
nor ( n17252 , n17250 , n17251 );
and ( n17253 , n17247 , n17252 );
not ( n17254 , n17247 );
not ( n17255 , n17252 );
and ( n17256 , n17254 , n17255 );
nor ( n17257 , n17253 , n17256 );
not ( n17258 , n16881 );
not ( n17259 , n17258 );
not ( n17260 , n13915 );
not ( n17261 , n17260 );
xor ( n17262 , n16823 , n16827 );
xor ( n17263 , n17262 , n16837 );
not ( n17264 , n17263 );
or ( n17265 , n17261 , n17264 );
or ( n17266 , n17263 , n17260 );
nand ( n17267 , n17265 , n17266 );
not ( n17268 , n17267 );
or ( n17269 , n17259 , n17268 );
or ( n17270 , n17267 , n17258 );
nand ( n17271 , n17269 , n17270 );
nand ( n17272 , n17257 , n17271 );
not ( n17273 , n17272 );
not ( n17274 , n11278 );
and ( n17275 , n17273 , n17274 );
and ( n17276 , n17272 , n11278 );
nor ( n17277 , n17275 , n17276 );
nor ( n17278 , n17246 , n17277 );
not ( n17279 , n17278 );
nand ( n17280 , n17246 , n17277 );
nand ( n17281 , n17279 , n17280 );
not ( n17282 , n17281 );
and ( n17283 , n17131 , n17282 );
and ( n17284 , n17130 , n17281 );
nor ( n17285 , n17283 , n17284 );
not ( n17286 , n17285 );
not ( n17287 , n17286 );
nand ( n17288 , n16997 , n17087 );
not ( n17289 , n17288 );
not ( n17290 , n10870 );
and ( n17291 , n17289 , n17290 );
and ( n17292 , n17288 , n10870 );
nor ( n17293 , n17291 , n17292 );
not ( n17294 , n17293 );
buf ( n17295 , n8246 );
not ( n17296 , n17295 );
buf ( n17297 , n5861 );
buf ( n17298 , n17297 );
not ( n17299 , n17298 );
not ( n17300 , n12406 );
not ( n17301 , n17300 );
or ( n17302 , n17299 , n17301 );
not ( n17303 , n17297 );
nand ( n17304 , n17303 , n12407 );
nand ( n17305 , n17302 , n17304 );
buf ( n17306 , n5862 );
not ( n17307 , n17306 );
and ( n17308 , n17305 , n17307 );
not ( n17309 , n17305 );
buf ( n17310 , n17306 );
and ( n17311 , n17309 , n17310 );
nor ( n17312 , n17308 , n17311 );
buf ( n17313 , n5863 );
nand ( n17314 , n7563 , n17313 );
buf ( n17315 , n5864 );
buf ( n17316 , n17315 );
and ( n17317 , n17314 , n17316 );
not ( n17318 , n17314 );
not ( n17319 , n17315 );
and ( n17320 , n17318 , n17319 );
nor ( n17321 , n17317 , n17320 );
xor ( n17322 , n17312 , n17321 );
buf ( n17323 , n5865 );
nand ( n17324 , n6515 , n17323 );
buf ( n17325 , n5866 );
not ( n17326 , n17325 );
and ( n17327 , n17324 , n17326 );
not ( n17328 , n17324 );
buf ( n17329 , n17325 );
and ( n17330 , n17328 , n17329 );
nor ( n17331 , n17327 , n17330 );
xnor ( n17332 , n17322 , n17331 );
buf ( n17333 , n17332 );
not ( n17334 , n17333 );
or ( n17335 , n17296 , n17334 );
not ( n17336 , n17321 );
not ( n17337 , n17331 );
or ( n17338 , n17336 , n17337 );
or ( n17339 , n17321 , n17331 );
nand ( n17340 , n17338 , n17339 );
not ( n17341 , n17312 );
and ( n17342 , n17340 , n17341 );
not ( n17343 , n17340 );
and ( n17344 , n17343 , n17312 );
nor ( n17345 , n17342 , n17344 );
not ( n17346 , n17345 );
not ( n17347 , n17346 );
nand ( n17348 , n17347 , n8247 );
nand ( n17349 , n17335 , n17348 );
and ( n17350 , n17349 , n8996 );
not ( n17351 , n17349 );
and ( n17352 , n17351 , n8992 );
nor ( n17353 , n17350 , n17352 );
not ( n17354 , n17353 );
buf ( n17355 , n5867 );
buf ( n17356 , n17355 );
xor ( n17357 , n12185 , n12195 );
xnor ( n17358 , n17357 , n12205 );
buf ( n17359 , n17358 );
xor ( n17360 , n17356 , n17359 );
not ( n17361 , n12236 );
xnor ( n17362 , n17360 , n17361 );
nand ( n17363 , n17354 , n17362 );
not ( n17364 , n10757 );
and ( n17365 , n17363 , n17364 );
not ( n17366 , n17363 );
and ( n17367 , n17366 , n10757 );
nor ( n17368 , n17365 , n17367 );
not ( n17369 , n17368 );
or ( n17370 , n17294 , n17369 );
or ( n17371 , n17368 , n17293 );
nand ( n17372 , n17370 , n17371 );
not ( n17373 , n17372 );
not ( n17374 , n17373 );
or ( n17375 , n17287 , n17374 );
nand ( n17376 , n17285 , n17372 );
nand ( n17377 , n17375 , n17376 );
not ( n17378 , n17377 );
or ( n17379 , n17094 , n17378 );
or ( n17380 , n17377 , n17093 );
nand ( n17381 , n17379 , n17380 );
xor ( n17382 , n8895 , n8904 );
xnor ( n17383 , n17382 , n8912 );
xor ( n17384 , n9784 , n17383 );
buf ( n17385 , n5868 );
buf ( n17386 , n17385 );
not ( n17387 , n17386 );
buf ( n17388 , n5869 );
not ( n17389 , n17388 );
not ( n17390 , n17389 );
or ( n17391 , n17387 , n17390 );
not ( n17392 , n17385 );
buf ( n17393 , n17388 );
nand ( n17394 , n17392 , n17393 );
nand ( n17395 , n17391 , n17394 );
not ( n17396 , n17115 );
and ( n17397 , n17395 , n17396 );
not ( n17398 , n17395 );
and ( n17399 , n17398 , n17116 );
nor ( n17400 , n17397 , n17399 );
xor ( n17401 , n17400 , n13686 );
buf ( n17402 , n5870 );
nand ( n17403 , n11688 , n17402 );
buf ( n17404 , n5871 );
not ( n17405 , n17404 );
and ( n17406 , n17403 , n17405 );
not ( n17407 , n17403 );
buf ( n17408 , n17404 );
and ( n17409 , n17407 , n17408 );
nor ( n17410 , n17406 , n17409 );
xnor ( n17411 , n17401 , n17410 );
not ( n17412 , n17411 );
xnor ( n17413 , n17384 , n17412 );
not ( n17414 , n17238 );
buf ( n17415 , n8824 );
not ( n17416 , n17415 );
xor ( n17417 , n17169 , n17188 );
not ( n17418 , n17178 );
xnor ( n17419 , n17417 , n17418 );
not ( n17420 , n17419 );
or ( n17421 , n17416 , n17420 );
or ( n17422 , n17419 , n17415 );
nand ( n17423 , n17421 , n17422 );
not ( n17424 , n17423 );
or ( n17425 , n17414 , n17424 );
buf ( n17426 , n17233 );
or ( n17427 , n17423 , n17426 );
nand ( n17428 , n17425 , n17427 );
nand ( n17429 , n17413 , n17428 );
not ( n17430 , n17429 );
not ( n17431 , n15856 );
not ( n17432 , n7539 );
or ( n17433 , n17431 , n17432 );
not ( n17434 , n15856 );
nand ( n17435 , n17434 , n8985 );
nand ( n17436 , n17433 , n17435 );
and ( n17437 , n17436 , n7580 );
not ( n17438 , n17436 );
not ( n17439 , n7580 );
and ( n17440 , n17438 , n17439 );
nor ( n17441 , n17437 , n17440 );
not ( n17442 , n17441 );
not ( n17443 , n17442 );
and ( n17444 , n17430 , n17443 );
and ( n17445 , n17429 , n17442 );
nor ( n17446 , n17444 , n17445 );
not ( n17447 , n13006 );
not ( n17448 , n14091 );
and ( n17449 , n17447 , n17448 );
and ( n17450 , n13006 , n14091 );
nor ( n17451 , n17449 , n17450 );
not ( n17452 , n16341 );
xor ( n17453 , n17452 , n16350 );
xnor ( n17454 , n17453 , n16357 );
buf ( n17455 , n17454 );
and ( n17456 , n17451 , n17455 );
not ( n17457 , n17451 );
and ( n17458 , n17457 , n16359 );
nor ( n17459 , n17456 , n17458 );
not ( n17460 , n9715 );
not ( n17461 , n6525 );
or ( n17462 , n17460 , n17461 );
or ( n17463 , n6525 , n9715 );
nand ( n17464 , n17462 , n17463 );
and ( n17465 , n17464 , n6572 );
not ( n17466 , n17464 );
and ( n17467 , n17466 , n16381 );
nor ( n17468 , n17465 , n17467 );
nor ( n17469 , n17459 , n17468 );
not ( n17470 , n17469 );
not ( n17471 , n10616 );
buf ( n17472 , n5872 );
buf ( n17473 , n17472 );
not ( n17474 , n17473 );
not ( n17475 , n12651 );
or ( n17476 , n17474 , n17475 );
or ( n17477 , n12651 , n17473 );
nand ( n17478 , n17476 , n17477 );
not ( n17479 , n17478 );
and ( n17480 , n17471 , n17479 );
and ( n17481 , n10616 , n17478 );
nor ( n17482 , n17480 , n17481 );
not ( n17483 , n17482 );
or ( n17484 , n17470 , n17483 );
not ( n17485 , n17469 );
not ( n17486 , n17482 );
nand ( n17487 , n17485 , n17486 );
nand ( n17488 , n17484 , n17487 );
xor ( n17489 , n17446 , n17488 );
not ( n17490 , n16992 );
buf ( n17491 , n15468 );
not ( n17492 , n17491 );
not ( n17493 , n16982 );
not ( n17494 , n17493 );
or ( n17495 , n17492 , n17494 );
not ( n17496 , n17491 );
nand ( n17497 , n17496 , n16983 );
nand ( n17498 , n17495 , n17497 );
not ( n17499 , n17498 );
and ( n17500 , n17490 , n17499 );
not ( n17501 , n16991 );
and ( n17502 , n17501 , n17498 );
nor ( n17503 , n17500 , n17502 );
not ( n17504 , n17503 );
buf ( n17505 , n7796 );
not ( n17506 , n17505 );
buf ( n17507 , n5873 );
buf ( n17508 , n17507 );
not ( n17509 , n17508 );
buf ( n17510 , n5874 );
not ( n17511 , n17510 );
not ( n17512 , n17511 );
or ( n17513 , n17509 , n17512 );
not ( n17514 , n17507 );
buf ( n17515 , n17510 );
nand ( n17516 , n17514 , n17515 );
nand ( n17517 , n17513 , n17516 );
buf ( n17518 , n5875 );
not ( n17519 , n17518 );
and ( n17520 , n17517 , n17519 );
not ( n17521 , n17517 );
buf ( n17522 , n17518 );
and ( n17523 , n17521 , n17522 );
nor ( n17524 , n17520 , n17523 );
buf ( n17525 , n5876 );
nand ( n17526 , n7247 , n17525 );
buf ( n17527 , n5877 );
buf ( n17528 , n17527 );
and ( n17529 , n17526 , n17528 );
not ( n17530 , n17526 );
not ( n17531 , n17527 );
and ( n17532 , n17530 , n17531 );
nor ( n17533 , n17529 , n17532 );
xor ( n17534 , n17524 , n17533 );
buf ( n17535 , n5878 );
nand ( n17536 , n7709 , n17535 );
buf ( n17537 , n5879 );
buf ( n17538 , n17537 );
and ( n17539 , n17536 , n17538 );
not ( n17540 , n17536 );
not ( n17541 , n17537 );
and ( n17542 , n17540 , n17541 );
nor ( n17543 , n17539 , n17542 );
xnor ( n17544 , n17534 , n17543 );
buf ( n17545 , n17544 );
not ( n17546 , n17545 );
not ( n17547 , n17546 );
or ( n17548 , n17506 , n17547 );
not ( n17549 , n17505 );
nand ( n17550 , n17549 , n17545 );
nand ( n17551 , n17548 , n17550 );
buf ( n17552 , n5880 );
buf ( n17553 , n17552 );
not ( n17554 , n17553 );
buf ( n17555 , n5881 );
not ( n17556 , n17555 );
not ( n17557 , n17556 );
or ( n17558 , n17554 , n17557 );
not ( n17559 , n17552 );
buf ( n17560 , n17555 );
nand ( n17561 , n17559 , n17560 );
nand ( n17562 , n17558 , n17561 );
and ( n17563 , n17562 , n8890 );
not ( n17564 , n17562 );
not ( n17565 , n8889 );
and ( n17566 , n17564 , n17565 );
nor ( n17567 , n17563 , n17566 );
buf ( n17568 , n5882 );
nand ( n17569 , n8375 , n17568 );
buf ( n17570 , n5883 );
not ( n17571 , n17570 );
and ( n17572 , n17569 , n17571 );
not ( n17573 , n17569 );
buf ( n17574 , n17570 );
and ( n17575 , n17573 , n17574 );
nor ( n17576 , n17572 , n17575 );
not ( n17577 , n17576 );
xor ( n17578 , n17567 , n17577 );
buf ( n17579 , n5884 );
nand ( n17580 , n11688 , n17579 );
buf ( n17581 , n5885 );
buf ( n17582 , n17581 );
and ( n17583 , n17580 , n17582 );
not ( n17584 , n17580 );
not ( n17585 , n17581 );
and ( n17586 , n17584 , n17585 );
nor ( n17587 , n17583 , n17586 );
buf ( n17588 , n17587 );
xnor ( n17589 , n17578 , n17588 );
buf ( n17590 , n17589 );
and ( n17591 , n17551 , n17590 );
not ( n17592 , n17551 );
not ( n17593 , n17587 );
not ( n17594 , n17576 );
or ( n17595 , n17593 , n17594 );
or ( n17596 , n17587 , n17576 );
nand ( n17597 , n17595 , n17596 );
and ( n17598 , n17597 , n17567 );
not ( n17599 , n17597 );
not ( n17600 , n17567 );
and ( n17601 , n17599 , n17600 );
nor ( n17602 , n17598 , n17601 );
buf ( n17603 , n17602 );
and ( n17604 , n17592 , n17603 );
nor ( n17605 , n17591 , n17604 );
nand ( n17606 , n17504 , n17605 );
not ( n17607 , n17606 );
buf ( n17608 , n5886 );
buf ( n17609 , n17608 );
not ( n17610 , n17609 );
not ( n17611 , n11858 );
not ( n17612 , n17611 );
or ( n17613 , n17610 , n17612 );
buf ( n17614 , n11858 );
not ( n17615 , n17608 );
nand ( n17616 , n17614 , n17615 );
nand ( n17617 , n17613 , n17616 );
and ( n17618 , n17617 , n13744 );
not ( n17619 , n17617 );
and ( n17620 , n17619 , n13731 );
nor ( n17621 , n17618 , n17620 );
not ( n17622 , n17621 );
and ( n17623 , n17607 , n17622 );
and ( n17624 , n17606 , n17621 );
nor ( n17625 , n17623 , n17624 );
xor ( n17626 , n17489 , n17625 );
not ( n17627 , n17410 );
nor ( n17628 , n17627 , n17112 );
not ( n17629 , n17628 );
not ( n17630 , n17410 );
nand ( n17631 , n17630 , n17112 );
nand ( n17632 , n17629 , n17631 );
and ( n17633 , n17632 , n13643 );
not ( n17634 , n17632 );
not ( n17635 , n13643 );
and ( n17636 , n17634 , n17635 );
nor ( n17637 , n17633 , n17636 );
not ( n17638 , n17637 );
not ( n17639 , n11346 );
buf ( n17640 , n5887 );
buf ( n17641 , n17640 );
not ( n17642 , n17641 );
buf ( n17643 , n5888 );
not ( n17644 , n17643 );
not ( n17645 , n17644 );
or ( n17646 , n17642 , n17645 );
not ( n17647 , n17640 );
buf ( n17648 , n17643 );
nand ( n17649 , n17647 , n17648 );
nand ( n17650 , n17646 , n17649 );
buf ( n17651 , n5889 );
not ( n17652 , n17651 );
and ( n17653 , n17650 , n17652 );
not ( n17654 , n17650 );
buf ( n17655 , n17651 );
and ( n17656 , n17654 , n17655 );
nor ( n17657 , n17653 , n17656 );
buf ( n17658 , n5890 );
nand ( n17659 , n6502 , n17658 );
buf ( n17660 , n5891 );
xor ( n17661 , n17659 , n17660 );
xor ( n17662 , n17657 , n17661 );
buf ( n17663 , n5892 );
nand ( n17664 , n7709 , n17663 );
buf ( n17665 , n5893 );
not ( n17666 , n17665 );
and ( n17667 , n17664 , n17666 );
not ( n17668 , n17664 );
buf ( n17669 , n17665 );
and ( n17670 , n17668 , n17669 );
nor ( n17671 , n17667 , n17670 );
xnor ( n17672 , n17662 , n17671 );
not ( n17673 , n17672 );
or ( n17674 , n17639 , n17673 );
not ( n17675 , n11346 );
not ( n17676 , n17672 );
nand ( n17677 , n17675 , n17676 );
nand ( n17678 , n17674 , n17677 );
and ( n17679 , n17678 , n17333 );
not ( n17680 , n17678 );
and ( n17681 , n17680 , n17347 );
nor ( n17682 , n17679 , n17681 );
not ( n17683 , n17682 );
nand ( n17684 , n17638 , n17683 );
buf ( n17685 , n5894 );
buf ( n17686 , n17685 );
xor ( n17687 , n17686 , n12811 );
buf ( n17688 , n12833 );
xor ( n17689 , n17687 , n17688 );
not ( n17690 , n17689 );
and ( n17691 , n17684 , n17690 );
not ( n17692 , n17684 );
and ( n17693 , n17692 , n17689 );
nor ( n17694 , n17691 , n17693 );
not ( n17695 , n17694 );
not ( n17696 , n17695 );
buf ( n17697 , n5895 );
nand ( n17698 , n11847 , n17697 );
buf ( n17699 , n5896 );
not ( n17700 , n17699 );
and ( n17701 , n17698 , n17700 );
not ( n17702 , n17698 );
buf ( n17703 , n17699 );
and ( n17704 , n17702 , n17703 );
nor ( n17705 , n17701 , n17704 );
buf ( n17706 , n17705 );
not ( n17707 , n15099 );
xor ( n17708 , n17706 , n17707 );
xnor ( n17709 , n17708 , n7993 );
not ( n17710 , n8091 );
buf ( n17711 , n9266 );
nor ( n17712 , n17710 , n17711 );
not ( n17713 , n17712 );
not ( n17714 , n8067 );
xor ( n17715 , n17714 , n8089 );
xnor ( n17716 , n17715 , n8079 );
buf ( n17717 , n17716 );
not ( n17718 , n17717 );
nand ( n17719 , n17711 , n17718 );
nand ( n17720 , n17713 , n17719 );
not ( n17721 , n8140 );
and ( n17722 , n17720 , n17721 );
not ( n17723 , n17720 );
not ( n17724 , n8136 );
and ( n17725 , n17723 , n17724 );
nor ( n17726 , n17722 , n17725 );
not ( n17727 , n17726 );
nand ( n17728 , n17709 , n17727 );
not ( n17729 , n16517 );
buf ( n17730 , n5897 );
buf ( n17731 , n17730 );
not ( n17732 , n17731 );
buf ( n17733 , n5898 );
not ( n17734 , n17733 );
not ( n17735 , n17734 );
or ( n17736 , n17732 , n17735 );
not ( n17737 , n17730 );
buf ( n17738 , n17733 );
nand ( n17739 , n17737 , n17738 );
nand ( n17740 , n17736 , n17739 );
buf ( n17741 , n5899 );
buf ( n17742 , n17741 );
and ( n17743 , n17740 , n17742 );
not ( n17744 , n17740 );
not ( n17745 , n17741 );
and ( n17746 , n17744 , n17745 );
nor ( n17747 , n17743 , n17746 );
buf ( n17748 , n5900 );
nand ( n17749 , n6557 , n17748 );
buf ( n17750 , n5901 );
not ( n17751 , n17750 );
and ( n17752 , n17749 , n17751 );
not ( n17753 , n17749 );
buf ( n17754 , n17750 );
and ( n17755 , n17753 , n17754 );
nor ( n17756 , n17752 , n17755 );
xor ( n17757 , n17747 , n17756 );
buf ( n17758 , n5902 );
nand ( n17759 , n7067 , n17758 );
buf ( n17760 , n5903 );
not ( n17761 , n17760 );
and ( n17762 , n17759 , n17761 );
not ( n17763 , n17759 );
buf ( n17764 , n17760 );
and ( n17765 , n17763 , n17764 );
nor ( n17766 , n17762 , n17765 );
xnor ( n17767 , n17757 , n17766 );
not ( n17768 , n17767 );
not ( n17769 , n17768 );
not ( n17770 , n17769 );
or ( n17771 , n17729 , n17770 );
not ( n17772 , n17767 );
not ( n17773 , n17772 );
or ( n17774 , n17773 , n16517 );
nand ( n17775 , n17771 , n17774 );
not ( n17776 , n14175 );
and ( n17777 , n17775 , n17776 );
not ( n17778 , n17775 );
and ( n17779 , n17778 , n14175 );
nor ( n17780 , n17777 , n17779 );
and ( n17781 , n17728 , n17780 );
not ( n17782 , n17728 );
not ( n17783 , n17780 );
and ( n17784 , n17782 , n17783 );
nor ( n17785 , n17781 , n17784 );
not ( n17786 , n17785 );
not ( n17787 , n17786 );
or ( n17788 , n17696 , n17787 );
nand ( n17789 , n17785 , n17694 );
nand ( n17790 , n17788 , n17789 );
and ( n17791 , n17626 , n17790 );
not ( n17792 , n17626 );
not ( n17793 , n17790 );
and ( n17794 , n17792 , n17793 );
nor ( n17795 , n17791 , n17794 );
not ( n17796 , n17795 );
not ( n17797 , n17796 );
and ( n17798 , n17381 , n17797 );
not ( n17799 , n17381 );
buf ( n17800 , n17795 );
not ( n17801 , n17800 );
and ( n17802 , n17799 , n17801 );
nor ( n17803 , n17798 , n17802 );
not ( n17804 , n17803 );
nand ( n17805 , n16952 , n17804 );
or ( n17806 , n15328 , n17805 );
buf ( n17807 , n13344 );
not ( n17808 , n17807 );
buf ( n17809 , n17808 );
not ( n17810 , n17809 );
nor ( n17811 , n15323 , n17810 );
nand ( n17812 , n17811 , n17805 );
buf ( n17813 , n13353 );
nand ( n17814 , n17813 , n13573 );
nand ( n17815 , n17806 , n17812 , n17814 );
buf ( n17816 , n17815 );
buf ( n17817 , n17816 );
not ( n17818 , n12738 );
buf ( n17819 , n13352 );
buf ( n17820 , n17819 );
not ( n17821 , n17820 );
or ( n17822 , n17818 , n17821 );
buf ( n17823 , n5904 );
buf ( n17824 , n17823 );
not ( n17825 , n17824 );
buf ( n17826 , n5905 );
not ( n17827 , n17826 );
not ( n17828 , n17827 );
or ( n17829 , n17825 , n17828 );
not ( n17830 , n17823 );
buf ( n17831 , n17826 );
nand ( n17832 , n17830 , n17831 );
nand ( n17833 , n17829 , n17832 );
buf ( n17834 , n5906 );
not ( n17835 , n17834 );
and ( n17836 , n17833 , n17835 );
not ( n17837 , n17833 );
buf ( n17838 , n17834 );
and ( n17839 , n17837 , n17838 );
nor ( n17840 , n17836 , n17839 );
buf ( n17841 , n5907 );
nand ( n17842 , n7258 , n17841 );
buf ( n17843 , n5908 );
buf ( n17844 , n17843 );
and ( n17845 , n17842 , n17844 );
not ( n17846 , n17842 );
not ( n17847 , n17843 );
and ( n17848 , n17846 , n17847 );
nor ( n17849 , n17845 , n17848 );
xor ( n17850 , n17840 , n17849 );
buf ( n17851 , n5909 );
nand ( n17852 , n7569 , n17851 );
buf ( n17853 , n5910 );
not ( n17854 , n17853 );
and ( n17855 , n17852 , n17854 );
not ( n17856 , n17852 );
buf ( n17857 , n17853 );
and ( n17858 , n17856 , n17857 );
nor ( n17859 , n17855 , n17858 );
xnor ( n17860 , n17850 , n17859 );
not ( n17861 , n17860 );
not ( n17862 , n17861 );
xor ( n17863 , n14183 , n17862 );
buf ( n17864 , n5911 );
not ( n17865 , n17864 );
buf ( n17866 , n5912 );
not ( n17867 , n17866 );
buf ( n17868 , n5913 );
buf ( n17869 , n17868 );
and ( n17870 , n17867 , n17869 );
not ( n17871 , n17867 );
not ( n17872 , n17868 );
and ( n17873 , n17871 , n17872 );
nor ( n17874 , n17870 , n17873 );
xor ( n17875 , n17865 , n17874 );
buf ( n17876 , n5914 );
buf ( n17877 , n5915 );
xor ( n17878 , n17876 , n17877 );
buf ( n17879 , n5916 );
nand ( n17880 , n6828 , n17879 );
xnor ( n17881 , n17878 , n17880 );
xnor ( n17882 , n17875 , n17881 );
buf ( n17883 , n17882 );
xnor ( n17884 , n17863 , n17883 );
buf ( n17885 , n5917 );
buf ( n17886 , n17885 );
not ( n17887 , n17886 );
not ( n17888 , n12707 );
or ( n17889 , n17887 , n17888 );
not ( n17890 , n17885 );
nand ( n17891 , n12713 , n17890 );
nand ( n17892 , n17889 , n17891 );
not ( n17893 , n12756 );
and ( n17894 , n17892 , n17893 );
not ( n17895 , n17892 );
and ( n17896 , n17895 , n12756 );
nor ( n17897 , n17894 , n17896 );
nand ( n17898 , n17884 , n17897 );
not ( n17899 , n16345 );
not ( n17900 , n13445 );
or ( n17901 , n17899 , n17900 );
xor ( n17902 , n13444 , n13412 );
buf ( n17903 , n13422 );
xnor ( n17904 , n17902 , n17903 );
or ( n17905 , n16345 , n17904 );
nand ( n17906 , n17901 , n17905 );
xor ( n17907 , n13377 , n13386 );
xnor ( n17908 , n17907 , n13397 );
and ( n17909 , n17906 , n17908 );
not ( n17910 , n17906 );
and ( n17911 , n17910 , n13399 );
nor ( n17912 , n17909 , n17911 );
not ( n17913 , n17912 );
and ( n17914 , n17898 , n17913 );
not ( n17915 , n17898 );
and ( n17916 , n17915 , n17912 );
nor ( n17917 , n17914 , n17916 );
not ( n17918 , n17917 );
not ( n17919 , n11747 );
buf ( n17920 , n5918 );
buf ( n17921 , n17920 );
not ( n17922 , n17921 );
buf ( n17923 , n5919 );
not ( n17924 , n17923 );
not ( n17925 , n17924 );
or ( n17926 , n17922 , n17925 );
not ( n17927 , n17920 );
buf ( n17928 , n17923 );
nand ( n17929 , n17927 , n17928 );
nand ( n17930 , n17926 , n17929 );
buf ( n17931 , n5920 );
not ( n17932 , n17931 );
and ( n17933 , n17930 , n17932 );
not ( n17934 , n17930 );
buf ( n17935 , n17931 );
and ( n17936 , n17934 , n17935 );
nor ( n17937 , n17933 , n17936 );
buf ( n17938 , n5921 );
nand ( n17939 , n6828 , n17938 );
buf ( n17940 , n5922 );
buf ( n17941 , n17940 );
and ( n17942 , n17939 , n17941 );
not ( n17943 , n17939 );
not ( n17944 , n17940 );
and ( n17945 , n17943 , n17944 );
nor ( n17946 , n17942 , n17945 );
xor ( n17947 , n17937 , n17946 );
buf ( n17948 , n5923 );
nand ( n17949 , n8675 , n17948 );
buf ( n17950 , n5924 );
not ( n17951 , n17950 );
and ( n17952 , n17949 , n17951 );
not ( n17953 , n17949 );
buf ( n17954 , n17950 );
and ( n17955 , n17953 , n17954 );
nor ( n17956 , n17952 , n17955 );
xnor ( n17957 , n17947 , n17956 );
not ( n17958 , n17957 );
not ( n17959 , n17958 );
not ( n17960 , n17959 );
or ( n17961 , n17919 , n17960 );
not ( n17962 , n11747 );
nand ( n17963 , n17962 , n17958 );
nand ( n17964 , n17961 , n17963 );
buf ( n17965 , n5925 );
buf ( n17966 , n17965 );
not ( n17967 , n17966 );
buf ( n17968 , n5926 );
not ( n17969 , n17968 );
not ( n17970 , n17969 );
or ( n17971 , n17967 , n17970 );
not ( n17972 , n17965 );
buf ( n17973 , n17968 );
nand ( n17974 , n17972 , n17973 );
nand ( n17975 , n17971 , n17974 );
buf ( n17976 , n5927 );
buf ( n17977 , n17976 );
and ( n17978 , n17975 , n17977 );
not ( n17979 , n17975 );
not ( n17980 , n17976 );
and ( n17981 , n17979 , n17980 );
nor ( n17982 , n17978 , n17981 );
buf ( n17983 , n5928 );
nand ( n17984 , n6502 , n17983 );
buf ( n17985 , n5929 );
not ( n17986 , n17985 );
and ( n17987 , n17984 , n17986 );
not ( n17988 , n17984 );
buf ( n17989 , n17985 );
and ( n17990 , n17988 , n17989 );
nor ( n17991 , n17987 , n17990 );
xor ( n17992 , n17982 , n17991 );
buf ( n17993 , n5930 );
nand ( n17994 , n6828 , n17993 );
buf ( n17995 , n5931 );
not ( n17996 , n17995 );
and ( n17997 , n17994 , n17996 );
not ( n17998 , n17994 );
buf ( n17999 , n17995 );
and ( n18000 , n17998 , n17999 );
nor ( n18001 , n17997 , n18000 );
xnor ( n18002 , n17992 , n18001 );
buf ( n18003 , n18002 );
not ( n18004 , n18003 );
and ( n18005 , n17964 , n18004 );
not ( n18006 , n17964 );
and ( n18007 , n18006 , n18003 );
nor ( n18008 , n18005 , n18007 );
not ( n18009 , n18008 );
not ( n18010 , n16036 );
not ( n18011 , n14174 );
or ( n18012 , n18010 , n18011 );
or ( n18013 , n14174 , n16036 );
nand ( n18014 , n18012 , n18013 );
not ( n18015 , n14151 );
and ( n18016 , n18014 , n18015 );
not ( n18017 , n18014 );
and ( n18018 , n18017 , n14152 );
nor ( n18019 , n18016 , n18018 );
not ( n18020 , n8722 );
not ( n18021 , n18020 );
buf ( n18022 , n5932 );
buf ( n18023 , n18022 );
not ( n18024 , n18023 );
and ( n18025 , n18021 , n18024 );
and ( n18026 , n18020 , n18023 );
nor ( n18027 , n18025 , n18026 );
not ( n18028 , n12010 );
and ( n18029 , n18027 , n18028 );
not ( n18030 , n18027 );
and ( n18031 , n18030 , n12011 );
nor ( n18032 , n18029 , n18031 );
nand ( n18033 , n18019 , n18032 );
not ( n18034 , n18033 );
or ( n18035 , n18009 , n18034 );
or ( n18036 , n18033 , n18008 );
nand ( n18037 , n18035 , n18036 );
not ( n18038 , n18037 );
not ( n18039 , n8760 );
not ( n18040 , n18039 );
buf ( n18041 , n5933 );
buf ( n18042 , n18041 );
not ( n18043 , n18042 );
buf ( n18044 , n5934 );
buf ( n18045 , n18044 );
not ( n18046 , n18045 );
buf ( n18047 , n5935 );
not ( n18048 , n18047 );
not ( n18049 , n18048 );
or ( n18050 , n18046 , n18049 );
not ( n18051 , n18044 );
buf ( n18052 , n18047 );
nand ( n18053 , n18051 , n18052 );
nand ( n18054 , n18050 , n18053 );
buf ( n18055 , n5936 );
buf ( n18056 , n18055 );
and ( n18057 , n18054 , n18056 );
not ( n18058 , n18054 );
not ( n18059 , n18055 );
and ( n18060 , n18058 , n18059 );
nor ( n18061 , n18057 , n18060 );
buf ( n18062 , n5937 );
nand ( n18063 , n8323 , n18062 );
buf ( n18064 , n5938 );
buf ( n18065 , n18064 );
and ( n18066 , n18063 , n18065 );
not ( n18067 , n18063 );
not ( n18068 , n18064 );
and ( n18069 , n18067 , n18068 );
nor ( n18070 , n18066 , n18069 );
xor ( n18071 , n18061 , n18070 );
buf ( n18072 , n5939 );
nand ( n18073 , n8675 , n18072 );
buf ( n18074 , n5940 );
buf ( n18075 , n18074 );
and ( n18076 , n18073 , n18075 );
not ( n18077 , n18073 );
not ( n18078 , n18074 );
and ( n18079 , n18077 , n18078 );
nor ( n18080 , n18076 , n18079 );
xnor ( n18081 , n18071 , n18080 );
buf ( n18082 , n18081 );
not ( n18083 , n18082 );
or ( n18084 , n18043 , n18083 );
or ( n18085 , n18082 , n18042 );
nand ( n18086 , n18084 , n18085 );
not ( n18087 , n18086 );
and ( n18088 , n18040 , n18087 );
and ( n18089 , n18039 , n18086 );
nor ( n18090 , n18088 , n18089 );
buf ( n18091 , n5941 );
buf ( n18092 , n18091 );
not ( n18093 , n18092 );
buf ( n18094 , n5942 );
not ( n18095 , n18094 );
not ( n18096 , n18095 );
or ( n18097 , n18093 , n18096 );
not ( n18098 , n18091 );
buf ( n18099 , n18094 );
nand ( n18100 , n18098 , n18099 );
nand ( n18101 , n18097 , n18100 );
xor ( n18102 , n9515 , n18101 );
buf ( n18103 , n5943 );
buf ( n18104 , n5944 );
not ( n18105 , n18104 );
xor ( n18106 , n18103 , n18105 );
buf ( n18107 , n5945 );
nand ( n18108 , n8375 , n18107 );
xnor ( n18109 , n18106 , n18108 );
xnor ( n18110 , n18102 , n18109 );
not ( n18111 , n18110 );
buf ( n18112 , n18111 );
not ( n18113 , n18112 );
buf ( n18114 , n5946 );
buf ( n18115 , n18114 );
not ( n18116 , n18115 );
buf ( n18117 , n5947 );
buf ( n18118 , n18117 );
not ( n18119 , n18118 );
buf ( n18120 , n5948 );
not ( n18121 , n18120 );
not ( n18122 , n18121 );
or ( n18123 , n18119 , n18122 );
not ( n18124 , n18117 );
buf ( n18125 , n18120 );
nand ( n18126 , n18124 , n18125 );
nand ( n18127 , n18123 , n18126 );
buf ( n18128 , n5949 );
buf ( n18129 , n18128 );
and ( n18130 , n18127 , n18129 );
not ( n18131 , n18127 );
not ( n18132 , n18128 );
and ( n18133 , n18131 , n18132 );
nor ( n18134 , n18130 , n18133 );
buf ( n18135 , n5950 );
nand ( n18136 , n6815 , n18135 );
buf ( n18137 , n5951 );
not ( n18138 , n18137 );
and ( n18139 , n18136 , n18138 );
not ( n18140 , n18136 );
buf ( n18141 , n18137 );
and ( n18142 , n18140 , n18141 );
nor ( n18143 , n18139 , n18142 );
xor ( n18144 , n18134 , n18143 );
buf ( n18145 , n5952 );
nand ( n18146 , n7014 , n18145 );
buf ( n18147 , n5953 );
buf ( n18148 , n18147 );
and ( n18149 , n18146 , n18148 );
not ( n18150 , n18146 );
not ( n18151 , n18147 );
and ( n18152 , n18150 , n18151 );
nor ( n18153 , n18149 , n18152 );
xor ( n18154 , n18144 , n18153 );
not ( n18155 , n18154 );
or ( n18156 , n18116 , n18155 );
or ( n18157 , n18154 , n18115 );
nand ( n18158 , n18156 , n18157 );
not ( n18159 , n18158 );
and ( n18160 , n18113 , n18159 );
and ( n18161 , n18112 , n18158 );
nor ( n18162 , n18160 , n18161 );
not ( n18163 , n18162 );
nand ( n18164 , n18090 , n18163 );
not ( n18165 , n18164 );
buf ( n18166 , n8046 );
not ( n18167 , n18166 );
buf ( n18168 , n15947 );
not ( n18169 , n18168 );
buf ( n18170 , n5954 );
buf ( n18171 , n18170 );
not ( n18172 , n18171 );
buf ( n18173 , n5955 );
not ( n18174 , n18173 );
not ( n18175 , n18174 );
or ( n18176 , n18172 , n18175 );
not ( n18177 , n18170 );
buf ( n18178 , n18173 );
nand ( n18179 , n18177 , n18178 );
nand ( n18180 , n18176 , n18179 );
buf ( n18181 , n5956 );
buf ( n18182 , n18181 );
and ( n18183 , n18180 , n18182 );
not ( n18184 , n18180 );
not ( n18185 , n18181 );
and ( n18186 , n18184 , n18185 );
nor ( n18187 , n18183 , n18186 );
buf ( n18188 , n5957 );
nand ( n18189 , n11946 , n18188 );
buf ( n18190 , n5958 );
buf ( n18191 , n18190 );
and ( n18192 , n18189 , n18191 );
not ( n18193 , n18189 );
not ( n18194 , n18190 );
and ( n18195 , n18193 , n18194 );
nor ( n18196 , n18192 , n18195 );
xor ( n18197 , n18187 , n18196 );
buf ( n18198 , n5959 );
nand ( n18199 , n7107 , n18198 );
buf ( n18200 , n5960 );
buf ( n18201 , n18200 );
and ( n18202 , n18199 , n18201 );
not ( n18203 , n18199 );
not ( n18204 , n18200 );
and ( n18205 , n18203 , n18204 );
nor ( n18206 , n18202 , n18205 );
xor ( n18207 , n18197 , n18206 );
not ( n18208 , n18207 );
not ( n18209 , n18208 );
or ( n18210 , n18169 , n18209 );
not ( n18211 , n18168 );
xor ( n18212 , n18187 , n18206 );
not ( n18213 , n18196 );
xnor ( n18214 , n18212 , n18213 );
nand ( n18215 , n18211 , n18214 );
nand ( n18216 , n18210 , n18215 );
not ( n18217 , n18216 );
or ( n18218 , n18167 , n18217 );
or ( n18219 , n18216 , n18166 );
nand ( n18220 , n18218 , n18219 );
not ( n18221 , n18220 );
and ( n18222 , n18165 , n18221 );
and ( n18223 , n18164 , n18220 );
nor ( n18224 , n18222 , n18223 );
not ( n18225 , n18224 );
or ( n18226 , n18038 , n18225 );
or ( n18227 , n18037 , n18224 );
nand ( n18228 , n18226 , n18227 );
not ( n18229 , n17884 );
nand ( n18230 , n18229 , n17913 );
not ( n18231 , n18230 );
not ( n18232 , n7365 );
not ( n18233 , n17233 );
or ( n18234 , n18232 , n18233 );
xor ( n18235 , n17212 , n17231 );
not ( n18236 , n17221 );
xnor ( n18237 , n18235 , n18236 );
nand ( n18238 , n18237 , n7364 );
nand ( n18239 , n18234 , n18238 );
not ( n18240 , n18239 );
buf ( n18241 , n5961 );
buf ( n18242 , n5962 );
buf ( n18243 , n18242 );
not ( n18244 , n18243 );
buf ( n18245 , n5963 );
not ( n18246 , n18245 );
not ( n18247 , n18246 );
or ( n18248 , n18244 , n18247 );
not ( n18249 , n18242 );
buf ( n18250 , n18245 );
nand ( n18251 , n18249 , n18250 );
nand ( n18252 , n18248 , n18251 );
xor ( n18253 , n18241 , n18252 );
buf ( n18254 , n5964 );
buf ( n18255 , n5965 );
xor ( n18256 , n18254 , n18255 );
buf ( n18257 , n5966 );
nand ( n18258 , n8455 , n18257 );
xnor ( n18259 , n18256 , n18258 );
xnor ( n18260 , n18253 , n18259 );
buf ( n18261 , n18260 );
not ( n18262 , n18261 );
and ( n18263 , n18240 , n18262 );
and ( n18264 , n18239 , n18261 );
nor ( n18265 , n18263 , n18264 );
not ( n18266 , n18265 );
not ( n18267 , n18266 );
and ( n18268 , n18231 , n18267 );
and ( n18269 , n18230 , n18266 );
nor ( n18270 , n18268 , n18269 );
not ( n18271 , n18270 );
and ( n18272 , n18228 , n18271 );
not ( n18273 , n18228 );
and ( n18274 , n18273 , n18270 );
nor ( n18275 , n18272 , n18274 );
not ( n18276 , n18275 );
not ( n18277 , n18276 );
not ( n18278 , n11128 );
not ( n18279 , n9788 );
or ( n18280 , n18278 , n18279 );
or ( n18281 , n9788 , n11128 );
nand ( n18282 , n18280 , n18281 );
not ( n18283 , n18282 );
not ( n18284 , n9839 );
or ( n18285 , n18283 , n18284 );
not ( n18286 , n9840 );
or ( n18287 , n18286 , n18282 );
nand ( n18288 , n18285 , n18287 );
not ( n18289 , n18288 );
buf ( n18290 , n5967 );
not ( n18291 , n18290 );
not ( n18292 , n8483 );
xor ( n18293 , n18292 , n8502 );
not ( n18294 , n8492 );
xnor ( n18295 , n18293 , n18294 );
not ( n18296 , n18295 );
not ( n18297 , n18296 );
not ( n18298 , n18297 );
or ( n18299 , n18291 , n18298 );
not ( n18300 , n18296 );
or ( n18301 , n18300 , n18290 );
nand ( n18302 , n18299 , n18301 );
and ( n18303 , n18302 , n8548 );
not ( n18304 , n18302 );
and ( n18305 , n18304 , n8549 );
nor ( n18306 , n18303 , n18305 );
not ( n18307 , n18306 );
nand ( n18308 , n18289 , n18307 );
not ( n18309 , n18308 );
xor ( n18310 , n12931 , n14052 );
buf ( n18311 , n5968 );
buf ( n18312 , n5969 );
not ( n18313 , n18312 );
buf ( n18314 , n5970 );
buf ( n18315 , n18314 );
and ( n18316 , n18313 , n18315 );
not ( n18317 , n18313 );
not ( n18318 , n18314 );
and ( n18319 , n18317 , n18318 );
nor ( n18320 , n18316 , n18319 );
xor ( n18321 , n18311 , n18320 );
buf ( n18322 , n5971 );
xor ( n18323 , n18322 , n10872 );
xnor ( n18324 , n18323 , n10876 );
xnor ( n18325 , n18321 , n18324 );
buf ( n18326 , n18325 );
xnor ( n18327 , n18310 , n18326 );
not ( n18328 , n18327 );
and ( n18329 , n18309 , n18328 );
and ( n18330 , n18308 , n18327 );
nor ( n18331 , n18329 , n18330 );
not ( n18332 , n18331 );
xor ( n18333 , n9579 , n10398 );
xnor ( n18334 , n18333 , n10679 );
buf ( n18335 , n5972 );
buf ( n18336 , n18335 );
not ( n18337 , n18336 );
buf ( n18338 , n5973 );
not ( n18339 , n18338 );
not ( n18340 , n18339 );
or ( n18341 , n18337 , n18340 );
not ( n18342 , n18335 );
buf ( n18343 , n18338 );
nand ( n18344 , n18342 , n18343 );
nand ( n18345 , n18341 , n18344 );
buf ( n18346 , n5974 );
buf ( n18347 , n18346 );
and ( n18348 , n18345 , n18347 );
not ( n18349 , n18345 );
not ( n18350 , n18346 );
and ( n18351 , n18349 , n18350 );
nor ( n18352 , n18348 , n18351 );
buf ( n18353 , n5975 );
nand ( n18354 , n7355 , n18353 );
buf ( n18355 , n5976 );
buf ( n18356 , n18355 );
and ( n18357 , n18354 , n18356 );
not ( n18358 , n18354 );
not ( n18359 , n18355 );
and ( n18360 , n18358 , n18359 );
nor ( n18361 , n18357 , n18360 );
xor ( n18362 , n18352 , n18361 );
buf ( n18363 , n5977 );
nand ( n18364 , n6647 , n18363 );
buf ( n18365 , n5978 );
not ( n18366 , n18365 );
and ( n18367 , n18364 , n18366 );
not ( n18368 , n18364 );
buf ( n18369 , n18365 );
and ( n18370 , n18368 , n18369 );
nor ( n18371 , n18367 , n18370 );
xnor ( n18372 , n18362 , n18371 );
and ( n18373 , n17055 , n18372 );
not ( n18374 , n17055 );
not ( n18375 , n18371 );
xor ( n18376 , n18352 , n18375 );
buf ( n18377 , n18361 );
xor ( n18378 , n18376 , n18377 );
not ( n18379 , n18378 );
and ( n18380 , n18374 , n18379 );
or ( n18381 , n18373 , n18380 );
not ( n18382 , n18381 );
not ( n18383 , n10271 );
or ( n18384 , n18382 , n18383 );
or ( n18385 , n10271 , n18381 );
nand ( n18386 , n18384 , n18385 );
buf ( n18387 , n18386 );
not ( n18388 , n18387 );
nand ( n18389 , n18334 , n18388 );
buf ( n18390 , n5979 );
nand ( n18391 , n8675 , n18390 );
buf ( n18392 , n5980 );
not ( n18393 , n18392 );
and ( n18394 , n18391 , n18393 );
not ( n18395 , n18391 );
buf ( n18396 , n18392 );
and ( n18397 , n18395 , n18396 );
nor ( n18398 , n18394 , n18397 );
buf ( n18399 , n18398 );
not ( n18400 , n18399 );
not ( n18401 , n17139 );
or ( n18402 , n18400 , n18401 );
not ( n18403 , n18399 );
nand ( n18404 , n18403 , n9898 );
nand ( n18405 , n18402 , n18404 );
and ( n18406 , n18405 , n9942 );
not ( n18407 , n18405 );
and ( n18408 , n18407 , n17146 );
nor ( n18409 , n18406 , n18408 );
and ( n18410 , n18389 , n18409 );
not ( n18411 , n18389 );
not ( n18412 , n18409 );
and ( n18413 , n18411 , n18412 );
nor ( n18414 , n18410 , n18413 );
not ( n18415 , n18414 );
or ( n18416 , n18332 , n18415 );
not ( n18417 , n18414 );
not ( n18418 , n18331 );
nand ( n18419 , n18417 , n18418 );
nand ( n18420 , n18416 , n18419 );
not ( n18421 , n18420 );
and ( n18422 , n18277 , n18421 );
and ( n18423 , n18276 , n18420 );
nor ( n18424 , n18422 , n18423 );
not ( n18425 , n18424 );
or ( n18426 , n17918 , n18425 );
not ( n18427 , n17917 );
not ( n18428 , n18275 );
not ( n18429 , n18420 );
not ( n18430 , n18429 );
or ( n18431 , n18428 , n18430 );
nand ( n18432 , n18276 , n18420 );
nand ( n18433 , n18431 , n18432 );
nand ( n18434 , n18427 , n18433 );
nand ( n18435 , n18426 , n18434 );
not ( n18436 , n16057 );
and ( n18437 , n15808 , n18436 );
not ( n18438 , n15808 );
and ( n18439 , n18438 , n16057 );
nor ( n18440 , n18437 , n18439 );
not ( n18441 , n18440 );
and ( n18442 , n16100 , n18441 );
not ( n18443 , n16100 );
and ( n18444 , n18443 , n18440 );
nor ( n18445 , n18442 , n18444 );
buf ( n18446 , n5981 );
nand ( n18447 , n6927 , n18446 );
buf ( n18448 , n5982 );
buf ( n18449 , n18448 );
and ( n18450 , n18447 , n18449 );
not ( n18451 , n18447 );
not ( n18452 , n18448 );
and ( n18453 , n18451 , n18452 );
nor ( n18454 , n18450 , n18453 );
buf ( n18455 , n18454 );
not ( n18456 , n18455 );
not ( n18457 , n15689 );
or ( n18458 , n18456 , n18457 );
xor ( n18459 , n15664 , n15683 );
not ( n18460 , n15673 );
xnor ( n18461 , n18459 , n18460 );
not ( n18462 , n18461 );
or ( n18463 , n18462 , n18455 );
nand ( n18464 , n18458 , n18463 );
buf ( n18465 , n12498 );
and ( n18466 , n18464 , n18465 );
not ( n18467 , n18464 );
and ( n18468 , n18467 , n15692 );
nor ( n18469 , n18466 , n18468 );
not ( n18470 , n18469 );
nand ( n18471 , n18445 , n18470 );
not ( n18472 , n18471 );
buf ( n18473 , n5983 );
buf ( n18474 , n18473 );
buf ( n18475 , n18082 );
xor ( n18476 , n18474 , n18475 );
xnor ( n18477 , n18476 , n7665 );
not ( n18478 , n18477 );
or ( n18479 , n18472 , n18478 );
or ( n18480 , n18477 , n18471 );
nand ( n18481 , n18479 , n18480 );
not ( n18482 , n18481 );
not ( n18483 , n18482 );
not ( n18484 , n12540 );
not ( n18485 , n10126 );
or ( n18486 , n18484 , n18485 );
not ( n18487 , n12540 );
nand ( n18488 , n18487 , n10491 );
nand ( n18489 , n18486 , n18488 );
buf ( n18490 , n5984 );
buf ( n18491 , n18490 );
not ( n18492 , n18491 );
not ( n18493 , n12663 );
not ( n18494 , n18493 );
or ( n18495 , n18492 , n18494 );
not ( n18496 , n18490 );
nand ( n18497 , n18496 , n12664 );
nand ( n18498 , n18495 , n18497 );
not ( n18499 , n18498 );
buf ( n18500 , n5985 );
nand ( n18501 , n7606 , n18500 );
buf ( n18502 , n5986 );
buf ( n18503 , n18502 );
and ( n18504 , n18501 , n18503 );
not ( n18505 , n18501 );
not ( n18506 , n18502 );
and ( n18507 , n18505 , n18506 );
nor ( n18508 , n18504 , n18507 );
xor ( n18509 , n17886 , n18508 );
buf ( n18510 , n5987 );
nand ( n18511 , n7709 , n18510 );
buf ( n18512 , n5988 );
not ( n18513 , n18512 );
and ( n18514 , n18511 , n18513 );
not ( n18515 , n18511 );
buf ( n18516 , n18512 );
and ( n18517 , n18515 , n18516 );
nor ( n18518 , n18514 , n18517 );
xnor ( n18519 , n18509 , n18518 );
not ( n18520 , n18519 );
not ( n18521 , n18520 );
or ( n18522 , n18499 , n18521 );
not ( n18523 , n18498 );
nand ( n18524 , n18523 , n18519 );
nand ( n18525 , n18522 , n18524 );
and ( n18526 , n18489 , n18525 );
not ( n18527 , n18489 );
not ( n18528 , n18525 );
and ( n18529 , n18527 , n18528 );
nor ( n18530 , n18526 , n18529 );
buf ( n18531 , n5989 );
buf ( n18532 , n18531 );
not ( n18533 , n18532 );
buf ( n18534 , n5990 );
not ( n18535 , n18534 );
not ( n18536 , n18535 );
or ( n18537 , n18533 , n18536 );
not ( n18538 , n18531 );
buf ( n18539 , n18534 );
nand ( n18540 , n18538 , n18539 );
nand ( n18541 , n18537 , n18540 );
buf ( n18542 , n5991 );
not ( n18543 , n18542 );
and ( n18544 , n18541 , n18543 );
not ( n18545 , n18541 );
buf ( n18546 , n18542 );
and ( n18547 , n18545 , n18546 );
nor ( n18548 , n18544 , n18547 );
xor ( n18549 , n18548 , n6586 );
buf ( n18550 , n5992 );
nand ( n18551 , n7247 , n18550 );
buf ( n18552 , n5993 );
not ( n18553 , n18552 );
and ( n18554 , n18551 , n18553 );
not ( n18555 , n18551 );
buf ( n18556 , n18552 );
and ( n18557 , n18555 , n18556 );
nor ( n18558 , n18554 , n18557 );
xor ( n18559 , n18549 , n18558 );
not ( n18560 , n18559 );
not ( n18561 , n18560 );
buf ( n18562 , n5994 );
not ( n18563 , n18562 );
not ( n18564 , n8233 );
not ( n18565 , n18564 );
or ( n18566 , n18563 , n18565 );
not ( n18567 , n8233 );
or ( n18568 , n18567 , n18562 );
nand ( n18569 , n18566 , n18568 );
not ( n18570 , n18569 );
or ( n18571 , n18561 , n18570 );
buf ( n18572 , n18559 );
not ( n18573 , n18572 );
or ( n18574 , n18569 , n18573 );
nand ( n18575 , n18571 , n18574 );
not ( n18576 , n18575 );
nand ( n18577 , n18530 , n18576 );
not ( n18578 , n18577 );
not ( n18579 , n13935 );
not ( n18580 , n9476 );
not ( n18581 , n13984 );
or ( n18582 , n18580 , n18581 );
not ( n18583 , n9476 );
nand ( n18584 , n18583 , n13991 );
nand ( n18585 , n18582 , n18584 );
xor ( n18586 , n18579 , n18585 );
buf ( n18587 , n18586 );
not ( n18588 , n18587 );
and ( n18589 , n18578 , n18588 );
and ( n18590 , n18577 , n18587 );
nor ( n18591 , n18589 , n18590 );
not ( n18592 , n18591 );
not ( n18593 , n18592 );
or ( n18594 , n18483 , n18593 );
nand ( n18595 , n18591 , n18481 );
nand ( n18596 , n18594 , n18595 );
not ( n18597 , n18596 );
buf ( n18598 , n5995 );
buf ( n18599 , n18598 );
not ( n18600 , n18599 );
not ( n18601 , n11501 );
or ( n18602 , n18600 , n18601 );
or ( n18603 , n11501 , n18599 );
nand ( n18604 , n18602 , n18603 );
and ( n18605 , n18604 , n15361 );
not ( n18606 , n18604 );
not ( n18607 , n15340 );
not ( n18608 , n15356 );
or ( n18609 , n18607 , n18608 );
or ( n18610 , n15356 , n15340 );
nand ( n18611 , n18609 , n18610 );
not ( n18612 , n18611 );
and ( n18613 , n18606 , n18612 );
or ( n18614 , n18605 , n18613 );
not ( n18615 , n9374 );
buf ( n18616 , n12830 );
xor ( n18617 , n18616 , n12827 );
not ( n18618 , n18617 );
not ( n18619 , n9321 );
or ( n18620 , n18618 , n18619 );
or ( n18621 , n9321 , n18617 );
nand ( n18622 , n18620 , n18621 );
not ( n18623 , n18622 );
or ( n18624 , n18615 , n18623 );
or ( n18625 , n18622 , n9374 );
nand ( n18626 , n18624 , n18625 );
nand ( n18627 , n18614 , n18626 );
not ( n18628 , n11310 );
not ( n18629 , n17672 );
or ( n18630 , n18628 , n18629 );
not ( n18631 , n17672 );
not ( n18632 , n18631 );
or ( n18633 , n18632 , n11310 );
nand ( n18634 , n18630 , n18633 );
not ( n18635 , n18634 );
not ( n18636 , n17333 );
and ( n18637 , n18635 , n18636 );
and ( n18638 , n18634 , n17333 );
nor ( n18639 , n18637 , n18638 );
and ( n18640 , n18627 , n18639 );
not ( n18641 , n18627 );
not ( n18642 , n18639 );
and ( n18643 , n18641 , n18642 );
nor ( n18644 , n18640 , n18643 );
not ( n18645 , n18644 );
buf ( n18646 , n6767 );
not ( n18647 , n18646 );
not ( n18648 , n12594 );
or ( n18649 , n18647 , n18648 );
not ( n18650 , n12591 );
or ( n18651 , n18650 , n18646 );
nand ( n18652 , n18649 , n18651 );
and ( n18653 , n18652 , n12636 );
not ( n18654 , n18652 );
not ( n18655 , n12636 );
and ( n18656 , n18654 , n18655 );
nor ( n18657 , n18653 , n18656 );
buf ( n18658 , n11003 );
not ( n18659 , n18658 );
not ( n18660 , n9694 );
or ( n18661 , n18659 , n18660 );
or ( n18662 , n9694 , n18658 );
nand ( n18663 , n18661 , n18662 );
buf ( n18664 , n6475 );
xor ( n18665 , n18664 , n9712 );
not ( n18666 , n9729 );
xnor ( n18667 , n18665 , n18666 );
buf ( n18668 , n18667 );
and ( n18669 , n18663 , n18668 );
not ( n18670 , n18663 );
and ( n18671 , n18670 , n9731 );
nor ( n18672 , n18669 , n18671 );
nand ( n18673 , n18657 , n18672 );
not ( n18674 , n18673 );
not ( n18675 , n10787 );
buf ( n18676 , n5996 );
buf ( n18677 , n18676 );
not ( n18678 , n18677 );
buf ( n18679 , n5997 );
not ( n18680 , n18679 );
not ( n18681 , n18680 );
or ( n18682 , n18678 , n18681 );
not ( n18683 , n18676 );
buf ( n18684 , n18679 );
nand ( n18685 , n18683 , n18684 );
nand ( n18686 , n18682 , n18685 );
buf ( n18687 , n5998 );
buf ( n18688 , n18687 );
and ( n18689 , n18686 , n18688 );
not ( n18690 , n18686 );
not ( n18691 , n18687 );
and ( n18692 , n18690 , n18691 );
nor ( n18693 , n18689 , n18692 );
buf ( n18694 , n5999 );
nand ( n18695 , n7355 , n18694 );
buf ( n18696 , n6000 );
buf ( n18697 , n18696 );
and ( n18698 , n18695 , n18697 );
not ( n18699 , n18695 );
not ( n18700 , n18696 );
and ( n18701 , n18699 , n18700 );
nor ( n18702 , n18698 , n18701 );
not ( n18703 , n18702 );
xor ( n18704 , n18693 , n18703 );
xnor ( n18705 , n18704 , n17705 );
not ( n18706 , n18705 );
or ( n18707 , n18675 , n18706 );
not ( n18708 , n10787 );
xor ( n18709 , n18693 , n18702 );
xnor ( n18710 , n18709 , n17705 );
nand ( n18711 , n18708 , n18710 );
nand ( n18712 , n18707 , n18711 );
not ( n18713 , n13294 );
not ( n18714 , n18713 );
and ( n18715 , n18712 , n18714 );
not ( n18716 , n18712 );
and ( n18717 , n18716 , n12342 );
nor ( n18718 , n18715 , n18717 );
not ( n18719 , n18718 );
not ( n18720 , n18719 );
not ( n18721 , n18720 );
and ( n18722 , n18674 , n18721 );
and ( n18723 , n18673 , n18720 );
nor ( n18724 , n18722 , n18723 );
not ( n18725 , n18724 );
and ( n18726 , n18645 , n18725 );
and ( n18727 , n18644 , n18724 );
nor ( n18728 , n18726 , n18727 );
xor ( n18729 , n8595 , n7025 );
buf ( n18730 , n6982 );
xnor ( n18731 , n18729 , n18730 );
not ( n18732 , n18731 );
not ( n18733 , n12713 );
buf ( n18734 , n18508 );
not ( n18735 , n18734 );
and ( n18736 , n18733 , n18735 );
and ( n18737 , n12713 , n18734 );
nor ( n18738 , n18736 , n18737 );
and ( n18739 , n18738 , n12755 );
not ( n18740 , n18738 );
and ( n18741 , n18740 , n17893 );
nor ( n18742 , n18739 , n18741 );
nand ( n18743 , n18732 , n18742 );
not ( n18744 , n7818 );
not ( n18745 , n17590 );
or ( n18746 , n18744 , n18745 );
nand ( n18747 , n17603 , n7814 );
nand ( n18748 , n18746 , n18747 );
and ( n18749 , n18748 , n10695 );
not ( n18750 , n18748 );
not ( n18751 , n10695 );
and ( n18752 , n18750 , n18751 );
nor ( n18753 , n18749 , n18752 );
buf ( n18754 , n18753 );
not ( n18755 , n18754 );
and ( n18756 , n18743 , n18755 );
not ( n18757 , n18743 );
and ( n18758 , n18757 , n18754 );
nor ( n18759 , n18756 , n18758 );
not ( n18760 , n18759 );
and ( n18761 , n18728 , n18760 );
not ( n18762 , n18728 );
and ( n18763 , n18762 , n18759 );
nor ( n18764 , n18761 , n18763 );
not ( n18765 , n18764 );
not ( n18766 , n18765 );
or ( n18767 , n18597 , n18766 );
not ( n18768 , n18596 );
nand ( n18769 , n18764 , n18768 );
nand ( n18770 , n18767 , n18769 );
buf ( n18771 , n18770 );
not ( n18772 , n18771 );
and ( n18773 , n18435 , n18772 );
not ( n18774 , n18435 );
and ( n18775 , n18774 , n18771 );
nor ( n18776 , n18773 , n18775 );
not ( n18777 , n18776 );
buf ( n18778 , n6001 );
nand ( n18779 , n11847 , n18778 );
buf ( n18780 , n6002 );
not ( n18781 , n18780 );
and ( n18782 , n18779 , n18781 );
not ( n18783 , n18779 );
buf ( n18784 , n18780 );
and ( n18785 , n18783 , n18784 );
nor ( n18786 , n18782 , n18785 );
xor ( n18787 , n18786 , n16149 );
xnor ( n18788 , n18787 , n11775 );
not ( n18789 , n18788 );
not ( n18790 , n18789 );
buf ( n18791 , n6003 );
buf ( n18792 , n18791 );
not ( n18793 , n18792 );
not ( n18794 , n7086 );
not ( n18795 , n18794 );
or ( n18796 , n18793 , n18795 );
not ( n18797 , n18791 );
nand ( n18798 , n18797 , n7087 );
nand ( n18799 , n18796 , n18798 );
buf ( n18800 , n6004 );
buf ( n18801 , n18800 );
and ( n18802 , n18799 , n18801 );
not ( n18803 , n18799 );
not ( n18804 , n18800 );
and ( n18805 , n18803 , n18804 );
nor ( n18806 , n18802 , n18805 );
buf ( n18807 , n6005 );
nand ( n18808 , n6927 , n18807 );
buf ( n18809 , n6006 );
xor ( n18810 , n18808 , n18809 );
xor ( n18811 , n18806 , n18810 );
buf ( n18812 , n6007 );
nand ( n18813 , n8260 , n18812 );
buf ( n18814 , n6008 );
buf ( n18815 , n18814 );
and ( n18816 , n18813 , n18815 );
not ( n18817 , n18813 );
not ( n18818 , n18814 );
and ( n18819 , n18817 , n18818 );
nor ( n18820 , n18816 , n18819 );
xnor ( n18821 , n18811 , n18820 );
buf ( n18822 , n18821 );
buf ( n18823 , n18822 );
not ( n18824 , n18823 );
buf ( n18825 , n6009 );
buf ( n18826 , n18825 );
not ( n18827 , n18826 );
buf ( n18828 , n6010 );
not ( n18829 , n18828 );
not ( n18830 , n18829 );
or ( n18831 , n18827 , n18830 );
not ( n18832 , n18825 );
buf ( n18833 , n18828 );
nand ( n18834 , n18832 , n18833 );
nand ( n18835 , n18831 , n18834 );
buf ( n18836 , n6011 );
buf ( n18837 , n18836 );
and ( n18838 , n18835 , n18837 );
not ( n18839 , n18835 );
not ( n18840 , n18836 );
and ( n18841 , n18839 , n18840 );
nor ( n18842 , n18838 , n18841 );
buf ( n18843 , n6012 );
nand ( n18844 , n6577 , n18843 );
buf ( n18845 , n6013 );
not ( n18846 , n18845 );
and ( n18847 , n18844 , n18846 );
not ( n18848 , n18844 );
buf ( n18849 , n18845 );
and ( n18850 , n18848 , n18849 );
nor ( n18851 , n18847 , n18850 );
xor ( n18852 , n18842 , n18851 );
buf ( n18853 , n6014 );
nand ( n18854 , n6515 , n18853 );
buf ( n18855 , n6015 );
not ( n18856 , n18855 );
and ( n18857 , n18854 , n18856 );
not ( n18858 , n18854 );
buf ( n18859 , n18855 );
and ( n18860 , n18858 , n18859 );
nor ( n18861 , n18857 , n18860 );
xor ( n18862 , n18852 , n18861 );
buf ( n18863 , n18862 );
xor ( n18864 , n7159 , n18863 );
not ( n18865 , n18864 );
or ( n18866 , n18824 , n18865 );
or ( n18867 , n18864 , n18823 );
nand ( n18868 , n18866 , n18867 );
buf ( n18869 , n6016 );
buf ( n18870 , n18869 );
not ( n18871 , n18870 );
not ( n18872 , n18461 );
or ( n18873 , n18871 , n18872 );
not ( n18874 , n18869 );
nand ( n18875 , n18462 , n18874 );
nand ( n18876 , n18873 , n18875 );
not ( n18877 , n18876 );
not ( n18878 , n18465 );
and ( n18879 , n18877 , n18878 );
and ( n18880 , n18876 , n18465 );
nor ( n18881 , n18879 , n18880 );
nor ( n18882 , n18868 , n18881 );
not ( n18883 , n18882 );
and ( n18884 , n18790 , n18883 );
and ( n18885 , n18789 , n18882 );
nor ( n18886 , n18884 , n18885 );
not ( n18887 , n18886 );
not ( n18888 , n18887 );
not ( n18889 , n7370 );
not ( n18890 , n18889 );
xor ( n18891 , n9460 , n18890 );
xnor ( n18892 , n18891 , n8843 );
not ( n18893 , n17560 );
not ( n18894 , n8888 );
or ( n18895 , n18893 , n18894 );
not ( n18896 , n17560 );
not ( n18897 , n8888 );
nand ( n18898 , n18896 , n18897 );
nand ( n18899 , n18895 , n18898 );
not ( n18900 , n18899 );
not ( n18901 , n8916 );
and ( n18902 , n18900 , n18901 );
and ( n18903 , n18899 , n8916 );
nor ( n18904 , n18902 , n18903 );
not ( n18905 , n18904 );
nand ( n18906 , n18892 , n18905 );
buf ( n18907 , n6017 );
nand ( n18908 , n6871 , n18907 );
buf ( n18909 , n6018 );
xor ( n18910 , n18908 , n18909 );
buf ( n18911 , n18910 );
not ( n18912 , n18911 );
not ( n18913 , n18912 );
not ( n18914 , n10581 );
or ( n18915 , n18913 , n18914 );
nand ( n18916 , n10587 , n18911 );
nand ( n18917 , n18915 , n18916 );
buf ( n18918 , n6019 );
buf ( n18919 , n18918 );
not ( n18920 , n18919 );
buf ( n18921 , n6020 );
not ( n18922 , n18921 );
not ( n18923 , n18922 );
or ( n18924 , n18920 , n18923 );
not ( n18925 , n18918 );
buf ( n18926 , n18921 );
nand ( n18927 , n18925 , n18926 );
nand ( n18928 , n18924 , n18927 );
buf ( n18929 , n6021 );
buf ( n18930 , n18929 );
and ( n18931 , n18928 , n18930 );
not ( n18932 , n18928 );
not ( n18933 , n18929 );
and ( n18934 , n18932 , n18933 );
nor ( n18935 , n18931 , n18934 );
buf ( n18936 , n6022 );
nand ( n18937 , n6646 , n18936 );
buf ( n18938 , n6023 );
buf ( n18939 , n18938 );
and ( n18940 , n18937 , n18939 );
not ( n18941 , n18937 );
not ( n18942 , n18938 );
and ( n18943 , n18941 , n18942 );
nor ( n18944 , n18940 , n18943 );
xor ( n18945 , n18935 , n18944 );
buf ( n18946 , n6024 );
nand ( n18947 , n10372 , n18946 );
buf ( n18948 , n6025 );
not ( n18949 , n18948 );
and ( n18950 , n18947 , n18949 );
not ( n18951 , n18947 );
buf ( n18952 , n18948 );
and ( n18953 , n18951 , n18952 );
nor ( n18954 , n18950 , n18953 );
xor ( n18955 , n18945 , n18954 );
buf ( n18956 , n18955 );
not ( n18957 , n18956 );
and ( n18958 , n18917 , n18957 );
not ( n18959 , n18917 );
and ( n18960 , n18959 , n18956 );
nor ( n18961 , n18958 , n18960 );
not ( n18962 , n18961 );
and ( n18963 , n18906 , n18962 );
not ( n18964 , n18906 );
and ( n18965 , n18964 , n18961 );
nor ( n18966 , n18963 , n18965 );
not ( n18967 , n18966 );
not ( n18968 , n18967 );
nand ( n18969 , n18789 , n18868 );
not ( n18970 , n18969 );
buf ( n18971 , n6026 );
nand ( n18972 , n8781 , n18971 );
not ( n18973 , n18972 );
buf ( n18974 , n6027 );
not ( n18975 , n18974 );
and ( n18976 , n18973 , n18975 );
and ( n18977 , n18972 , n18974 );
nor ( n18978 , n18976 , n18977 );
xor ( n18979 , n18978 , n17614 );
xnor ( n18980 , n18979 , n13547 );
not ( n18981 , n18980 );
not ( n18982 , n18981 );
and ( n18983 , n18970 , n18982 );
and ( n18984 , n18969 , n18981 );
nor ( n18985 , n18983 , n18984 );
not ( n18986 , n18985 );
not ( n18987 , n18986 );
or ( n18988 , n18968 , n18987 );
nand ( n18989 , n18985 , n18966 );
nand ( n18990 , n18988 , n18989 );
not ( n18991 , n18990 );
buf ( n18992 , n6028 );
nand ( n18993 , n6605 , n18992 );
buf ( n18994 , n6029 );
not ( n18995 , n18994 );
and ( n18996 , n18993 , n18995 );
not ( n18997 , n18993 );
buf ( n18998 , n18994 );
and ( n18999 , n18997 , n18998 );
nor ( n19000 , n18996 , n18999 );
not ( n19001 , n19000 );
not ( n19002 , n19001 );
not ( n19003 , n19002 );
buf ( n19004 , n12348 );
xor ( n19005 , n19004 , n12358 );
xnor ( n19006 , n19005 , n12374 );
not ( n19007 , n19006 );
not ( n19008 , n19007 );
or ( n19009 , n19003 , n19008 );
not ( n19010 , n19002 );
nand ( n19011 , n19010 , n19006 );
nand ( n19012 , n19009 , n19011 );
buf ( n19013 , n6030 );
buf ( n19014 , n19013 );
not ( n19015 , n19014 );
buf ( n19016 , n6031 );
not ( n19017 , n19016 );
not ( n19018 , n19017 );
or ( n19019 , n19015 , n19018 );
not ( n19020 , n19013 );
buf ( n19021 , n19016 );
nand ( n19022 , n19020 , n19021 );
nand ( n19023 , n19019 , n19022 );
buf ( n19024 , n6032 );
buf ( n19025 , n19024 );
and ( n19026 , n19023 , n19025 );
not ( n19027 , n19023 );
not ( n19028 , n19024 );
and ( n19029 , n19027 , n19028 );
nor ( n19030 , n19026 , n19029 );
xor ( n19031 , n19030 , n18910 );
buf ( n19032 , n6033 );
nand ( n19033 , n7569 , n19032 );
buf ( n19034 , n6034 );
not ( n19035 , n19034 );
and ( n19036 , n19033 , n19035 );
not ( n19037 , n19033 );
buf ( n19038 , n19034 );
and ( n19039 , n19037 , n19038 );
nor ( n19040 , n19036 , n19039 );
xor ( n19041 , n19031 , n19040 );
not ( n19042 , n19041 );
and ( n19043 , n19012 , n19042 );
not ( n19044 , n19012 );
buf ( n19045 , n19041 );
and ( n19046 , n19044 , n19045 );
nor ( n19047 , n19043 , n19046 );
not ( n19048 , n19047 );
not ( n19049 , n10306 );
not ( n19050 , n7848 );
and ( n19051 , n19049 , n19050 );
and ( n19052 , n10306 , n7848 );
nor ( n19053 , n19051 , n19052 );
not ( n19054 , n19053 );
not ( n19055 , n10296 );
or ( n19056 , n19054 , n19055 );
or ( n19057 , n10296 , n19053 );
nand ( n19058 , n19056 , n19057 );
and ( n19059 , n19058 , n9322 );
not ( n19060 , n19058 );
buf ( n19061 , n9321 );
and ( n19062 , n19060 , n19061 );
nor ( n19063 , n19059 , n19062 );
not ( n19064 , n19063 );
not ( n19065 , n12205 );
buf ( n19066 , n6035 );
buf ( n19067 , n19066 );
not ( n19068 , n19067 );
buf ( n19069 , n6036 );
not ( n19070 , n19069 );
not ( n19071 , n19070 );
or ( n19072 , n19068 , n19071 );
not ( n19073 , n19066 );
buf ( n19074 , n19069 );
nand ( n19075 , n19073 , n19074 );
nand ( n19076 , n19072 , n19075 );
and ( n19077 , n19076 , n17686 );
not ( n19078 , n19076 );
not ( n19079 , n17685 );
and ( n19080 , n19078 , n19079 );
nor ( n19081 , n19077 , n19080 );
buf ( n19082 , n6037 );
nand ( n19083 , n6719 , n19082 );
buf ( n19084 , n6038 );
buf ( n19085 , n19084 );
and ( n19086 , n19083 , n19085 );
not ( n19087 , n19083 );
not ( n19088 , n19084 );
and ( n19089 , n19087 , n19088 );
nor ( n19090 , n19086 , n19089 );
not ( n19091 , n19090 );
xor ( n19092 , n19081 , n19091 );
xnor ( n19093 , n19092 , n12771 );
not ( n19094 , n19093 );
or ( n19095 , n19065 , n19094 );
not ( n19096 , n12205 );
xor ( n19097 , n19081 , n19090 );
xnor ( n19098 , n19097 , n12771 );
nand ( n19099 , n19096 , n19098 );
nand ( n19100 , n19095 , n19099 );
buf ( n19101 , n9694 );
not ( n19102 , n19101 );
and ( n19103 , n19100 , n19102 );
not ( n19104 , n19100 );
not ( n19105 , n9695 );
and ( n19106 , n19104 , n19105 );
nor ( n19107 , n19103 , n19106 );
nand ( n19108 , n19064 , n19107 );
not ( n19109 , n19108 );
and ( n19110 , n19048 , n19109 );
and ( n19111 , n19108 , n19047 );
nor ( n19112 , n19110 , n19111 );
not ( n19113 , n19112 );
not ( n19114 , n19113 );
buf ( n19115 , n6039 );
buf ( n19116 , n19115 );
not ( n19117 , n19116 );
buf ( n19118 , n6040 );
buf ( n19119 , n19118 );
not ( n19120 , n19119 );
buf ( n19121 , n6041 );
not ( n19122 , n19121 );
not ( n19123 , n19122 );
or ( n19124 , n19120 , n19123 );
not ( n19125 , n19118 );
buf ( n19126 , n19121 );
nand ( n19127 , n19125 , n19126 );
nand ( n19128 , n19124 , n19127 );
not ( n19129 , n19128 );
not ( n19130 , n19129 );
or ( n19131 , n19117 , n19130 );
not ( n19132 , n19115 );
nand ( n19133 , n19128 , n19132 );
nand ( n19134 , n19131 , n19133 );
not ( n19135 , n19134 );
buf ( n19136 , n6042 );
buf ( n19137 , n6043 );
nand ( n19138 , n6815 , n19137 );
buf ( n19139 , n6044 );
buf ( n19140 , n19139 );
and ( n19141 , n19138 , n19140 );
not ( n19142 , n19138 );
not ( n19143 , n19139 );
and ( n19144 , n19142 , n19143 );
nor ( n19145 , n19141 , n19144 );
xor ( n19146 , n19136 , n19145 );
buf ( n19147 , n6045 );
nand ( n19148 , n7247 , n19147 );
buf ( n19149 , n6046 );
buf ( n19150 , n19149 );
and ( n19151 , n19148 , n19150 );
not ( n19152 , n19148 );
not ( n19153 , n19149 );
and ( n19154 , n19152 , n19153 );
nor ( n19155 , n19151 , n19154 );
xnor ( n19156 , n19146 , n19155 );
buf ( n19157 , n19156 );
not ( n19158 , n19157 );
or ( n19159 , n19135 , n19158 );
or ( n19160 , n19157 , n19134 );
nand ( n19161 , n19159 , n19160 );
buf ( n19162 , n6047 );
buf ( n19163 , n19162 );
not ( n19164 , n19163 );
buf ( n19165 , n6048 );
not ( n19166 , n19165 );
not ( n19167 , n19166 );
or ( n19168 , n19164 , n19167 );
not ( n19169 , n19162 );
buf ( n19170 , n19165 );
nand ( n19171 , n19169 , n19170 );
nand ( n19172 , n19168 , n19171 );
buf ( n19173 , n6049 );
not ( n19174 , n19173 );
and ( n19175 , n19172 , n19174 );
not ( n19176 , n19172 );
buf ( n19177 , n19173 );
and ( n19178 , n19176 , n19177 );
nor ( n19179 , n19175 , n19178 );
buf ( n19180 , n6050 );
nand ( n19181 , n9812 , n19180 );
buf ( n19182 , n6051 );
buf ( n19183 , n19182 );
and ( n19184 , n19181 , n19183 );
not ( n19185 , n19181 );
not ( n19186 , n19182 );
and ( n19187 , n19185 , n19186 );
nor ( n19188 , n19184 , n19187 );
xor ( n19189 , n19179 , n19188 );
buf ( n19190 , n6052 );
nand ( n19191 , n8675 , n19190 );
buf ( n19192 , n6053 );
not ( n19193 , n19192 );
and ( n19194 , n19191 , n19193 );
not ( n19195 , n19191 );
buf ( n19196 , n19192 );
and ( n19197 , n19195 , n19196 );
nor ( n19198 , n19194 , n19197 );
xnor ( n19199 , n19189 , n19198 );
buf ( n19200 , n19199 );
and ( n19201 , n19161 , n19200 );
not ( n19202 , n19161 );
xor ( n19203 , n19179 , n19188 );
xor ( n19204 , n19203 , n19198 );
and ( n19205 , n19202 , n19204 );
nor ( n19206 , n19201 , n19205 );
buf ( n19207 , n6054 );
buf ( n19208 , n19207 );
not ( n19209 , n19208 );
buf ( n19210 , n6055 );
not ( n19211 , n19210 );
buf ( n19212 , n6056 );
buf ( n19213 , n19212 );
and ( n19214 , n19211 , n19213 );
not ( n19215 , n19211 );
not ( n19216 , n19212 );
and ( n19217 , n19215 , n19216 );
nor ( n19218 , n19214 , n19217 );
not ( n19219 , n19218 );
or ( n19220 , n19209 , n19219 );
or ( n19221 , n19218 , n19208 );
nand ( n19222 , n19220 , n19221 );
not ( n19223 , n19222 );
buf ( n19224 , n6057 );
not ( n19225 , n19224 );
xor ( n19226 , n13789 , n19225 );
buf ( n19227 , n6058 );
nand ( n19228 , n6916 , n19227 );
buf ( n19229 , n6059 );
not ( n19230 , n19229 );
and ( n19231 , n19228 , n19230 );
not ( n19232 , n19228 );
buf ( n19233 , n19229 );
and ( n19234 , n19232 , n19233 );
nor ( n19235 , n19231 , n19234 );
xnor ( n19236 , n19226 , n19235 );
not ( n19237 , n19236 );
not ( n19238 , n19237 );
or ( n19239 , n19223 , n19238 );
or ( n19240 , n19237 , n19222 );
nand ( n19241 , n19239 , n19240 );
not ( n19242 , n19241 );
buf ( n19243 , n11226 );
not ( n19244 , n19243 );
and ( n19245 , n19242 , n19244 );
and ( n19246 , n19241 , n11228 );
nor ( n19247 , n19245 , n19246 );
not ( n19248 , n19247 );
nand ( n19249 , n19206 , n19248 );
not ( n19250 , n19249 );
buf ( n19251 , n13161 );
xor ( n19252 , n19251 , n13642 );
buf ( n19253 , n6060 );
buf ( n19254 , n6061 );
buf ( n19255 , n19254 );
not ( n19256 , n19255 );
buf ( n19257 , n6062 );
not ( n19258 , n19257 );
not ( n19259 , n19258 );
or ( n19260 , n19256 , n19259 );
not ( n19261 , n19254 );
buf ( n19262 , n19257 );
nand ( n19263 , n19261 , n19262 );
nand ( n19264 , n19260 , n19263 );
xor ( n19265 , n19253 , n19264 );
buf ( n19266 , n6063 );
buf ( n19267 , n6064 );
not ( n19268 , n19267 );
xor ( n19269 , n19266 , n19268 );
buf ( n19270 , n6065 );
nand ( n19271 , n8032 , n19270 );
xnor ( n19272 , n19269 , n19271 );
xnor ( n19273 , n19265 , n19272 );
buf ( n19274 , n19273 );
and ( n19275 , n19252 , n19274 );
not ( n19276 , n19252 );
not ( n19277 , n19274 );
and ( n19278 , n19276 , n19277 );
nor ( n19279 , n19275 , n19278 );
not ( n19280 , n19279 );
or ( n19281 , n19250 , n19280 );
or ( n19282 , n19279 , n19249 );
nand ( n19283 , n19281 , n19282 );
not ( n19284 , n19283 );
not ( n19285 , n19284 );
or ( n19286 , n19114 , n19285 );
nand ( n19287 , n19283 , n19112 );
nand ( n19288 , n19286 , n19287 );
not ( n19289 , n13925 );
buf ( n19290 , n16838 );
not ( n19291 , n19290 );
or ( n19292 , n19289 , n19291 );
buf ( n19293 , n17263 );
nand ( n19294 , n19293 , n13921 );
nand ( n19295 , n19292 , n19294 );
not ( n19296 , n19295 );
not ( n19297 , n16881 );
buf ( n19298 , n19297 );
not ( n19299 , n19298 );
and ( n19300 , n19296 , n19299 );
and ( n19301 , n19295 , n19298 );
nor ( n19302 , n19300 , n19301 );
not ( n19303 , n19302 );
buf ( n19304 , n6066 );
not ( n19305 , n15251 );
buf ( n19306 , n6067 );
not ( n19307 , n19306 );
not ( n19308 , n19307 );
or ( n19309 , n19305 , n19308 );
not ( n19310 , n15250 );
buf ( n19311 , n19306 );
nand ( n19312 , n19310 , n19311 );
nand ( n19313 , n19309 , n19312 );
xor ( n19314 , n19304 , n19313 );
buf ( n19315 , n6068 );
buf ( n19316 , n6069 );
not ( n19317 , n19316 );
xor ( n19318 , n19315 , n19317 );
buf ( n19319 , n6070 );
nand ( n19320 , n7912 , n19319 );
xnor ( n19321 , n19318 , n19320 );
xnor ( n19322 , n19314 , n19321 );
buf ( n19323 , n19322 );
not ( n19324 , n19323 );
not ( n19325 , n19324 );
not ( n19326 , n17903 );
buf ( n19327 , n6071 );
buf ( n19328 , n19327 );
not ( n19329 , n19328 );
buf ( n19330 , n6072 );
not ( n19331 , n19330 );
not ( n19332 , n19331 );
or ( n19333 , n19329 , n19332 );
not ( n19334 , n19327 );
buf ( n19335 , n19330 );
nand ( n19336 , n19334 , n19335 );
nand ( n19337 , n19333 , n19336 );
buf ( n19338 , n6073 );
not ( n19339 , n19338 );
and ( n19340 , n19337 , n19339 );
not ( n19341 , n19337 );
buf ( n19342 , n19338 );
and ( n19343 , n19341 , n19342 );
nor ( n19344 , n19340 , n19343 );
buf ( n19345 , n6074 );
nand ( n19346 , n7698 , n19345 );
buf ( n19347 , n6075 );
not ( n19348 , n19347 );
and ( n19349 , n19346 , n19348 );
not ( n19350 , n19346 );
buf ( n19351 , n19347 );
and ( n19352 , n19350 , n19351 );
nor ( n19353 , n19349 , n19352 );
xor ( n19354 , n19344 , n19353 );
buf ( n19355 , n6076 );
nand ( n19356 , n11946 , n19355 );
buf ( n19357 , n6077 );
not ( n19358 , n19357 );
and ( n19359 , n19356 , n19358 );
not ( n19360 , n19356 );
buf ( n19361 , n19357 );
and ( n19362 , n19360 , n19361 );
nor ( n19363 , n19359 , n19362 );
xnor ( n19364 , n19354 , n19363 );
buf ( n19365 , n19364 );
not ( n19366 , n19365 );
not ( n19367 , n19366 );
or ( n19368 , n19326 , n19367 );
not ( n19369 , n17903 );
not ( n19370 , n19364 );
not ( n19371 , n19370 );
nand ( n19372 , n19369 , n19371 );
nand ( n19373 , n19368 , n19372 );
not ( n19374 , n19373 );
or ( n19375 , n19325 , n19374 );
or ( n19376 , n19324 , n19373 );
nand ( n19377 , n19375 , n19376 );
not ( n19378 , n19377 );
nand ( n19379 , n19303 , n19378 );
not ( n19380 , n19379 );
not ( n19381 , n12009 );
not ( n19382 , n16910 );
or ( n19383 , n19381 , n19382 );
not ( n19384 , n12009 );
nand ( n19385 , n19384 , n10824 );
nand ( n19386 , n19383 , n19385 );
xor ( n19387 , n19386 , n16917 );
not ( n19388 , n19387 );
not ( n19389 , n19388 );
and ( n19390 , n19380 , n19389 );
and ( n19391 , n19379 , n19388 );
nor ( n19392 , n19390 , n19391 );
and ( n19393 , n19288 , n19392 );
not ( n19394 , n19288 );
not ( n19395 , n19392 );
and ( n19396 , n19394 , n19395 );
nor ( n19397 , n19393 , n19396 );
not ( n19398 , n19397 );
and ( n19399 , n18991 , n19398 );
and ( n19400 , n18990 , n19397 );
nor ( n19401 , n19399 , n19400 );
not ( n19402 , n19401 );
or ( n19403 , n18888 , n19402 );
not ( n19404 , n18887 );
not ( n19405 , n19397 );
and ( n19406 , n18990 , n19405 );
not ( n19407 , n18990 );
and ( n19408 , n19407 , n19397 );
nor ( n19409 , n19406 , n19408 );
nand ( n19410 , n19404 , n19409 );
nand ( n19411 , n19403 , n19410 );
xor ( n19412 , n16043 , n14152 );
xnor ( n19413 , n19412 , n14175 );
not ( n19414 , n19413 );
not ( n19415 , n7217 );
buf ( n19416 , n6078 );
buf ( n19417 , n19416 );
not ( n19418 , n19417 );
buf ( n19419 , n6079 );
not ( n19420 , n19419 );
not ( n19421 , n19420 );
or ( n19422 , n19418 , n19421 );
not ( n19423 , n19416 );
buf ( n19424 , n19419 );
nand ( n19425 , n19423 , n19424 );
nand ( n19426 , n19422 , n19425 );
and ( n19427 , n19426 , n18599 );
not ( n19428 , n19426 );
not ( n19429 , n18598 );
and ( n19430 , n19428 , n19429 );
nor ( n19431 , n19427 , n19430 );
xor ( n19432 , n19431 , n15372 );
buf ( n19433 , n6080 );
nand ( n19434 , n7107 , n19433 );
buf ( n19435 , n6081 );
buf ( n19436 , n19435 );
and ( n19437 , n19434 , n19436 );
not ( n19438 , n19434 );
not ( n19439 , n19435 );
and ( n19440 , n19438 , n19439 );
nor ( n19441 , n19437 , n19440 );
xnor ( n19442 , n19432 , n19441 );
buf ( n19443 , n19442 );
not ( n19444 , n19443 );
or ( n19445 , n19415 , n19444 );
not ( n19446 , n19442 );
buf ( n19447 , n19446 );
nand ( n19448 , n19447 , n7213 );
nand ( n19449 , n19445 , n19448 );
not ( n19450 , n18862 );
buf ( n19451 , n19450 );
xor ( n19452 , n19449 , n19451 );
nand ( n19453 , n19414 , n19452 );
buf ( n19454 , n6082 );
buf ( n19455 , n6083 );
buf ( n19456 , n19455 );
not ( n19457 , n19456 );
buf ( n19458 , n6084 );
not ( n19459 , n19458 );
not ( n19460 , n19459 );
or ( n19461 , n19457 , n19460 );
not ( n19462 , n19455 );
buf ( n19463 , n19458 );
nand ( n19464 , n19462 , n19463 );
nand ( n19465 , n19461 , n19464 );
not ( n19466 , n19465 );
xor ( n19467 , n19454 , n19466 );
xor ( n19468 , n11791 , n18974 );
xnor ( n19469 , n19468 , n18972 );
xnor ( n19470 , n19467 , n19469 );
not ( n19471 , n19470 );
xor ( n19472 , n16165 , n19471 );
xnor ( n19473 , n19472 , n10351 );
not ( n19474 , n19473 );
and ( n19475 , n19453 , n19474 );
not ( n19476 , n19453 );
and ( n19477 , n19476 , n19473 );
nor ( n19478 , n19475 , n19477 );
not ( n19479 , n19478 );
buf ( n19480 , n14373 );
not ( n19481 , n19480 );
not ( n19482 , n7097 );
buf ( n19483 , n6085 );
nand ( n19484 , n8323 , n19483 );
buf ( n19485 , n6086 );
buf ( n19486 , n19485 );
and ( n19487 , n19484 , n19486 );
not ( n19488 , n19484 );
not ( n19489 , n19485 );
and ( n19490 , n19488 , n19489 );
nor ( n19491 , n19487 , n19490 );
not ( n19492 , n19491 );
buf ( n19493 , n6087 );
nand ( n19494 , n6502 , n19493 );
buf ( n19495 , n6088 );
not ( n19496 , n19495 );
and ( n19497 , n19494 , n19496 );
not ( n19498 , n19494 );
buf ( n19499 , n19495 );
and ( n19500 , n19498 , n19499 );
nor ( n19501 , n19497 , n19500 );
not ( n19502 , n19501 );
or ( n19503 , n19492 , n19502 );
or ( n19504 , n19491 , n19501 );
nand ( n19505 , n19503 , n19504 );
buf ( n19506 , n6089 );
buf ( n19507 , n19506 );
not ( n19508 , n19507 );
not ( n19509 , n13011 );
or ( n19510 , n19508 , n19509 );
not ( n19511 , n19506 );
buf ( n19512 , n13010 );
nand ( n19513 , n19511 , n19512 );
nand ( n19514 , n19510 , n19513 );
buf ( n19515 , n6090 );
not ( n19516 , n19515 );
and ( n19517 , n19514 , n19516 );
not ( n19518 , n19514 );
buf ( n19519 , n19515 );
and ( n19520 , n19518 , n19519 );
nor ( n19521 , n19517 , n19520 );
and ( n19522 , n19505 , n19521 );
not ( n19523 , n19505 );
not ( n19524 , n19521 );
and ( n19525 , n19523 , n19524 );
nor ( n19526 , n19522 , n19525 );
buf ( n19527 , n19526 );
not ( n19528 , n19527 );
or ( n19529 , n19482 , n19528 );
or ( n19530 , n19527 , n7097 );
nand ( n19531 , n19529 , n19530 );
not ( n19532 , n19531 );
and ( n19533 , n19481 , n19532 );
and ( n19534 , n19480 , n19531 );
nor ( n19535 , n19533 , n19534 );
not ( n19536 , n19535 );
not ( n19537 , n19536 );
not ( n19538 , n10059 );
not ( n19539 , n15428 );
or ( n19540 , n19538 , n19539 );
not ( n19541 , n15424 );
nand ( n19542 , n19541 , n10055 );
nand ( n19543 , n19540 , n19542 );
and ( n19544 , n19543 , n15475 );
not ( n19545 , n19543 );
and ( n19546 , n19545 , n15471 );
or ( n19547 , n19544 , n19546 );
not ( n19548 , n19547 );
not ( n19549 , n7666 );
xor ( n19550 , n7605 , n7625 );
not ( n19551 , n7615 );
xnor ( n19552 , n19550 , n19551 );
buf ( n19553 , n6091 );
not ( n19554 , n19553 );
and ( n19555 , n19552 , n19554 );
not ( n19556 , n19552 );
buf ( n19557 , n19553 );
and ( n19558 , n19556 , n19557 );
nor ( n19559 , n19555 , n19558 );
not ( n19560 , n19559 );
and ( n19561 , n19549 , n19560 );
and ( n19562 , n7666 , n19559 );
nor ( n19563 , n19561 , n19562 );
not ( n19564 , n19563 );
nand ( n19565 , n19548 , n19564 );
not ( n19566 , n19565 );
or ( n19567 , n19537 , n19566 );
or ( n19568 , n19565 , n19536 );
nand ( n19569 , n19567 , n19568 );
not ( n19570 , n19569 );
and ( n19571 , n19479 , n19570 );
and ( n19572 , n19478 , n19569 );
nor ( n19573 , n19571 , n19572 );
not ( n19574 , n19573 );
not ( n19575 , n13758 );
buf ( n19576 , n6092 );
not ( n19577 , n19576 );
buf ( n19578 , n6093 );
not ( n19579 , n19578 );
buf ( n19580 , n6094 );
buf ( n19581 , n19580 );
nand ( n19582 , n19579 , n19581 );
not ( n19583 , n19580 );
buf ( n19584 , n19578 );
nand ( n19585 , n19583 , n19584 );
and ( n19586 , n19582 , n19585 );
xor ( n19587 , n19577 , n19586 );
buf ( n19588 , n6095 );
buf ( n19589 , n6096 );
xor ( n19590 , n19588 , n19589 );
buf ( n19591 , n6097 );
nand ( n19592 , n8608 , n19591 );
xnor ( n19593 , n19590 , n19592 );
xor ( n19594 , n19587 , n19593 );
not ( n19595 , n19594 );
not ( n19596 , n19595 );
or ( n19597 , n19575 , n19596 );
or ( n19598 , n19595 , n13758 );
nand ( n19599 , n19597 , n19598 );
not ( n19600 , n11910 );
not ( n19601 , n11914 );
and ( n19602 , n19600 , n19601 );
and ( n19603 , n11910 , n11914 );
nor ( n19604 , n19602 , n19603 );
buf ( n19605 , n19604 );
and ( n19606 , n19599 , n19605 );
not ( n19607 , n19599 );
buf ( n19608 , n11916 );
and ( n19609 , n19607 , n19608 );
nor ( n19610 , n19606 , n19609 );
not ( n19611 , n19610 );
not ( n19612 , n19611 );
not ( n19613 , n11054 );
not ( n19614 , n14717 );
and ( n19615 , n19613 , n19614 );
and ( n19616 , n11054 , n14717 );
nor ( n19617 , n19615 , n19616 );
not ( n19618 , n16756 );
buf ( n19619 , n19618 );
and ( n19620 , n19617 , n19619 );
not ( n19621 , n19617 );
not ( n19622 , n19618 );
and ( n19623 , n19621 , n19622 );
nor ( n19624 , n19620 , n19623 );
not ( n19625 , n19624 );
not ( n19626 , n11985 );
not ( n19627 , n16907 );
or ( n19628 , n19626 , n19627 );
not ( n19629 , n16906 );
or ( n19630 , n19629 , n11985 );
nand ( n19631 , n19628 , n19630 );
and ( n19632 , n19631 , n16914 );
not ( n19633 , n19631 );
and ( n19634 , n19633 , n14311 );
nor ( n19635 , n19632 , n19634 );
nand ( n19636 , n19625 , n19635 );
not ( n19637 , n19636 );
or ( n19638 , n19612 , n19637 );
buf ( n19639 , n19635 );
nand ( n19640 , n19625 , n19639 );
or ( n19641 , n19640 , n19611 );
nand ( n19642 , n19638 , n19641 );
not ( n19643 , n19642 );
buf ( n19644 , n6098 );
buf ( n19645 , n19644 );
not ( n19646 , n19645 );
buf ( n19647 , n6099 );
not ( n19648 , n19647 );
not ( n19649 , n19648 );
or ( n19650 , n19646 , n19649 );
not ( n19651 , n19644 );
buf ( n19652 , n19647 );
nand ( n19653 , n19651 , n19652 );
nand ( n19654 , n19650 , n19653 );
and ( n19655 , n19654 , n17134 );
not ( n19656 , n19654 );
not ( n19657 , n17133 );
and ( n19658 , n19656 , n19657 );
nor ( n19659 , n19655 , n19658 );
not ( n19660 , n19659 );
xor ( n19661 , n19660 , n9851 );
xnor ( n19662 , n19661 , n18398 );
and ( n19663 , n9143 , n19662 );
not ( n19664 , n9143 );
xor ( n19665 , n19659 , n9851 );
xnor ( n19666 , n19665 , n18398 );
and ( n19667 , n19664 , n19666 );
nor ( n19668 , n19663 , n19667 );
not ( n19669 , n19668 );
not ( n19670 , n19669 );
buf ( n19671 , n6100 );
not ( n19672 , n19671 );
buf ( n19673 , n6101 );
not ( n19674 , n19673 );
buf ( n19675 , n6102 );
buf ( n19676 , n19675 );
and ( n19677 , n19674 , n19676 );
not ( n19678 , n19674 );
not ( n19679 , n19675 );
and ( n19680 , n19678 , n19679 );
nor ( n19681 , n19677 , n19680 );
xor ( n19682 , n19672 , n19681 );
buf ( n19683 , n6103 );
buf ( n19684 , n6104 );
xor ( n19685 , n19683 , n19684 );
buf ( n19686 , n6105 );
nand ( n19687 , n6973 , n19686 );
xnor ( n19688 , n19685 , n19687 );
xnor ( n19689 , n19682 , n19688 );
not ( n19690 , n19689 );
or ( n19691 , n19670 , n19690 );
not ( n19692 , n19689 );
nand ( n19693 , n19692 , n19668 );
nand ( n19694 , n19691 , n19693 );
not ( n19695 , n19694 );
not ( n19696 , n12635 );
buf ( n19697 , n6106 );
not ( n19698 , n19697 );
and ( n19699 , n19696 , n19698 );
and ( n19700 , n12635 , n19697 );
nor ( n19701 , n19699 , n19700 );
buf ( n19702 , n6107 );
buf ( n19703 , n19702 );
not ( n19704 , n19703 );
buf ( n19705 , n6108 );
not ( n19706 , n19705 );
not ( n19707 , n19706 );
or ( n19708 , n19704 , n19707 );
not ( n19709 , n19702 );
buf ( n19710 , n19705 );
nand ( n19711 , n19709 , n19710 );
nand ( n19712 , n19708 , n19711 );
buf ( n19713 , n6109 );
not ( n19714 , n19713 );
and ( n19715 , n19712 , n19714 );
not ( n19716 , n19712 );
buf ( n19717 , n19713 );
and ( n19718 , n19716 , n19717 );
nor ( n19719 , n19715 , n19718 );
buf ( n19720 , n6110 );
nand ( n19721 , n7197 , n19720 );
buf ( n19722 , n6111 );
buf ( n19723 , n19722 );
and ( n19724 , n19721 , n19723 );
not ( n19725 , n19721 );
not ( n19726 , n19722 );
and ( n19727 , n19725 , n19726 );
nor ( n19728 , n19724 , n19727 );
xor ( n19729 , n19719 , n19728 );
buf ( n19730 , n6112 );
nand ( n19731 , n7067 , n19730 );
buf ( n19732 , n6113 );
not ( n19733 , n19732 );
and ( n19734 , n19731 , n19733 );
not ( n19735 , n19731 );
buf ( n19736 , n19732 );
and ( n19737 , n19735 , n19736 );
nor ( n19738 , n19734 , n19737 );
xnor ( n19739 , n19729 , n19738 );
not ( n19740 , n19739 );
not ( n19741 , n19740 );
and ( n19742 , n19701 , n19741 );
not ( n19743 , n19701 );
not ( n19744 , n19728 );
xor ( n19745 , n19719 , n19744 );
xnor ( n19746 , n19745 , n19738 );
buf ( n19747 , n19746 );
and ( n19748 , n19743 , n19747 );
nor ( n19749 , n19742 , n19748 );
nand ( n19750 , n19695 , n19749 );
not ( n19751 , n19750 );
not ( n19752 , n16621 );
not ( n19753 , n12206 );
or ( n19754 , n19752 , n19753 );
or ( n19755 , n12206 , n16621 );
nand ( n19756 , n19754 , n19755 );
not ( n19757 , n19756 );
not ( n19758 , n16250 );
and ( n19759 , n19757 , n19758 );
and ( n19760 , n19756 , n16250 );
nor ( n19761 , n19759 , n19760 );
not ( n19762 , n19761 );
not ( n19763 , n19762 );
and ( n19764 , n19751 , n19763 );
and ( n19765 , n19750 , n19762 );
nor ( n19766 , n19764 , n19765 );
not ( n19767 , n19766 );
or ( n19768 , n19643 , n19767 );
or ( n19769 , n19766 , n19642 );
nand ( n19770 , n19768 , n19769 );
not ( n19771 , n19770 );
not ( n19772 , n7891 );
not ( n19773 , n10270 );
not ( n19774 , n19773 );
not ( n19775 , n19774 );
or ( n19776 , n19772 , n19775 );
or ( n19777 , n10271 , n7891 );
nand ( n19778 , n19776 , n19777 );
and ( n19779 , n19778 , n10314 );
not ( n19780 , n19778 );
and ( n19781 , n19780 , n10311 );
nor ( n19782 , n19779 , n19781 );
not ( n19783 , n19782 );
buf ( n19784 , n15161 );
not ( n19785 , n19784 );
buf ( n19786 , n6114 );
buf ( n19787 , n19786 );
not ( n19788 , n19787 );
not ( n19789 , n19207 );
not ( n19790 , n19789 );
or ( n19791 , n19788 , n19790 );
not ( n19792 , n19786 );
nand ( n19793 , n19792 , n19208 );
nand ( n19794 , n19791 , n19793 );
buf ( n19795 , n6115 );
not ( n19796 , n19795 );
and ( n19797 , n19794 , n19796 );
not ( n19798 , n19794 );
buf ( n19799 , n19795 );
and ( n19800 , n19798 , n19799 );
nor ( n19801 , n19797 , n19800 );
buf ( n19802 , n6116 );
nand ( n19803 , n6770 , n19802 );
buf ( n19804 , n6117 );
not ( n19805 , n19804 );
and ( n19806 , n19803 , n19805 );
not ( n19807 , n19803 );
buf ( n19808 , n19804 );
and ( n19809 , n19807 , n19808 );
nor ( n19810 , n19806 , n19809 );
xor ( n19811 , n19801 , n19810 );
buf ( n19812 , n6118 );
nand ( n19813 , n7259 , n19812 );
buf ( n19814 , n6119 );
not ( n19815 , n19814 );
and ( n19816 , n19813 , n19815 );
not ( n19817 , n19813 );
buf ( n19818 , n19814 );
and ( n19819 , n19817 , n19818 );
nor ( n19820 , n19816 , n19819 );
xnor ( n19821 , n19811 , n19820 );
not ( n19822 , n19821 );
not ( n19823 , n19822 );
or ( n19824 , n19785 , n19823 );
not ( n19825 , n19784 );
not ( n19826 , n19822 );
nand ( n19827 , n19825 , n19826 );
nand ( n19828 , n19824 , n19827 );
buf ( n19829 , n13595 );
buf ( n19830 , n19829 );
and ( n19831 , n19828 , n19830 );
not ( n19832 , n19828 );
buf ( n19833 , n13591 );
buf ( n19834 , n19833 );
and ( n19835 , n19832 , n19834 );
nor ( n19836 , n19831 , n19835 );
nand ( n19837 , n19783 , n19836 );
not ( n19838 , n19837 );
not ( n19839 , n7580 );
nor ( n19840 , n7539 , n15863 );
not ( n19841 , n19840 );
nand ( n19842 , n7539 , n15863 );
nand ( n19843 , n19841 , n19842 );
not ( n19844 , n19843 );
or ( n19845 , n19839 , n19844 );
or ( n19846 , n19843 , n7580 );
nand ( n19847 , n19845 , n19846 );
not ( n19848 , n19847 );
and ( n19849 , n19838 , n19848 );
and ( n19850 , n19837 , n19847 );
nor ( n19851 , n19849 , n19850 );
not ( n19852 , n19851 );
or ( n19853 , n19771 , n19852 );
or ( n19854 , n19851 , n19770 );
nand ( n19855 , n19853 , n19854 );
not ( n19856 , n19855 );
or ( n19857 , n19574 , n19856 );
or ( n19858 , n19855 , n19573 );
nand ( n19859 , n19857 , n19858 );
buf ( n19860 , n19859 );
buf ( n19861 , n19860 );
not ( n19862 , n19861 );
and ( n19863 , n19411 , n19862 );
not ( n19864 , n19411 );
not ( n19865 , n19860 );
not ( n19866 , n19865 );
and ( n19867 , n19864 , n19866 );
nor ( n19868 , n19863 , n19867 );
nand ( n19869 , n18777 , n19868 );
buf ( n19870 , n10665 );
not ( n19871 , n19870 );
not ( n19872 , n13905 );
or ( n19873 , n19871 , n19872 );
buf ( n19874 , n13905 );
or ( n19875 , n19874 , n19870 );
nand ( n19876 , n19873 , n19875 );
not ( n19877 , n19876 );
not ( n19878 , n7803 );
or ( n19879 , n19877 , n19878 );
not ( n19880 , n7802 );
or ( n19881 , n19880 , n19876 );
nand ( n19882 , n19879 , n19881 );
not ( n19883 , n19882 );
not ( n19884 , n16716 );
not ( n19885 , n8354 );
buf ( n19886 , n16755 );
not ( n19887 , n19886 );
or ( n19888 , n19885 , n19887 );
or ( n19889 , n19886 , n8354 );
nand ( n19890 , n19888 , n19889 );
not ( n19891 , n19890 );
or ( n19892 , n19884 , n19891 );
or ( n19893 , n19890 , n16716 );
nand ( n19894 , n19892 , n19893 );
buf ( n19895 , n13627 );
not ( n19896 , n19895 );
not ( n19897 , n13722 );
buf ( n19898 , n6120 );
not ( n19899 , n19898 );
not ( n19900 , n19899 );
or ( n19901 , n19897 , n19900 );
not ( n19902 , n13721 );
buf ( n19903 , n19898 );
nand ( n19904 , n19902 , n19903 );
nand ( n19905 , n19901 , n19904 );
and ( n19906 , n19905 , n17615 );
not ( n19907 , n19905 );
and ( n19908 , n19907 , n17609 );
nor ( n19909 , n19906 , n19908 );
buf ( n19910 , n6121 );
nand ( n19911 , n7563 , n19910 );
buf ( n19912 , n6122 );
buf ( n19913 , n19912 );
and ( n19914 , n19911 , n19913 );
not ( n19915 , n19911 );
not ( n19916 , n19912 );
and ( n19917 , n19915 , n19916 );
nor ( n19918 , n19914 , n19917 );
xor ( n19919 , n19909 , n19918 );
buf ( n19920 , n6123 );
nand ( n19921 , n14573 , n19920 );
buf ( n19922 , n6124 );
not ( n19923 , n19922 );
and ( n19924 , n19921 , n19923 );
not ( n19925 , n19921 );
buf ( n19926 , n19922 );
and ( n19927 , n19925 , n19926 );
nor ( n19928 , n19924 , n19927 );
xnor ( n19929 , n19919 , n19928 );
not ( n19930 , n19929 );
not ( n19931 , n19930 );
or ( n19932 , n19896 , n19931 );
or ( n19933 , n19930 , n19895 );
nand ( n19934 , n19932 , n19933 );
not ( n19935 , n12899 );
buf ( n19936 , n6125 );
not ( n19937 , n19936 );
not ( n19938 , n19937 );
or ( n19939 , n19935 , n19938 );
not ( n19940 , n12898 );
buf ( n19941 , n19936 );
nand ( n19942 , n19940 , n19941 );
nand ( n19943 , n19939 , n19942 );
buf ( n19944 , n6126 );
not ( n19945 , n19944 );
and ( n19946 , n19943 , n19945 );
not ( n19947 , n19943 );
buf ( n19948 , n19944 );
and ( n19949 , n19947 , n19948 );
nor ( n19950 , n19946 , n19949 );
buf ( n19951 , n6127 );
nand ( n19952 , n7977 , n19951 );
buf ( n19953 , n6128 );
buf ( n19954 , n19953 );
and ( n19955 , n19952 , n19954 );
not ( n19956 , n19952 );
not ( n19957 , n19953 );
and ( n19958 , n19956 , n19957 );
nor ( n19959 , n19955 , n19958 );
xor ( n19960 , n19950 , n19959 );
buf ( n19961 , n6129 );
nand ( n19962 , n6816 , n19961 );
buf ( n19963 , n6130 );
not ( n19964 , n19963 );
and ( n19965 , n19962 , n19964 );
not ( n19966 , n19962 );
buf ( n19967 , n19963 );
and ( n19968 , n19966 , n19967 );
nor ( n19969 , n19965 , n19968 );
xnor ( n19970 , n19960 , n19969 );
not ( n19971 , n19970 );
not ( n19972 , n19971 );
xor ( n19973 , n19934 , n19972 );
nand ( n19974 , n19894 , n19973 );
not ( n19975 , n19974 );
or ( n19976 , n19883 , n19975 );
or ( n19977 , n19882 , n19974 );
nand ( n19978 , n19976 , n19977 );
not ( n19979 , n19978 );
buf ( n19980 , n6131 );
nand ( n19981 , n6577 , n19980 );
buf ( n19982 , n6132 );
buf ( n19983 , n19982 );
and ( n19984 , n19981 , n19983 );
not ( n19985 , n19981 );
not ( n19986 , n19982 );
and ( n19987 , n19985 , n19986 );
nor ( n19988 , n19984 , n19987 );
buf ( n19989 , n19988 );
and ( n19990 , n19989 , n10749 );
not ( n19991 , n19989 );
and ( n19992 , n19991 , n10744 );
nor ( n19993 , n19990 , n19992 );
not ( n19994 , n19993 );
and ( n19995 , n9067 , n19994 );
not ( n19996 , n9067 );
and ( n19997 , n19996 , n19993 );
nor ( n19998 , n19995 , n19997 );
not ( n19999 , n10252 );
buf ( n20000 , n6133 );
buf ( n20001 , n20000 );
not ( n20002 , n20001 );
buf ( n20003 , n6134 );
not ( n20004 , n20003 );
not ( n20005 , n20004 );
or ( n20006 , n20002 , n20005 );
not ( n20007 , n20000 );
buf ( n20008 , n20003 );
nand ( n20009 , n20007 , n20008 );
nand ( n20010 , n20006 , n20009 );
buf ( n20011 , n6135 );
not ( n20012 , n20011 );
and ( n20013 , n20010 , n20012 );
not ( n20014 , n20010 );
buf ( n20015 , n20011 );
and ( n20016 , n20014 , n20015 );
nor ( n20017 , n20013 , n20016 );
buf ( n20018 , n6136 );
nand ( n20019 , n7563 , n20018 );
buf ( n20020 , n6137 );
buf ( n20021 , n20020 );
and ( n20022 , n20019 , n20021 );
not ( n20023 , n20019 );
not ( n20024 , n20020 );
and ( n20025 , n20023 , n20024 );
nor ( n20026 , n20022 , n20025 );
xor ( n20027 , n20017 , n20026 );
buf ( n20028 , n6138 );
nand ( n20029 , n7709 , n20028 );
buf ( n20030 , n6139 );
not ( n20031 , n20030 );
and ( n20032 , n20029 , n20031 );
not ( n20033 , n20029 );
buf ( n20034 , n20030 );
and ( n20035 , n20033 , n20034 );
nor ( n20036 , n20032 , n20035 );
xnor ( n20037 , n20027 , n20036 );
not ( n20038 , n20037 );
not ( n20039 , n20038 );
not ( n20040 , n20039 );
or ( n20041 , n19999 , n20040 );
not ( n20042 , n10252 );
nand ( n20043 , n20042 , n20038 );
nand ( n20044 , n20041 , n20043 );
buf ( n20045 , n6140 );
buf ( n20046 , n20045 );
not ( n20047 , n20046 );
buf ( n20048 , n6141 );
not ( n20049 , n20048 );
not ( n20050 , n20049 );
or ( n20051 , n20047 , n20050 );
not ( n20052 , n20045 );
buf ( n20053 , n20048 );
nand ( n20054 , n20052 , n20053 );
nand ( n20055 , n20051 , n20054 );
and ( n20056 , n20055 , n17356 );
not ( n20057 , n20055 );
not ( n20058 , n17355 );
and ( n20059 , n20057 , n20058 );
nor ( n20060 , n20056 , n20059 );
buf ( n20061 , n6142 );
nand ( n20062 , n6828 , n20061 );
buf ( n20063 , n6143 );
buf ( n20064 , n20063 );
and ( n20065 , n20062 , n20064 );
not ( n20066 , n20062 );
not ( n20067 , n20063 );
and ( n20068 , n20066 , n20067 );
nor ( n20069 , n20065 , n20068 );
xor ( n20070 , n20060 , n20069 );
xor ( n20071 , n20070 , n12167 );
not ( n20072 , n20071 );
not ( n20073 , n20072 );
and ( n20074 , n20044 , n20073 );
not ( n20075 , n20044 );
xor ( n20076 , n20060 , n12167 );
xnor ( n20077 , n20076 , n20069 );
buf ( n20078 , n20077 );
and ( n20079 , n20075 , n20078 );
nor ( n20080 , n20074 , n20079 );
nand ( n20081 , n19998 , n20080 );
not ( n20082 , n20081 );
not ( n20083 , n19128 );
not ( n20084 , n19156 );
or ( n20085 , n20083 , n20084 );
not ( n20086 , n19156 );
nand ( n20087 , n20086 , n19129 );
nand ( n20088 , n20085 , n20087 );
not ( n20089 , n20088 );
not ( n20090 , n20089 );
not ( n20091 , n12732 );
not ( n20092 , n15833 );
or ( n20093 , n20091 , n20092 );
nand ( n20094 , n15839 , n12729 );
nand ( n20095 , n20093 , n20094 );
not ( n20096 , n20095 );
and ( n20097 , n20090 , n20096 );
and ( n20098 , n20089 , n20095 );
nor ( n20099 , n20097 , n20098 );
not ( n20100 , n20099 );
not ( n20101 , n20100 );
and ( n20102 , n20082 , n20101 );
and ( n20103 , n20081 , n20100 );
nor ( n20104 , n20102 , n20103 );
not ( n20105 , n20104 );
not ( n20106 , n20105 );
not ( n20107 , n11686 );
not ( n20108 , n20107 );
not ( n20109 , n16796 );
or ( n20110 , n20108 , n20109 );
not ( n20111 , n20107 );
nand ( n20112 , n20111 , n16795 );
nand ( n20113 , n20110 , n20112 );
and ( n20114 , n20113 , n16804 );
not ( n20115 , n20113 );
and ( n20116 , n20115 , n16801 );
nor ( n20117 , n20114 , n20116 );
not ( n20118 , n20117 );
buf ( n20119 , n9978 );
not ( n20120 , n20119 );
buf ( n20121 , n17095 );
not ( n20122 , n20121 );
buf ( n20123 , n6144 );
not ( n20124 , n20123 );
not ( n20125 , n20124 );
or ( n20126 , n20122 , n20125 );
buf ( n20127 , n20123 );
nand ( n20128 , n17096 , n20127 );
nand ( n20129 , n20126 , n20128 );
and ( n20130 , n20129 , n15115 );
not ( n20131 , n20129 );
buf ( n20132 , n15114 );
and ( n20133 , n20131 , n20132 );
nor ( n20134 , n20130 , n20133 );
buf ( n20135 , n6145 );
nand ( n20136 , n8781 , n20135 );
buf ( n20137 , n6146 );
not ( n20138 , n20137 );
and ( n20139 , n20136 , n20138 );
not ( n20140 , n20136 );
buf ( n20141 , n20137 );
and ( n20142 , n20140 , n20141 );
nor ( n20143 , n20139 , n20142 );
xor ( n20144 , n20134 , n20143 );
buf ( n20145 , n6147 );
nand ( n20146 , n10570 , n20145 );
buf ( n20147 , n6148 );
not ( n20148 , n20147 );
and ( n20149 , n20146 , n20148 );
not ( n20150 , n20146 );
buf ( n20151 , n20147 );
and ( n20152 , n20150 , n20151 );
nor ( n20153 , n20149 , n20152 );
xnor ( n20154 , n20144 , n20153 );
not ( n20155 , n20154 );
or ( n20156 , n20120 , n20155 );
or ( n20157 , n20154 , n20119 );
nand ( n20158 , n20156 , n20157 );
buf ( n20159 , n6149 );
buf ( n20160 , n20159 );
not ( n20161 , n20160 );
buf ( n20162 , n6150 );
not ( n20163 , n20162 );
not ( n20164 , n20163 );
or ( n20165 , n20161 , n20164 );
not ( n20166 , n20159 );
buf ( n20167 , n20162 );
nand ( n20168 , n20166 , n20167 );
nand ( n20169 , n20165 , n20168 );
buf ( n20170 , n6151 );
buf ( n20171 , n20170 );
and ( n20172 , n20169 , n20171 );
not ( n20173 , n20169 );
not ( n20174 , n20170 );
and ( n20175 , n20173 , n20174 );
nor ( n20176 , n20172 , n20175 );
buf ( n20177 , n6152 );
nand ( n20178 , n8781 , n20177 );
buf ( n20179 , n6153 );
not ( n20180 , n20179 );
and ( n20181 , n20178 , n20180 );
not ( n20182 , n20178 );
buf ( n20183 , n20179 );
and ( n20184 , n20182 , n20183 );
nor ( n20185 , n20181 , n20184 );
xor ( n20186 , n20176 , n20185 );
buf ( n20187 , n6154 );
nand ( n20188 , n14573 , n20187 );
buf ( n20189 , n6155 );
not ( n20190 , n20189 );
and ( n20191 , n20188 , n20190 );
not ( n20192 , n20188 );
buf ( n20193 , n20189 );
and ( n20194 , n20192 , n20193 );
nor ( n20195 , n20191 , n20194 );
xnor ( n20196 , n20186 , n20195 );
not ( n20197 , n20196 );
not ( n20198 , n20197 );
not ( n20199 , n20198 );
and ( n20200 , n20158 , n20199 );
not ( n20201 , n20158 );
not ( n20202 , n20196 );
not ( n20203 , n20202 );
and ( n20204 , n20201 , n20203 );
nor ( n20205 , n20200 , n20204 );
nand ( n20206 , n20118 , n20205 );
not ( n20207 , n11734 );
buf ( n20208 , n17957 );
not ( n20209 , n20208 );
or ( n20210 , n20207 , n20209 );
or ( n20211 , n20208 , n11734 );
nand ( n20212 , n20210 , n20211 );
and ( n20213 , n20212 , n18003 );
not ( n20214 , n20212 );
and ( n20215 , n20214 , n18004 );
nor ( n20216 , n20213 , n20215 );
buf ( n20217 , n20216 );
xor ( n20218 , n20206 , n20217 );
not ( n20219 , n20218 );
not ( n20220 , n20219 );
or ( n20221 , n20106 , n20220 );
nand ( n20222 , n20218 , n20104 );
nand ( n20223 , n20221 , n20222 );
not ( n20224 , n16093 );
not ( n20225 , n18015 );
or ( n20226 , n20224 , n20225 );
not ( n20227 , n16093 );
nand ( n20228 , n20227 , n14151 );
nand ( n20229 , n20226 , n20228 );
xor ( n20230 , n11670 , n11638 );
xnor ( n20231 , n20230 , n11648 );
buf ( n20232 , n20231 );
xnor ( n20233 , n20229 , n20232 );
buf ( n20234 , n6156 );
nand ( n20235 , n6828 , n20234 );
buf ( n20236 , n6157 );
buf ( n20237 , n20236 );
and ( n20238 , n20235 , n20237 );
not ( n20239 , n20235 );
not ( n20240 , n20236 );
and ( n20241 , n20239 , n20240 );
nor ( n20242 , n20238 , n20241 );
buf ( n20243 , n20242 );
not ( n20244 , n20243 );
buf ( n20245 , n6158 );
buf ( n20246 , n20245 );
not ( n20247 , n20246 );
buf ( n20248 , n6159 );
not ( n20249 , n20248 );
not ( n20250 , n20249 );
or ( n20251 , n20247 , n20250 );
not ( n20252 , n20245 );
buf ( n20253 , n20248 );
nand ( n20254 , n20252 , n20253 );
nand ( n20255 , n20251 , n20254 );
buf ( n20256 , n6160 );
buf ( n20257 , n20256 );
and ( n20258 , n20255 , n20257 );
not ( n20259 , n20255 );
not ( n20260 , n20256 );
and ( n20261 , n20259 , n20260 );
nor ( n20262 , n20258 , n20261 );
buf ( n20263 , n6161 );
nand ( n20264 , n8364 , n20263 );
buf ( n20265 , n6162 );
not ( n20266 , n20265 );
and ( n20267 , n20264 , n20266 );
not ( n20268 , n20264 );
buf ( n20269 , n20265 );
and ( n20270 , n20268 , n20269 );
nor ( n20271 , n20267 , n20270 );
xor ( n20272 , n20262 , n20271 );
xnor ( n20273 , n20272 , n11366 );
not ( n20274 , n20273 );
not ( n20275 , n20274 );
or ( n20276 , n20244 , n20275 );
or ( n20277 , n20274 , n20243 );
nand ( n20278 , n20276 , n20277 );
buf ( n20279 , n6163 );
buf ( n20280 , n6164 );
buf ( n20281 , n20280 );
not ( n20282 , n20281 );
buf ( n20283 , n6165 );
not ( n20284 , n20283 );
not ( n20285 , n20284 );
or ( n20286 , n20282 , n20285 );
not ( n20287 , n20280 );
buf ( n20288 , n20283 );
nand ( n20289 , n20287 , n20288 );
nand ( n20290 , n20286 , n20289 );
xor ( n20291 , n20279 , n20290 );
buf ( n20292 , n6166 );
buf ( n20293 , n6167 );
not ( n20294 , n20293 );
xor ( n20295 , n20292 , n20294 );
buf ( n20296 , n6168 );
nand ( n20297 , n6558 , n20296 );
xnor ( n20298 , n20295 , n20297 );
xnor ( n20299 , n20291 , n20298 );
not ( n20300 , n20299 );
not ( n20301 , n20300 );
and ( n20302 , n20278 , n20301 );
not ( n20303 , n20278 );
buf ( n20304 , n20300 );
and ( n20305 , n20303 , n20304 );
nor ( n20306 , n20302 , n20305 );
buf ( n20307 , n20306 );
nand ( n20308 , n20233 , n20307 );
not ( n20309 , n17522 );
not ( n20310 , n13857 );
buf ( n20311 , n6169 );
not ( n20312 , n20311 );
not ( n20313 , n20312 );
or ( n20314 , n20310 , n20313 );
not ( n20315 , n13856 );
buf ( n20316 , n20311 );
nand ( n20317 , n20315 , n20316 );
nand ( n20318 , n20314 , n20317 );
buf ( n20319 , n6170 );
buf ( n20320 , n20319 );
and ( n20321 , n20318 , n20320 );
not ( n20322 , n20318 );
not ( n20323 , n20319 );
and ( n20324 , n20322 , n20323 );
nor ( n20325 , n20321 , n20324 );
xor ( n20326 , n20325 , n9574 );
buf ( n20327 , n6171 );
nand ( n20328 , n9310 , n20327 );
buf ( n20329 , n6172 );
not ( n20330 , n20329 );
and ( n20331 , n20328 , n20330 );
not ( n20332 , n20328 );
buf ( n20333 , n20329 );
and ( n20334 , n20332 , n20333 );
nor ( n20335 , n20331 , n20334 );
xnor ( n20336 , n20326 , n20335 );
buf ( n20337 , n20336 );
buf ( n20338 , n20337 );
not ( n20339 , n20338 );
or ( n20340 , n20309 , n20339 );
not ( n20341 , n20338 );
nand ( n20342 , n20341 , n17519 );
nand ( n20343 , n20340 , n20342 );
buf ( n20344 , n8888 );
not ( n20345 , n20344 );
and ( n20346 , n20343 , n20345 );
not ( n20347 , n20343 );
and ( n20348 , n20347 , n20344 );
nor ( n20349 , n20346 , n20348 );
not ( n20350 , n20349 );
and ( n20351 , n20308 , n20350 );
not ( n20352 , n20308 );
and ( n20353 , n20352 , n20349 );
nor ( n20354 , n20351 , n20353 );
and ( n20355 , n20223 , n20354 );
not ( n20356 , n20223 );
not ( n20357 , n20354 );
and ( n20358 , n20356 , n20357 );
nor ( n20359 , n20355 , n20358 );
not ( n20360 , n20359 );
not ( n20361 , n14800 );
buf ( n20362 , n13277 );
buf ( n20363 , n13273 );
and ( n20364 , n20362 , n20363 );
not ( n20365 , n20362 );
and ( n20366 , n20365 , n13274 );
nor ( n20367 , n20364 , n20366 );
not ( n20368 , n20367 );
buf ( n20369 , n6173 );
buf ( n20370 , n20369 );
not ( n20371 , n20370 );
buf ( n20372 , n6174 );
not ( n20373 , n20372 );
not ( n20374 , n20373 );
or ( n20375 , n20371 , n20374 );
not ( n20376 , n20369 );
buf ( n20377 , n20372 );
nand ( n20378 , n20376 , n20377 );
nand ( n20379 , n20375 , n20378 );
buf ( n20380 , n6175 );
not ( n20381 , n20380 );
and ( n20382 , n20379 , n20381 );
not ( n20383 , n20379 );
buf ( n20384 , n20380 );
and ( n20385 , n20383 , n20384 );
nor ( n20386 , n20382 , n20385 );
buf ( n20387 , n6176 );
nand ( n20388 , n6828 , n20387 );
buf ( n20389 , n6177 );
buf ( n20390 , n20389 );
and ( n20391 , n20388 , n20390 );
not ( n20392 , n20388 );
not ( n20393 , n20389 );
and ( n20394 , n20392 , n20393 );
nor ( n20395 , n20391 , n20394 );
xor ( n20396 , n20386 , n20395 );
buf ( n20397 , n6178 );
nand ( n20398 , n8966 , n20397 );
buf ( n20399 , n6179 );
buf ( n20400 , n20399 );
and ( n20401 , n20398 , n20400 );
not ( n20402 , n20398 );
not ( n20403 , n20399 );
and ( n20404 , n20402 , n20403 );
nor ( n20405 , n20401 , n20404 );
not ( n20406 , n20405 );
xor ( n20407 , n20396 , n20406 );
not ( n20408 , n20407 );
or ( n20409 , n20368 , n20408 );
buf ( n20410 , n20407 );
or ( n20411 , n20410 , n20367 );
nand ( n20412 , n20409 , n20411 );
not ( n20413 , n20412 );
or ( n20414 , n20361 , n20413 );
buf ( n20415 , n14794 );
or ( n20416 , n20412 , n20415 );
nand ( n20417 , n20414 , n20416 );
not ( n20418 , n20417 );
buf ( n20419 , n6180 );
nand ( n20420 , n7709 , n20419 );
buf ( n20421 , n6181 );
not ( n20422 , n20421 );
and ( n20423 , n20420 , n20422 );
not ( n20424 , n20420 );
buf ( n20425 , n20421 );
and ( n20426 , n20424 , n20425 );
nor ( n20427 , n20423 , n20426 );
not ( n20428 , n18082 );
xor ( n20429 , n20427 , n20428 );
xnor ( n20430 , n20429 , n7665 );
not ( n20431 , n20430 );
nand ( n20432 , n20418 , n20431 );
not ( n20433 , n20432 );
not ( n20434 , n11414 );
not ( n20435 , n6792 );
or ( n20436 , n20434 , n20435 );
xor ( n20437 , n6769 , n6789 );
xnor ( n20438 , n20437 , n6779 );
buf ( n20439 , n20438 );
nand ( n20440 , n20439 , n11411 );
nand ( n20441 , n20436 , n20440 );
not ( n20442 , n20441 );
buf ( n20443 , n6182 );
buf ( n20444 , n20443 );
not ( n20445 , n20444 );
buf ( n20446 , n6183 );
not ( n20447 , n20446 );
not ( n20448 , n20447 );
or ( n20449 , n20445 , n20448 );
not ( n20450 , n20443 );
buf ( n20451 , n20446 );
nand ( n20452 , n20450 , n20451 );
nand ( n20453 , n20449 , n20452 );
xor ( n20454 , n19697 , n20453 );
buf ( n20455 , n6184 );
buf ( n20456 , n6185 );
not ( n20457 , n20456 );
xor ( n20458 , n20455 , n20457 );
buf ( n20459 , n6186 );
nand ( n20460 , n6647 , n20459 );
xnor ( n20461 , n20458 , n20460 );
xnor ( n20462 , n20454 , n20461 );
buf ( n20463 , n20462 );
not ( n20464 , n20463 );
not ( n20465 , n20464 );
and ( n20466 , n20442 , n20465 );
and ( n20467 , n20464 , n20441 );
nor ( n20468 , n20466 , n20467 );
not ( n20469 , n20468 );
not ( n20470 , n20469 );
and ( n20471 , n20433 , n20470 );
and ( n20472 , n20432 , n20469 );
nor ( n20473 , n20471 , n20472 );
not ( n20474 , n20473 );
not ( n20475 , n19882 );
not ( n20476 , n19973 );
nand ( n20477 , n20475 , n20476 );
not ( n20478 , n20477 );
buf ( n20479 , n6187 );
buf ( n20480 , n20479 );
not ( n20481 , n20480 );
buf ( n20482 , n6188 );
not ( n20483 , n20482 );
not ( n20484 , n20483 );
or ( n20485 , n20481 , n20484 );
not ( n20486 , n20479 );
buf ( n20487 , n20482 );
nand ( n20488 , n20486 , n20487 );
nand ( n20489 , n20485 , n20488 );
buf ( n20490 , n6189 );
buf ( n20491 , n20490 );
and ( n20492 , n20489 , n20491 );
not ( n20493 , n20489 );
not ( n20494 , n20490 );
and ( n20495 , n20493 , n20494 );
nor ( n20496 , n20492 , n20495 );
buf ( n20497 , n6190 );
nand ( n20498 , n8781 , n20497 );
buf ( n20499 , n6191 );
buf ( n20500 , n20499 );
and ( n20501 , n20498 , n20500 );
not ( n20502 , n20498 );
not ( n20503 , n20499 );
and ( n20504 , n20502 , n20503 );
nor ( n20505 , n20501 , n20504 );
xor ( n20506 , n20496 , n20505 );
buf ( n20507 , n6192 );
nand ( n20508 , n6719 , n20507 );
buf ( n20509 , n6193 );
buf ( n20510 , n20509 );
and ( n20511 , n20508 , n20510 );
not ( n20512 , n20508 );
not ( n20513 , n20509 );
and ( n20514 , n20512 , n20513 );
nor ( n20515 , n20511 , n20514 );
not ( n20516 , n20515 );
xnor ( n20517 , n20506 , n20516 );
buf ( n20518 , n20517 );
xor ( n20519 , n16856 , n20518 );
not ( n20520 , n15874 );
not ( n20521 , n20520 );
buf ( n20522 , n20521 );
xnor ( n20523 , n20519 , n20522 );
not ( n20524 , n20523 );
or ( n20525 , n20478 , n20524 );
or ( n20526 , n20523 , n20477 );
nand ( n20527 , n20525 , n20526 );
not ( n20528 , n20527 );
and ( n20529 , n20474 , n20528 );
and ( n20530 , n20473 , n20527 );
nor ( n20531 , n20529 , n20530 );
not ( n20532 , n20531 );
and ( n20533 , n20360 , n20532 );
not ( n20534 , n20360 );
and ( n20535 , n20534 , n20531 );
nor ( n20536 , n20533 , n20535 );
not ( n20537 , n20536 );
or ( n20538 , n19979 , n20537 );
not ( n20539 , n19978 );
not ( n20540 , n20531 );
not ( n20541 , n20359 );
or ( n20542 , n20540 , n20541 );
nand ( n20543 , n20360 , n20532 );
nand ( n20544 , n20542 , n20543 );
nand ( n20545 , n20539 , n20544 );
nand ( n20546 , n20538 , n20545 );
not ( n20547 , n9756 );
not ( n20548 , n8916 );
or ( n20549 , n20547 , n20548 );
not ( n20550 , n9756 );
nand ( n20551 , n20550 , n8913 );
nand ( n20552 , n20549 , n20551 );
buf ( n20553 , n17411 );
not ( n20554 , n20553 );
and ( n20555 , n20552 , n20554 );
not ( n20556 , n20552 );
buf ( n20557 , n17412 );
not ( n20558 , n20557 );
and ( n20559 , n20556 , n20558 );
nor ( n20560 , n20555 , n20559 );
not ( n20561 , n20560 );
not ( n20562 , n11190 );
xor ( n20563 , n13767 , n13776 );
xor ( n20564 , n20563 , n13784 );
not ( n20565 , n20564 );
not ( n20566 , n20565 );
or ( n20567 , n20562 , n20566 );
not ( n20568 , n11190 );
nand ( n20569 , n20568 , n20564 );
nand ( n20570 , n20567 , n20569 );
buf ( n20571 , n14684 );
not ( n20572 , n20571 );
and ( n20573 , n20570 , n20572 );
not ( n20574 , n20570 );
buf ( n20575 , n14683 );
not ( n20576 , n20575 );
and ( n20577 , n20574 , n20576 );
nor ( n20578 , n20573 , n20577 );
nand ( n20579 , n20561 , n20578 );
not ( n20580 , n20579 );
not ( n20581 , n12218 );
buf ( n20582 , n6194 );
buf ( n20583 , n20582 );
not ( n20584 , n20583 );
buf ( n20585 , n6195 );
not ( n20586 , n20585 );
not ( n20587 , n20586 );
or ( n20588 , n20584 , n20587 );
not ( n20589 , n20582 );
buf ( n20590 , n20585 );
nand ( n20591 , n20589 , n20590 );
nand ( n20592 , n20588 , n20591 );
buf ( n20593 , n6196 );
not ( n20594 , n20593 );
and ( n20595 , n20592 , n20594 );
not ( n20596 , n20592 );
buf ( n20597 , n20593 );
and ( n20598 , n20596 , n20597 );
nor ( n20599 , n20595 , n20598 );
buf ( n20600 , n6197 );
nand ( n20601 , n7014 , n20600 );
buf ( n20602 , n6198 );
buf ( n20603 , n20602 );
and ( n20604 , n20601 , n20603 );
not ( n20605 , n20601 );
not ( n20606 , n20602 );
and ( n20607 , n20605 , n20606 );
nor ( n20608 , n20604 , n20607 );
xor ( n20609 , n20599 , n20608 );
buf ( n20610 , n6199 );
nand ( n20611 , n7344 , n20610 );
buf ( n20612 , n6200 );
buf ( n20613 , n20612 );
and ( n20614 , n20611 , n20613 );
not ( n20615 , n20611 );
not ( n20616 , n20612 );
and ( n20617 , n20615 , n20616 );
nor ( n20618 , n20614 , n20617 );
xor ( n20619 , n20609 , n20618 );
not ( n20620 , n20619 );
or ( n20621 , n20581 , n20620 );
not ( n20622 , n12218 );
xor ( n20623 , n20599 , n20618 );
buf ( n20624 , n20608 );
xnor ( n20625 , n20623 , n20624 );
nand ( n20626 , n20622 , n20625 );
nand ( n20627 , n20621 , n20626 );
buf ( n20628 , n19098 );
and ( n20629 , n20627 , n20628 );
not ( n20630 , n20627 );
buf ( n20631 , n19093 );
and ( n20632 , n20630 , n20631 );
nor ( n20633 , n20629 , n20632 );
not ( n20634 , n20633 );
and ( n20635 , n20580 , n20634 );
and ( n20636 , n20579 , n20633 );
nor ( n20637 , n20635 , n20636 );
xor ( n20638 , n13259 , n13270 );
xnor ( n20639 , n20638 , n13278 );
not ( n20640 , n20639 );
not ( n20641 , n20640 );
not ( n20642 , n7688 );
buf ( n20643 , n6201 );
buf ( n20644 , n20643 );
not ( n20645 , n20644 );
buf ( n20646 , n6202 );
not ( n20647 , n20646 );
not ( n20648 , n20647 );
or ( n20649 , n20645 , n20648 );
not ( n20650 , n20643 );
buf ( n20651 , n20646 );
nand ( n20652 , n20650 , n20651 );
nand ( n20653 , n20649 , n20652 );
buf ( n20654 , n6203 );
buf ( n20655 , n20654 );
and ( n20656 , n20653 , n20655 );
not ( n20657 , n20653 );
not ( n20658 , n20654 );
and ( n20659 , n20657 , n20658 );
nor ( n20660 , n20656 , n20659 );
buf ( n20661 , n6204 );
nand ( n20662 , n6828 , n20661 );
buf ( n20663 , n6205 );
buf ( n20664 , n20663 );
and ( n20665 , n20662 , n20664 );
not ( n20666 , n20662 );
not ( n20667 , n20663 );
and ( n20668 , n20666 , n20667 );
nor ( n20669 , n20665 , n20668 );
xor ( n20670 , n20660 , n20669 );
buf ( n20671 , n6206 );
nand ( n20672 , n6916 , n20671 );
buf ( n20673 , n6207 );
buf ( n20674 , n20673 );
and ( n20675 , n20672 , n20674 );
not ( n20676 , n20672 );
not ( n20677 , n20673 );
and ( n20678 , n20676 , n20677 );
nor ( n20679 , n20675 , n20678 );
not ( n20680 , n20679 );
xor ( n20681 , n20670 , n20680 );
not ( n20682 , n20681 );
or ( n20683 , n20642 , n20682 );
or ( n20684 , n20681 , n7688 );
nand ( n20685 , n20683 , n20684 );
not ( n20686 , n20685 );
or ( n20687 , n20641 , n20686 );
or ( n20688 , n20685 , n20640 );
nand ( n20689 , n20687 , n20688 );
buf ( n20690 , n20689 );
not ( n20691 , n20690 );
buf ( n20692 , n6208 );
buf ( n20693 , n20692 );
not ( n20694 , n20693 );
not ( n20695 , n8234 );
not ( n20696 , n20695 );
or ( n20697 , n20694 , n20696 );
not ( n20698 , n20692 );
nand ( n20699 , n8234 , n20698 );
nand ( n20700 , n20697 , n20699 );
buf ( n20701 , n18560 );
not ( n20702 , n20701 );
and ( n20703 , n20700 , n20702 );
not ( n20704 , n20700 );
and ( n20705 , n20704 , n18573 );
nor ( n20706 , n20703 , n20705 );
nand ( n20707 , n20691 , n20706 );
not ( n20708 , n20707 );
buf ( n20709 , n12890 );
not ( n20710 , n20709 );
not ( n20711 , n6942 );
or ( n20712 , n20710 , n20711 );
or ( n20713 , n6942 , n20709 );
nand ( n20714 , n20712 , n20713 );
and ( n20715 , n20714 , n6893 );
not ( n20716 , n20714 );
and ( n20717 , n20716 , n6892 );
nor ( n20718 , n20715 , n20717 );
not ( n20719 , n20718 );
not ( n20720 , n20719 );
and ( n20721 , n20708 , n20720 );
and ( n20722 , n20707 , n20719 );
nor ( n20723 , n20721 , n20722 );
not ( n20724 , n20723 );
not ( n20725 , n6623 );
not ( n20726 , n10446 );
or ( n20727 , n20725 , n20726 );
not ( n20728 , n6623 );
nand ( n20729 , n20728 , n10443 );
nand ( n20730 , n20727 , n20729 );
buf ( n20731 , n6209 );
nand ( n20732 , n9160 , n20731 );
buf ( n20733 , n6210 );
buf ( n20734 , n20733 );
and ( n20735 , n20732 , n20734 );
not ( n20736 , n20732 );
not ( n20737 , n20733 );
and ( n20738 , n20736 , n20737 );
nor ( n20739 , n20735 , n20738 );
not ( n20740 , n20739 );
buf ( n20741 , n6211 );
nand ( n20742 , n7107 , n20741 );
buf ( n20743 , n6212 );
not ( n20744 , n20743 );
and ( n20745 , n20742 , n20744 );
not ( n20746 , n20742 );
buf ( n20747 , n20743 );
and ( n20748 , n20746 , n20747 );
nor ( n20749 , n20745 , n20748 );
not ( n20750 , n20749 );
or ( n20751 , n20740 , n20750 );
or ( n20752 , n20739 , n20749 );
nand ( n20753 , n20751 , n20752 );
buf ( n20754 , n6213 );
buf ( n20755 , n20754 );
not ( n20756 , n20755 );
buf ( n20757 , n6214 );
not ( n20758 , n20757 );
not ( n20759 , n20758 );
or ( n20760 , n20756 , n20759 );
not ( n20761 , n20754 );
buf ( n20762 , n20757 );
nand ( n20763 , n20761 , n20762 );
nand ( n20764 , n20760 , n20763 );
buf ( n20765 , n6215 );
not ( n20766 , n20765 );
and ( n20767 , n20764 , n20766 );
not ( n20768 , n20764 );
buf ( n20769 , n20765 );
and ( n20770 , n20768 , n20769 );
nor ( n20771 , n20767 , n20770 );
not ( n20772 , n20771 );
and ( n20773 , n20753 , n20772 );
not ( n20774 , n20753 );
and ( n20775 , n20774 , n20771 );
nor ( n20776 , n20773 , n20775 );
not ( n20777 , n20776 );
not ( n20778 , n20777 );
and ( n20779 , n20730 , n20778 );
not ( n20780 , n20730 );
xor ( n20781 , n20771 , n20739 );
xnor ( n20782 , n20781 , n20749 );
not ( n20783 , n20782 );
buf ( n20784 , n20783 );
not ( n20785 , n20784 );
and ( n20786 , n20780 , n20785 );
nor ( n20787 , n20779 , n20786 );
not ( n20788 , n20787 );
not ( n20789 , n13963 );
buf ( n20790 , n6216 );
buf ( n20791 , n20790 );
not ( n20792 , n20791 );
buf ( n20793 , n6217 );
not ( n20794 , n20793 );
not ( n20795 , n20794 );
or ( n20796 , n20792 , n20795 );
not ( n20797 , n20790 );
buf ( n20798 , n20793 );
nand ( n20799 , n20797 , n20798 );
nand ( n20800 , n20796 , n20799 );
buf ( n20801 , n6218 );
buf ( n20802 , n20801 );
and ( n20803 , n20800 , n20802 );
not ( n20804 , n20800 );
not ( n20805 , n20801 );
and ( n20806 , n20804 , n20805 );
nor ( n20807 , n20803 , n20806 );
buf ( n20808 , n6219 );
nand ( n20809 , n9160 , n20808 );
buf ( n20810 , n6220 );
buf ( n20811 , n20810 );
and ( n20812 , n20809 , n20811 );
not ( n20813 , n20809 );
not ( n20814 , n20810 );
and ( n20815 , n20813 , n20814 );
nor ( n20816 , n20812 , n20815 );
xor ( n20817 , n20807 , n20816 );
buf ( n20818 , n6221 );
nand ( n20819 , n8323 , n20818 );
buf ( n20820 , n6222 );
not ( n20821 , n20820 );
and ( n20822 , n20819 , n20821 );
not ( n20823 , n20819 );
buf ( n20824 , n20820 );
and ( n20825 , n20823 , n20824 );
nor ( n20826 , n20822 , n20825 );
xor ( n20827 , n20817 , n20826 );
not ( n20828 , n20827 );
not ( n20829 , n20828 );
not ( n20830 , n20829 );
or ( n20831 , n20789 , n20830 );
or ( n20832 , n20829 , n13963 );
nand ( n20833 , n20831 , n20832 );
and ( n20834 , n20833 , n19293 );
not ( n20835 , n20833 );
not ( n20836 , n19290 );
not ( n20837 , n20836 );
and ( n20838 , n20835 , n20837 );
nor ( n20839 , n20834 , n20838 );
nand ( n20840 , n20788 , n20839 );
not ( n20841 , n20840 );
xor ( n20842 , n16490 , n16009 );
not ( n20843 , n15937 );
xor ( n20844 , n15969 , n20843 );
xnor ( n20845 , n20844 , n18168 );
buf ( n20846 , n20845 );
xnor ( n20847 , n20842 , n20846 );
not ( n20848 , n20847 );
not ( n20849 , n20848 );
and ( n20850 , n20841 , n20849 );
and ( n20851 , n20840 , n20848 );
nor ( n20852 , n20850 , n20851 );
not ( n20853 , n20852 );
not ( n20854 , n20853 );
or ( n20855 , n20724 , n20854 );
not ( n20856 , n20723 );
nand ( n20857 , n20856 , n20852 );
nand ( n20858 , n20855 , n20857 );
xor ( n20859 , n20637 , n20858 );
not ( n20860 , n18926 );
not ( n20861 , n13457 );
or ( n20862 , n20860 , n20861 );
nand ( n20863 , n9989 , n18922 );
nand ( n20864 , n20862 , n20863 );
not ( n20865 , n20864 );
buf ( n20866 , n13832 );
not ( n20867 , n20866 );
and ( n20868 , n20865 , n20867 );
and ( n20869 , n20864 , n20866 );
nor ( n20870 , n20868 , n20869 );
and ( n20871 , n9283 , n16658 );
not ( n20872 , n9283 );
not ( n20873 , n16658 );
and ( n20874 , n20872 , n20873 );
nor ( n20875 , n20871 , n20874 );
and ( n20876 , n20875 , n16685 );
not ( n20877 , n20875 );
not ( n20878 , n16681 );
and ( n20879 , n20877 , n20878 );
nor ( n20880 , n20876 , n20879 );
not ( n20881 , n20880 );
nand ( n20882 , n20870 , n20881 );
buf ( n20883 , n15171 );
not ( n20884 , n20883 );
not ( n20885 , n19821 );
or ( n20886 , n20884 , n20885 );
or ( n20887 , n19826 , n20883 );
nand ( n20888 , n20886 , n20887 );
and ( n20889 , n20888 , n19829 );
not ( n20890 , n20888 );
and ( n20891 , n20890 , n19833 );
nor ( n20892 , n20889 , n20891 );
not ( n20893 , n20892 );
and ( n20894 , n20882 , n20893 );
not ( n20895 , n20882 );
and ( n20896 , n20895 , n20892 );
nor ( n20897 , n20894 , n20896 );
not ( n20898 , n20897 );
not ( n20899 , n20898 );
buf ( n20900 , n6223 );
buf ( n20901 , n20900 );
not ( n20902 , n20901 );
not ( n20903 , n12375 );
not ( n20904 , n20903 );
or ( n20905 , n20902 , n20904 );
not ( n20906 , n20901 );
nand ( n20907 , n20906 , n19006 );
nand ( n20908 , n20905 , n20907 );
not ( n20909 , n19045 );
and ( n20910 , n20908 , n20909 );
not ( n20911 , n20908 );
not ( n20912 , n19041 );
not ( n20913 , n20912 );
and ( n20914 , n20911 , n20913 );
nor ( n20915 , n20910 , n20914 );
not ( n20916 , n7963 );
not ( n20917 , n14540 );
not ( n20918 , n20917 );
or ( n20919 , n20916 , n20918 );
or ( n20920 , n20917 , n7963 );
nand ( n20921 , n20919 , n20920 );
and ( n20922 , n20921 , n15701 );
not ( n20923 , n20921 );
and ( n20924 , n20923 , n14508 );
nor ( n20925 , n20922 , n20924 );
buf ( n20926 , n20925 );
nand ( n20927 , n20915 , n20926 );
not ( n20928 , n20927 );
buf ( n20929 , n11435 );
and ( n20930 , n20929 , n6791 );
not ( n20931 , n20929 );
and ( n20932 , n20931 , n20438 );
nor ( n20933 , n20930 , n20932 );
not ( n20934 , n20933 );
not ( n20935 , n20462 );
or ( n20936 , n20934 , n20935 );
not ( n20937 , n20462 );
not ( n20938 , n20937 );
or ( n20939 , n20938 , n20933 );
nand ( n20940 , n20936 , n20939 );
buf ( n20941 , n20940 );
not ( n20942 , n20941 );
and ( n20943 , n20928 , n20942 );
and ( n20944 , n20927 , n20941 );
nor ( n20945 , n20943 , n20944 );
not ( n20946 , n20945 );
not ( n20947 , n20946 );
or ( n20948 , n20899 , n20947 );
nand ( n20949 , n20945 , n20897 );
nand ( n20950 , n20948 , n20949 );
xor ( n20951 , n20859 , n20950 );
buf ( n20952 , n20951 );
and ( n20953 , n20546 , n20952 );
not ( n20954 , n20546 );
not ( n20955 , n20858 );
not ( n20956 , n20955 );
not ( n20957 , n20637 );
and ( n20958 , n20950 , n20957 );
not ( n20959 , n20950 );
and ( n20960 , n20959 , n20637 );
nor ( n20961 , n20958 , n20960 );
not ( n20962 , n20961 );
or ( n20963 , n20956 , n20962 );
not ( n20964 , n20961 );
nand ( n20965 , n20964 , n20858 );
nand ( n20966 , n20963 , n20965 );
buf ( n20967 , n20966 );
and ( n20968 , n20954 , n20967 );
nor ( n20969 , n20953 , n20968 );
not ( n20970 , n20969 );
and ( n20971 , n19869 , n20970 );
not ( n20972 , n19869 );
and ( n20973 , n20972 , n20969 );
nor ( n20974 , n20971 , n20973 );
buf ( n20975 , n15324 );
buf ( n20976 , n20975 );
buf ( n20977 , n20976 );
or ( n20978 , n20974 , n20977 );
nand ( n20979 , n17822 , n20978 );
buf ( n20980 , n20979 );
buf ( n20981 , n20980 );
not ( n20982 , n15207 );
buf ( n20983 , n13352 );
buf ( n20984 , n20983 );
not ( n20985 , n20984 );
or ( n20986 , n20982 , n20985 );
buf ( n20987 , n14435 );
not ( n20988 , n20987 );
not ( n20989 , n20988 );
not ( n20990 , n8186 );
or ( n20991 , n20989 , n20990 );
nand ( n20992 , n8192 , n20987 );
nand ( n20993 , n20991 , n20992 );
not ( n20994 , n20993 );
not ( n20995 , n8233 );
not ( n20996 , n20995 );
and ( n20997 , n20994 , n20996 );
and ( n20998 , n20993 , n20995 );
nor ( n20999 , n20997 , n20998 );
not ( n21000 , n20999 );
nand ( n21001 , n10404 , n21000 );
not ( n21002 , n21001 );
not ( n21003 , n10316 );
not ( n21004 , n21003 );
or ( n21005 , n21002 , n21004 );
or ( n21006 , n21003 , n21001 );
nand ( n21007 , n21005 , n21006 );
not ( n21008 , n21007 );
not ( n21009 , n10463 );
or ( n21010 , n21008 , n21009 );
not ( n21011 , n21007 );
nand ( n21012 , n21011 , n10472 );
nand ( n21013 , n21010 , n21012 );
and ( n21014 , n21013 , n11293 );
not ( n21015 , n21013 );
and ( n21016 , n21015 , n11302 );
nor ( n21017 , n21014 , n21016 );
not ( n21018 , n21017 );
not ( n21019 , n9518 );
not ( n21020 , n21019 );
not ( n21021 , n18129 );
not ( n21022 , n16147 );
or ( n21023 , n21021 , n21022 );
or ( n21024 , n16147 , n18129 );
nand ( n21025 , n21023 , n21024 );
not ( n21026 , n21025 );
or ( n21027 , n21020 , n21026 );
or ( n21028 , n21025 , n21019 );
nand ( n21029 , n21027 , n21028 );
not ( n21030 , n21029 );
not ( n21031 , n13550 );
buf ( n21032 , n6224 );
nand ( n21033 , n8675 , n21032 );
buf ( n21034 , n6225 );
buf ( n21035 , n21034 );
and ( n21036 , n21033 , n21035 );
not ( n21037 , n21033 );
not ( n21038 , n21034 );
and ( n21039 , n21037 , n21038 );
nor ( n21040 , n21036 , n21039 );
buf ( n21041 , n21040 );
not ( n21042 , n21041 );
not ( n21043 , n21042 );
not ( n21044 , n13591 );
or ( n21045 , n21043 , n21044 );
nand ( n21046 , n13595 , n21041 );
nand ( n21047 , n21045 , n21046 );
not ( n21048 , n21047 );
and ( n21049 , n21031 , n21048 );
and ( n21050 , n13550 , n21047 );
nor ( n21051 , n21049 , n21050 );
not ( n21052 , n21051 );
nand ( n21053 , n21030 , n21052 );
not ( n21054 , n21053 );
not ( n21055 , n9099 );
not ( n21056 , n19199 );
or ( n21057 , n21055 , n21056 );
or ( n21058 , n19199 , n9099 );
nand ( n21059 , n21057 , n21058 );
buf ( n21060 , n19662 );
and ( n21061 , n21059 , n21060 );
not ( n21062 , n21059 );
buf ( n21063 , n19666 );
and ( n21064 , n21062 , n21063 );
nor ( n21065 , n21061 , n21064 );
not ( n21066 , n21065 );
not ( n21067 , n21066 );
and ( n21068 , n21054 , n21067 );
and ( n21069 , n21053 , n21066 );
nor ( n21070 , n21068 , n21069 );
not ( n21071 , n21070 );
nand ( n21072 , n21065 , n21029 );
not ( n21073 , n21072 );
not ( n21074 , n12206 );
not ( n21075 , n20053 );
not ( n21076 , n12216 );
or ( n21077 , n21075 , n21076 );
or ( n21078 , n12216 , n20053 );
nand ( n21079 , n21077 , n21078 );
not ( n21080 , n21079 );
not ( n21081 , n12231 );
not ( n21082 , n21081 );
or ( n21083 , n21080 , n21082 );
or ( n21084 , n21081 , n21079 );
nand ( n21085 , n21083 , n21084 );
not ( n21086 , n21085 );
and ( n21087 , n21074 , n21086 );
and ( n21088 , n21085 , n12206 );
nor ( n21089 , n21087 , n21088 );
not ( n21090 , n21089 );
not ( n21091 , n21090 );
and ( n21092 , n21073 , n21091 );
and ( n21093 , n21072 , n21090 );
nor ( n21094 , n21092 , n21093 );
not ( n21095 , n21094 );
buf ( n21096 , n6226 );
buf ( n21097 , n21096 );
not ( n21098 , n21097 );
not ( n21099 , n8042 );
or ( n21100 , n21098 , n21099 );
or ( n21101 , n8042 , n21097 );
nand ( n21102 , n21100 , n21101 );
not ( n21103 , n21102 );
not ( n21104 , n21103 );
not ( n21105 , n7992 );
or ( n21106 , n21104 , n21105 );
nand ( n21107 , n7993 , n21102 );
nand ( n21108 , n21106 , n21107 );
not ( n21109 , n21108 );
not ( n21110 , n14092 );
not ( n21111 , n21110 );
not ( n21112 , n6668 );
and ( n21113 , n21111 , n21112 );
and ( n21114 , n21110 , n6668 );
nor ( n21115 , n21113 , n21114 );
buf ( n21116 , n6227 );
buf ( n21117 , n21116 );
not ( n21118 , n21117 );
buf ( n21119 , n6228 );
not ( n21120 , n21119 );
not ( n21121 , n21120 );
or ( n21122 , n21118 , n21121 );
not ( n21123 , n21116 );
buf ( n21124 , n21119 );
nand ( n21125 , n21123 , n21124 );
nand ( n21126 , n21122 , n21125 );
buf ( n21127 , n6229 );
not ( n21128 , n21127 );
and ( n21129 , n21126 , n21128 );
not ( n21130 , n21126 );
buf ( n21131 , n21127 );
and ( n21132 , n21130 , n21131 );
nor ( n21133 , n21129 , n21132 );
xor ( n21134 , n21133 , n16298 );
buf ( n21135 , n6230 );
nand ( n21136 , n10165 , n21135 );
buf ( n21137 , n6231 );
buf ( n21138 , n21137 );
and ( n21139 , n21136 , n21138 );
not ( n21140 , n21136 );
not ( n21141 , n21137 );
and ( n21142 , n21140 , n21141 );
nor ( n21143 , n21139 , n21142 );
not ( n21144 , n21143 );
xnor ( n21145 , n21134 , n21144 );
buf ( n21146 , n21145 );
and ( n21147 , n21115 , n21146 );
not ( n21148 , n21115 );
not ( n21149 , n21145 );
and ( n21150 , n21148 , n21149 );
nor ( n21151 , n21147 , n21150 );
nand ( n21152 , n21109 , n21151 );
not ( n21153 , n20089 );
and ( n21154 , n12725 , n15833 );
not ( n21155 , n12725 );
and ( n21156 , n21155 , n15839 );
nor ( n21157 , n21154 , n21156 );
not ( n21158 , n21157 );
not ( n21159 , n21158 );
or ( n21160 , n21153 , n21159 );
nand ( n21161 , n21157 , n20088 );
nand ( n21162 , n21160 , n21161 );
not ( n21163 , n21162 );
and ( n21164 , n21152 , n21163 );
not ( n21165 , n21152 );
and ( n21166 , n21165 , n21162 );
nor ( n21167 , n21164 , n21166 );
not ( n21168 , n21167 );
or ( n21169 , n21095 , n21168 );
or ( n21170 , n21167 , n21094 );
nand ( n21171 , n21169 , n21170 );
not ( n21172 , n12505 );
not ( n21173 , n10126 );
or ( n21174 , n21172 , n21173 );
not ( n21175 , n12505 );
nand ( n21176 , n21175 , n10491 );
nand ( n21177 , n21174 , n21176 );
not ( n21178 , n21177 );
not ( n21179 , n18528 );
and ( n21180 , n21178 , n21179 );
and ( n21181 , n21177 , n18528 );
nor ( n21182 , n21180 , n21181 );
buf ( n21183 , n6232 );
buf ( n21184 , n21183 );
nor ( n21185 , n7923 , n21184 );
not ( n21186 , n21185 );
nand ( n21187 , n7927 , n21184 );
nand ( n21188 , n21186 , n21187 );
not ( n21189 , n7879 );
and ( n21190 , n21188 , n21189 );
not ( n21191 , n21188 );
and ( n21192 , n21191 , n7879 );
nor ( n21193 , n21190 , n21192 );
nand ( n21194 , n21182 , n21193 );
not ( n21195 , n20451 );
not ( n21196 , n12636 );
or ( n21197 , n21195 , n21196 );
or ( n21198 , n12636 , n20451 );
nand ( n21199 , n21197 , n21198 );
buf ( n21200 , n19747 );
and ( n21201 , n21199 , n21200 );
not ( n21202 , n21199 );
buf ( n21203 , n19739 );
and ( n21204 , n21202 , n21203 );
nor ( n21205 , n21201 , n21204 );
not ( n21206 , n21205 );
and ( n21207 , n21194 , n21206 );
not ( n21208 , n21194 );
and ( n21209 , n21208 , n21205 );
nor ( n21210 , n21207 , n21209 );
and ( n21211 , n21171 , n21210 );
not ( n21212 , n21171 );
not ( n21213 , n21210 );
and ( n21214 , n21212 , n21213 );
nor ( n21215 , n21211 , n21214 );
not ( n21216 , n21215 );
not ( n21217 , n15291 );
xor ( n21218 , n19328 , n21217 );
buf ( n21219 , n6233 );
buf ( n21220 , n21219 );
not ( n21221 , n21220 );
buf ( n21222 , n6234 );
not ( n21223 , n21222 );
not ( n21224 , n21223 );
or ( n21225 , n21221 , n21224 );
not ( n21226 , n21219 );
buf ( n21227 , n21222 );
nand ( n21228 , n21226 , n21227 );
nand ( n21229 , n21225 , n21228 );
not ( n21230 , n21229 );
buf ( n21231 , n6235 );
nand ( n21232 , n6634 , n21231 );
buf ( n21233 , n6236 );
buf ( n21234 , n21233 );
and ( n21235 , n21232 , n21234 );
not ( n21236 , n21232 );
not ( n21237 , n21233 );
and ( n21238 , n21236 , n21237 );
nor ( n21239 , n21235 , n21238 );
not ( n21240 , n21239 );
buf ( n21241 , n6237 );
nand ( n21242 , n6647 , n21241 );
buf ( n21243 , n6238 );
buf ( n21244 , n21243 );
and ( n21245 , n21242 , n21244 );
not ( n21246 , n21242 );
not ( n21247 , n21243 );
and ( n21248 , n21246 , n21247 );
nor ( n21249 , n21245 , n21248 );
not ( n21250 , n21249 );
not ( n21251 , n21250 );
or ( n21252 , n21240 , n21251 );
not ( n21253 , n21239 );
nand ( n21254 , n21249 , n21253 );
nand ( n21255 , n21252 , n21254 );
buf ( n21256 , n6239 );
buf ( n21257 , n21256 );
and ( n21258 , n21255 , n21257 );
not ( n21259 , n21255 );
not ( n21260 , n21256 );
and ( n21261 , n21259 , n21260 );
nor ( n21262 , n21258 , n21261 );
and ( n21263 , n21230 , n21262 );
not ( n21264 , n21230 );
not ( n21265 , n21262 );
and ( n21266 , n21264 , n21265 );
nor ( n21267 , n21263 , n21266 );
not ( n21268 , n21267 );
xnor ( n21269 , n21218 , n21268 );
not ( n21270 , n11307 );
not ( n21271 , n21270 );
not ( n21272 , n8524 );
not ( n21273 , n11348 );
or ( n21274 , n21272 , n21273 );
or ( n21275 , n11348 , n8524 );
nand ( n21276 , n21274 , n21275 );
not ( n21277 , n21276 );
or ( n21278 , n21271 , n21277 );
or ( n21279 , n21276 , n21270 );
nand ( n21280 , n21278 , n21279 );
nand ( n21281 , n21269 , n21280 );
not ( n21282 , n21281 );
not ( n21283 , n13246 );
not ( n21284 , n14794 );
or ( n21285 , n21283 , n21284 );
nand ( n21286 , n14799 , n13242 );
nand ( n21287 , n21285 , n21286 );
not ( n21288 , n21287 );
not ( n21289 , n14847 );
and ( n21290 , n21288 , n21289 );
and ( n21291 , n21287 , n14847 );
nor ( n21292 , n21290 , n21291 );
not ( n21293 , n21292 );
not ( n21294 , n21293 );
and ( n21295 , n21282 , n21294 );
nand ( n21296 , n21269 , n21280 );
and ( n21297 , n21296 , n21293 );
nor ( n21298 , n21295 , n21297 );
not ( n21299 , n21298 );
buf ( n21300 , n6240 );
buf ( n21301 , n21300 );
xor ( n21302 , n21301 , n20428 );
not ( n21303 , n7665 );
not ( n21304 , n21303 );
xor ( n21305 , n21302 , n21304 );
not ( n21306 , n14564 );
not ( n21307 , n7720 );
or ( n21308 , n21306 , n21307 );
not ( n21309 , n7719 );
nand ( n21310 , n21309 , n14558 );
nand ( n21311 , n21308 , n21310 );
not ( n21312 , n21311 );
not ( n21313 , n15237 );
not ( n21314 , n21313 );
and ( n21315 , n21312 , n21314 );
and ( n21316 , n21311 , n21313 );
nor ( n21317 , n21315 , n21316 );
nand ( n21318 , n21305 , n21317 );
not ( n21319 , n17098 );
not ( n21320 , n21319 );
not ( n21321 , n21320 );
buf ( n21322 , n6241 );
buf ( n21323 , n21322 );
not ( n21324 , n21323 );
buf ( n21325 , n6242 );
not ( n21326 , n21325 );
not ( n21327 , n21326 );
or ( n21328 , n21324 , n21327 );
not ( n21329 , n21322 );
buf ( n21330 , n21325 );
nand ( n21331 , n21329 , n21330 );
nand ( n21332 , n21328 , n21331 );
buf ( n21333 , n6243 );
not ( n21334 , n21333 );
and ( n21335 , n21332 , n21334 );
not ( n21336 , n21332 );
buf ( n21337 , n21333 );
and ( n21338 , n21336 , n21337 );
nor ( n21339 , n21335 , n21338 );
buf ( n21340 , n6244 );
nand ( n21341 , n7202 , n21340 );
buf ( n21342 , n6245 );
buf ( n21343 , n21342 );
and ( n21344 , n21341 , n21343 );
not ( n21345 , n21341 );
not ( n21346 , n21342 );
and ( n21347 , n21345 , n21346 );
nor ( n21348 , n21344 , n21347 );
xor ( n21349 , n21339 , n21348 );
buf ( n21350 , n6246 );
nand ( n21351 , n6605 , n21350 );
buf ( n21352 , n6247 );
not ( n21353 , n21352 );
and ( n21354 , n21351 , n21353 );
not ( n21355 , n21351 );
buf ( n21356 , n21352 );
and ( n21357 , n21355 , n21356 );
nor ( n21358 , n21354 , n21357 );
xnor ( n21359 , n21349 , n21358 );
not ( n21360 , n21359 );
not ( n21361 , n21360 );
not ( n21362 , n21361 );
buf ( n21363 , n6248 );
buf ( n21364 , n21363 );
not ( n21365 , n21364 );
and ( n21366 , n21362 , n21365 );
and ( n21367 , n21361 , n21364 );
nor ( n21368 , n21366 , n21367 );
not ( n21369 , n21368 );
and ( n21370 , n21321 , n21369 );
and ( n21371 , n21320 , n21368 );
nor ( n21372 , n21370 , n21371 );
and ( n21373 , n21318 , n21372 );
not ( n21374 , n21318 );
not ( n21375 , n21372 );
and ( n21376 , n21374 , n21375 );
nor ( n21377 , n21373 , n21376 );
not ( n21378 , n21377 );
nand ( n21379 , n21299 , n21378 );
nand ( n21380 , n21298 , n21377 );
nand ( n21381 , n21379 , n21380 );
not ( n21382 , n21381 );
not ( n21383 , n21382 );
or ( n21384 , n21216 , n21383 );
not ( n21385 , n21215 );
nand ( n21386 , n21385 , n21381 );
nand ( n21387 , n21384 , n21386 );
not ( n21388 , n21387 );
or ( n21389 , n21071 , n21388 );
or ( n21390 , n21387 , n21070 );
nand ( n21391 , n21389 , n21390 );
not ( n21392 , n13977 );
not ( n21393 , n20827 );
or ( n21394 , n21392 , n21393 );
not ( n21395 , n13977 );
not ( n21396 , n20827 );
nand ( n21397 , n21395 , n21396 );
nand ( n21398 , n21394 , n21397 );
and ( n21399 , n21398 , n19290 );
not ( n21400 , n21398 );
and ( n21401 , n21400 , n19293 );
nor ( n21402 , n21399 , n21401 );
not ( n21403 , n21402 );
not ( n21404 , n21403 );
not ( n21405 , n14683 );
buf ( n21406 , n11270 );
not ( n21407 , n21406 );
and ( n21408 , n21405 , n21407 );
and ( n21409 , n14683 , n21406 );
nor ( n21410 , n21408 , n21409 );
xor ( n21411 , n14651 , n21410 );
buf ( n21412 , n18705 );
not ( n21413 , n21412 );
not ( n21414 , n10842 );
not ( n21415 , n21414 );
not ( n21416 , n21097 );
buf ( n21417 , n6249 );
not ( n21418 , n21417 );
not ( n21419 , n21418 );
or ( n21420 , n21416 , n21419 );
not ( n21421 , n21096 );
buf ( n21422 , n21417 );
nand ( n21423 , n21421 , n21422 );
nand ( n21424 , n21420 , n21423 );
buf ( n21425 , n6250 );
not ( n21426 , n21425 );
and ( n21427 , n21424 , n21426 );
not ( n21428 , n21424 );
buf ( n21429 , n21425 );
and ( n21430 , n21428 , n21429 );
nor ( n21431 , n21427 , n21430 );
buf ( n21432 , n6251 );
nand ( n21433 , n7606 , n21432 );
buf ( n21434 , n6252 );
buf ( n21435 , n21434 );
and ( n21436 , n21433 , n21435 );
not ( n21437 , n21433 );
not ( n21438 , n21434 );
and ( n21439 , n21437 , n21438 );
nor ( n21440 , n21436 , n21439 );
xor ( n21441 , n21431 , n21440 );
xnor ( n21442 , n21441 , n8002 );
not ( n21443 , n21442 );
not ( n21444 , n21443 );
not ( n21445 , n21444 );
or ( n21446 , n21415 , n21445 );
not ( n21447 , n21442 );
nand ( n21448 , n21447 , n10843 );
nand ( n21449 , n21446 , n21448 );
not ( n21450 , n21449 );
or ( n21451 , n21413 , n21450 );
not ( n21452 , n18705 );
not ( n21453 , n21452 );
or ( n21454 , n21449 , n21453 );
nand ( n21455 , n21451 , n21454 );
nand ( n21456 , n21411 , n21455 );
not ( n21457 , n21456 );
or ( n21458 , n21404 , n21457 );
or ( n21459 , n21456 , n21403 );
nand ( n21460 , n21458 , n21459 );
not ( n21461 , n21460 );
buf ( n21462 , n8535 );
not ( n21463 , n21462 );
not ( n21464 , n11335 );
xor ( n21465 , n11326 , n21464 );
xnor ( n21466 , n21465 , n11346 );
not ( n21467 , n21466 );
or ( n21468 , n21463 , n21467 );
or ( n21469 , n21466 , n21462 );
nand ( n21470 , n21468 , n21469 );
xor ( n21471 , n11307 , n21470 );
buf ( n21472 , n15904 );
not ( n21473 , n21472 );
not ( n21474 , n10036 );
or ( n21475 , n21473 , n21474 );
not ( n21476 , n21472 );
nand ( n21477 , n21476 , n8977 );
nand ( n21478 , n21475 , n21477 );
and ( n21479 , n21478 , n7540 );
not ( n21480 , n21478 );
and ( n21481 , n21480 , n8986 );
nor ( n21482 , n21479 , n21481 );
nand ( n21483 , n21471 , n21482 );
not ( n21484 , n21483 );
not ( n21485 , n10276 );
not ( n21486 , n20077 );
or ( n21487 , n21485 , n21486 );
not ( n21488 , n10276 );
nand ( n21489 , n21488 , n20071 );
nand ( n21490 , n21487 , n21489 );
buf ( n21491 , n16661 );
and ( n21492 , n21490 , n21491 );
not ( n21493 , n21490 );
not ( n21494 , n21491 );
and ( n21495 , n21493 , n21494 );
nor ( n21496 , n21492 , n21495 );
not ( n21497 , n21496 );
and ( n21498 , n21484 , n21497 );
and ( n21499 , n21483 , n21496 );
nor ( n21500 , n21498 , n21499 );
not ( n21501 , n21500 );
or ( n21502 , n21461 , n21501 );
or ( n21503 , n21460 , n21500 );
nand ( n21504 , n21502 , n21503 );
buf ( n21505 , n6253 );
buf ( n21506 , n21505 );
not ( n21507 , n21506 );
not ( n21508 , n7881 );
not ( n21509 , n21508 );
or ( n21510 , n21507 , n21509 );
not ( n21511 , n21505 );
nand ( n21512 , n21511 , n7882 );
nand ( n21513 , n21510 , n21512 );
xor ( n21514 , n21184 , n21513 );
buf ( n21515 , n6254 );
nand ( n21516 , n8537 , n21515 );
buf ( n21517 , n6255 );
buf ( n21518 , n21517 );
and ( n21519 , n21516 , n21518 );
not ( n21520 , n21516 );
not ( n21521 , n21517 );
and ( n21522 , n21520 , n21521 );
nor ( n21523 , n21519 , n21522 );
not ( n21524 , n21523 );
buf ( n21525 , n6256 );
nand ( n21526 , n6815 , n21525 );
buf ( n21527 , n6257 );
buf ( n21528 , n21527 );
and ( n21529 , n21526 , n21528 );
not ( n21530 , n21526 );
not ( n21531 , n21527 );
and ( n21532 , n21530 , n21531 );
nor ( n21533 , n21529 , n21532 );
not ( n21534 , n21533 );
not ( n21535 , n21534 );
or ( n21536 , n21524 , n21535 );
not ( n21537 , n21523 );
nand ( n21538 , n21533 , n21537 );
nand ( n21539 , n21536 , n21538 );
xnor ( n21540 , n21514 , n21539 );
not ( n21541 , n21540 );
buf ( n21542 , n7578 );
not ( n21543 , n21542 );
not ( n21544 , n14942 );
or ( n21545 , n21543 , n21544 );
or ( n21546 , n14942 , n21542 );
nand ( n21547 , n21545 , n21546 );
not ( n21548 , n21547 );
or ( n21549 , n21541 , n21548 );
or ( n21550 , n21547 , n21540 );
nand ( n21551 , n21549 , n21550 );
not ( n21552 , n21551 );
not ( n21553 , n9124 );
not ( n21554 , n19204 );
or ( n21555 , n21553 , n21554 );
or ( n21556 , n19204 , n9124 );
nand ( n21557 , n21555 , n21556 );
and ( n21558 , n21557 , n21060 );
not ( n21559 , n21557 );
and ( n21560 , n21559 , n21063 );
nor ( n21561 , n21558 , n21560 );
not ( n21562 , n21561 );
nand ( n21563 , n21552 , n21562 );
not ( n21564 , n21563 );
not ( n21565 , n17452 );
not ( n21566 , n13445 );
not ( n21567 , n21566 );
or ( n21568 , n21565 , n21567 );
or ( n21569 , n21566 , n17452 );
nand ( n21570 , n21568 , n21569 );
and ( n21571 , n21570 , n17908 );
not ( n21572 , n21570 );
and ( n21573 , n21572 , n13399 );
nor ( n21574 , n21571 , n21573 );
buf ( n21575 , n21574 );
not ( n21576 , n21575 );
and ( n21577 , n21564 , n21576 );
and ( n21578 , n21563 , n21575 );
nor ( n21579 , n21577 , n21578 );
and ( n21580 , n21504 , n21579 );
not ( n21581 , n21504 );
not ( n21582 , n21579 );
and ( n21583 , n21581 , n21582 );
nor ( n21584 , n21580 , n21583 );
not ( n21585 , n21584 );
buf ( n21586 , n6837 );
not ( n21587 , n12591 );
xor ( n21588 , n21586 , n21587 );
xnor ( n21589 , n21588 , n14393 );
not ( n21590 , n21589 );
not ( n21591 , n19589 );
not ( n21592 , n19592 );
or ( n21593 , n21591 , n21592 );
or ( n21594 , n19592 , n19589 );
nand ( n21595 , n21593 , n21594 );
not ( n21596 , n21595 );
buf ( n21597 , n6258 );
buf ( n21598 , n21597 );
not ( n21599 , n21598 );
not ( n21600 , n13596 );
or ( n21601 , n21599 , n21600 );
not ( n21602 , n21597 );
nand ( n21603 , n21602 , n13553 );
nand ( n21604 , n21601 , n21603 );
buf ( n21605 , n6259 );
not ( n21606 , n21605 );
and ( n21607 , n21604 , n21606 );
not ( n21608 , n21604 );
buf ( n21609 , n21605 );
and ( n21610 , n21608 , n21609 );
nor ( n21611 , n21607 , n21610 );
buf ( n21612 , n6260 );
nand ( n21613 , n6577 , n21612 );
buf ( n21614 , n6261 );
buf ( n21615 , n21614 );
and ( n21616 , n21613 , n21615 );
not ( n21617 , n21613 );
not ( n21618 , n21614 );
and ( n21619 , n21617 , n21618 );
nor ( n21620 , n21616 , n21619 );
xor ( n21621 , n21611 , n21620 );
xnor ( n21622 , n21621 , n21040 );
nor ( n21623 , n21596 , n21622 );
not ( n21624 , n21623 );
not ( n21625 , n21595 );
nand ( n21626 , n21625 , n21622 );
nand ( n21627 , n21624 , n21626 );
buf ( n21628 , n11175 );
not ( n21629 , n21628 );
and ( n21630 , n21627 , n21629 );
not ( n21631 , n21627 );
not ( n21632 , n11174 );
and ( n21633 , n21631 , n21632 );
nor ( n21634 , n21630 , n21633 );
not ( n21635 , n21634 );
nand ( n21636 , n21590 , n21635 );
not ( n21637 , n17310 );
not ( n21638 , n12442 );
or ( n21639 , n21637 , n21638 );
or ( n21640 , n12442 , n17310 );
nand ( n21641 , n21639 , n21640 );
and ( n21642 , n21641 , n12462 );
not ( n21643 , n21641 );
and ( n21644 , n21643 , n12466 );
nor ( n21645 , n21642 , n21644 );
xor ( n21646 , n21636 , n21645 );
not ( n21647 , n21646 );
buf ( n21648 , n15974 );
xor ( n21649 , n16474 , n21648 );
not ( n21650 , n16009 );
xnor ( n21651 , n21649 , n21650 );
not ( n21652 , n21651 );
not ( n21653 , n21652 );
xor ( n21654 , n16744 , n21309 );
xor ( n21655 , n21654 , n7756 );
not ( n21656 , n21655 );
buf ( n21657 , n21533 );
not ( n21658 , n21657 );
not ( n21659 , n7926 );
or ( n21660 , n21658 , n21659 );
or ( n21661 , n7926 , n21657 );
nand ( n21662 , n21660 , n21661 );
not ( n21663 , n21662 );
not ( n21664 , n7879 );
and ( n21665 , n21663 , n21664 );
and ( n21666 , n21662 , n7879 );
nor ( n21667 , n21665 , n21666 );
nand ( n21668 , n21656 , n21667 );
not ( n21669 , n21668 );
or ( n21670 , n21653 , n21669 );
not ( n21671 , n21667 );
not ( n21672 , n21671 );
nand ( n21673 , n21672 , n21656 );
or ( n21674 , n21673 , n21652 );
nand ( n21675 , n21670 , n21674 );
not ( n21676 , n21675 );
or ( n21677 , n21647 , n21676 );
or ( n21678 , n21675 , n21646 );
nand ( n21679 , n21677 , n21678 );
not ( n21680 , n21679 );
and ( n21681 , n21585 , n21680 );
and ( n21682 , n21584 , n21679 );
nor ( n21683 , n21681 , n21682 );
buf ( n21684 , n21683 );
buf ( n21685 , n21684 );
and ( n21686 , n21391 , n21685 );
not ( n21687 , n21391 );
not ( n21688 , n21685 );
and ( n21689 , n21687 , n21688 );
nor ( n21690 , n21686 , n21689 );
nand ( n21691 , n21018 , n21690 );
not ( n21692 , n21691 );
not ( n21693 , n13549 );
not ( n21694 , n21693 );
not ( n21695 , n21453 );
not ( n21696 , n10829 );
not ( n21697 , n21447 );
or ( n21698 , n21696 , n21697 );
not ( n21699 , n21447 );
not ( n21700 , n10828 );
nand ( n21701 , n21699 , n21700 );
nand ( n21702 , n21698 , n21701 );
not ( n21703 , n21702 );
or ( n21704 , n21695 , n21703 );
buf ( n21705 , n18705 );
or ( n21706 , n21702 , n21705 );
nand ( n21707 , n21704 , n21706 );
nand ( n21708 , n13602 , n21707 );
not ( n21709 , n21708 );
or ( n21710 , n21694 , n21709 );
or ( n21711 , n21708 , n21693 );
nand ( n21712 , n21710 , n21711 );
not ( n21713 , n21712 );
not ( n21714 , n21713 );
not ( n21715 , n14334 );
not ( n21716 , n21715 );
or ( n21717 , n21714 , n21716 );
not ( n21718 , n14334 );
or ( n21719 , n21718 , n21713 );
nand ( n21720 , n21717 , n21719 );
and ( n21721 , n21720 , n15319 );
not ( n21722 , n21720 );
not ( n21723 , n15313 );
not ( n21724 , n14863 );
or ( n21725 , n21723 , n21724 );
or ( n21726 , n14863 , n15313 );
nand ( n21727 , n21725 , n21726 );
buf ( n21728 , n21727 );
and ( n21729 , n21722 , n21728 );
nor ( n21730 , n21721 , n21729 );
not ( n21731 , n21730 );
not ( n21732 , n21731 );
and ( n21733 , n21692 , n21732 );
and ( n21734 , n21691 , n21731 );
nor ( n21735 , n21733 , n21734 );
not ( n21736 , n15324 );
buf ( n21737 , n21736 );
not ( n21738 , n21737 );
or ( n21739 , n21735 , n21738 );
nand ( n21740 , n20986 , n21739 );
buf ( n21741 , n21740 );
buf ( n21742 , n21741 );
not ( n21743 , n12124 );
buf ( n21744 , n13353 );
not ( n21745 , n21744 );
or ( n21746 , n21743 , n21745 );
buf ( n21747 , n12624 );
not ( n21748 , n21747 );
buf ( n21749 , n6262 );
buf ( n21750 , n21749 );
not ( n21751 , n21750 );
not ( n21752 , n18874 );
or ( n21753 , n21751 , n21752 );
not ( n21754 , n21749 );
nand ( n21755 , n21754 , n18870 );
nand ( n21756 , n21753 , n21755 );
not ( n21757 , n15644 );
and ( n21758 , n21756 , n21757 );
not ( n21759 , n21756 );
and ( n21760 , n21759 , n15645 );
nor ( n21761 , n21758 , n21760 );
buf ( n21762 , n6263 );
nand ( n21763 , n10372 , n21762 );
buf ( n21764 , n6264 );
buf ( n21765 , n21764 );
and ( n21766 , n21763 , n21765 );
not ( n21767 , n21763 );
not ( n21768 , n21764 );
and ( n21769 , n21767 , n21768 );
nor ( n21770 , n21766 , n21769 );
xor ( n21771 , n21761 , n21770 );
xnor ( n21772 , n21771 , n18454 );
not ( n21773 , n21772 );
or ( n21774 , n21748 , n21773 );
or ( n21775 , n21772 , n21747 );
nand ( n21776 , n21774 , n21775 );
not ( n21777 , n21776 );
not ( n21778 , n21777 );
buf ( n21779 , n6265 );
buf ( n21780 , n21779 );
not ( n21781 , n12469 );
buf ( n21782 , n6266 );
buf ( n21783 , n21782 );
and ( n21784 , n21781 , n21783 );
not ( n21785 , n21781 );
not ( n21786 , n21782 );
and ( n21787 , n21785 , n21786 );
nor ( n21788 , n21784 , n21787 );
xor ( n21789 , n21780 , n21788 );
buf ( n21790 , n6267 );
buf ( n21791 , n6268 );
xor ( n21792 , n21790 , n21791 );
buf ( n21793 , n6269 );
nand ( n21794 , n11337 , n21793 );
xnor ( n21795 , n21792 , n21794 );
xnor ( n21796 , n21789 , n21795 );
buf ( n21797 , n21796 );
not ( n21798 , n21797 );
or ( n21799 , n21778 , n21798 );
not ( n21800 , n21779 );
xor ( n21801 , n21800 , n21788 );
xnor ( n21802 , n21801 , n21795 );
buf ( n21803 , n21802 );
nand ( n21804 , n21803 , n21776 );
nand ( n21805 , n21799 , n21804 );
nand ( n21806 , n21805 , n9946 );
not ( n21807 , n21806 );
not ( n21808 , n9846 );
or ( n21809 , n21807 , n21808 );
or ( n21810 , n9846 , n21806 );
nand ( n21811 , n21809 , n21810 );
not ( n21812 , n21811 );
not ( n21813 , n10463 );
or ( n21814 , n21812 , n21813 );
not ( n21815 , n21811 );
nand ( n21816 , n21815 , n10472 );
nand ( n21817 , n21814 , n21816 );
and ( n21818 , n21817 , n11293 );
not ( n21819 , n21817 );
and ( n21820 , n21819 , n11302 );
nor ( n21821 , n21818 , n21820 );
not ( n21822 , n21821 );
xor ( n21823 , n15606 , n14714 );
not ( n21824 , n14755 );
xnor ( n21825 , n21823 , n21824 );
not ( n21826 , n21825 );
not ( n21827 , n21826 );
not ( n21828 , n9915 );
not ( n21829 , n12654 );
buf ( n21830 , n6270 );
not ( n21831 , n21830 );
not ( n21832 , n21831 );
or ( n21833 , n21829 , n21832 );
not ( n21834 , n12653 );
buf ( n21835 , n21830 );
nand ( n21836 , n21834 , n21835 );
nand ( n21837 , n21833 , n21836 );
not ( n21838 , n17472 );
and ( n21839 , n21837 , n21838 );
not ( n21840 , n21837 );
and ( n21841 , n21840 , n17473 );
nor ( n21842 , n21839 , n21841 );
buf ( n21843 , n6271 );
nand ( n21844 , n8454 , n21843 );
buf ( n21845 , n6272 );
buf ( n21846 , n21845 );
and ( n21847 , n21844 , n21846 );
not ( n21848 , n21844 );
not ( n21849 , n21845 );
and ( n21850 , n21848 , n21849 );
nor ( n21851 , n21847 , n21850 );
xor ( n21852 , n21842 , n21851 );
xnor ( n21853 , n21852 , n10626 );
not ( n21854 , n21853 );
not ( n21855 , n21854 );
or ( n21856 , n21828 , n21855 );
buf ( n21857 , n21853 );
nand ( n21858 , n21857 , n9918 );
nand ( n21859 , n21856 , n21858 );
buf ( n21860 , n9598 );
xor ( n21861 , n21859 , n21860 );
not ( n21862 , n7660 );
not ( n21863 , n21862 );
not ( n21864 , n16458 );
not ( n21865 , n21864 );
or ( n21866 , n21863 , n21865 );
or ( n21867 , n21864 , n21862 );
nand ( n21868 , n21866 , n21867 );
not ( n21869 , n16493 );
and ( n21870 , n21868 , n21869 );
not ( n21871 , n21868 );
not ( n21872 , n16497 );
and ( n21873 , n21871 , n21872 );
nor ( n21874 , n21870 , n21873 );
nand ( n21875 , n21861 , n21874 );
not ( n21876 , n21875 );
and ( n21877 , n21827 , n21876 );
and ( n21878 , n21826 , n21875 );
nor ( n21879 , n21877 , n21878 );
not ( n21880 , n21879 );
not ( n21881 , n21880 );
not ( n21882 , n13606 );
buf ( n21883 , n19929 );
not ( n21884 , n21883 );
or ( n21885 , n21882 , n21884 );
not ( n21886 , n13605 );
nand ( n21887 , n19930 , n21886 );
nand ( n21888 , n21885 , n21887 );
not ( n21889 , n21888 );
not ( n21890 , n19972 );
and ( n21891 , n21889 , n21890 );
not ( n21892 , n19970 );
not ( n21893 , n21892 );
buf ( n21894 , n21893 );
and ( n21895 , n21888 , n21894 );
nor ( n21896 , n21891 , n21895 );
not ( n21897 , n21896 );
not ( n21898 , n15045 );
not ( n21899 , n13050 );
and ( n21900 , n21898 , n21899 );
and ( n21901 , n15045 , n13050 );
nor ( n21902 , n21900 , n21901 );
buf ( n21903 , n20274 );
not ( n21904 , n21903 );
and ( n21905 , n21902 , n21904 );
not ( n21906 , n21902 );
and ( n21907 , n21906 , n21903 );
nor ( n21908 , n21905 , n21907 );
not ( n21909 , n21908 );
nand ( n21910 , n21897 , n21909 );
not ( n21911 , n21910 );
xor ( n21912 , n12448 , n12457 );
xnor ( n21913 , n21912 , n12461 );
xor ( n21914 , n7237 , n21913 );
buf ( n21915 , n6273 );
buf ( n21916 , n21915 );
not ( n21917 , n21916 );
not ( n21918 , n10860 );
or ( n21919 , n21917 , n21918 );
not ( n21920 , n21915 );
nand ( n21921 , n21920 , n10855 );
nand ( n21922 , n21919 , n21921 );
not ( n21923 , n8579 );
and ( n21924 , n21922 , n21923 );
not ( n21925 , n21922 );
and ( n21926 , n21925 , n8580 );
nor ( n21927 , n21924 , n21926 );
buf ( n21928 , n6274 );
nand ( n21929 , n7197 , n21928 );
buf ( n21930 , n6275 );
buf ( n21931 , n21930 );
and ( n21932 , n21929 , n21931 );
not ( n21933 , n21929 );
not ( n21934 , n21930 );
and ( n21935 , n21933 , n21934 );
nor ( n21936 , n21932 , n21935 );
xor ( n21937 , n21927 , n21936 );
buf ( n21938 , n6276 );
nand ( n21939 , n8032 , n21938 );
buf ( n21940 , n6277 );
not ( n21941 , n21940 );
and ( n21942 , n21939 , n21941 );
not ( n21943 , n21939 );
buf ( n21944 , n21940 );
and ( n21945 , n21943 , n21944 );
nor ( n21946 , n21942 , n21945 );
xnor ( n21947 , n21937 , n21946 );
not ( n21948 , n21947 );
buf ( n21949 , n21948 );
xnor ( n21950 , n21914 , n21949 );
not ( n21951 , n21950 );
not ( n21952 , n21951 );
and ( n21953 , n21911 , n21952 );
nand ( n21954 , n21897 , n21909 );
and ( n21955 , n21954 , n21951 );
nor ( n21956 , n21953 , n21955 );
not ( n21957 , n21956 );
not ( n21958 , n9277 );
not ( n21959 , n10884 );
not ( n21960 , n9235 );
or ( n21961 , n21959 , n21960 );
or ( n21962 , n9235 , n10884 );
nand ( n21963 , n21961 , n21962 );
not ( n21964 , n21963 );
or ( n21965 , n21958 , n21964 );
not ( n21966 , n21963 );
nand ( n21967 , n21966 , n9272 );
nand ( n21968 , n21965 , n21967 );
not ( n21969 , n21968 );
not ( n21970 , n16666 );
not ( n21971 , n16250 );
or ( n21972 , n21970 , n21971 );
not ( n21973 , n16666 );
nand ( n21974 , n21973 , n11015 );
nand ( n21975 , n21972 , n21974 );
and ( n21976 , n21975 , n16257 );
not ( n21977 , n21975 );
and ( n21978 , n21977 , n16258 );
nor ( n21979 , n21976 , n21978 );
not ( n21980 , n21979 );
nand ( n21981 , n21969 , n21980 );
not ( n21982 , n12091 );
not ( n21983 , n7188 );
not ( n21984 , n21983 );
or ( n21985 , n21982 , n21984 );
not ( n21986 , n12091 );
xor ( n21987 , n7168 , n7177 );
xnor ( n21988 , n21987 , n7187 );
nand ( n21989 , n21986 , n21988 );
nand ( n21990 , n21985 , n21989 );
not ( n21991 , n14992 );
buf ( n21992 , n21991 );
and ( n21993 , n21990 , n21992 );
not ( n21994 , n21990 );
and ( n21995 , n21994 , n14997 );
nor ( n21996 , n21993 , n21995 );
buf ( n21997 , n21996 );
and ( n21998 , n21981 , n21997 );
not ( n21999 , n21981 );
not ( n22000 , n21997 );
and ( n22001 , n21999 , n22000 );
nor ( n22002 , n21998 , n22001 );
not ( n22003 , n22002 );
or ( n22004 , n21957 , n22003 );
or ( n22005 , n22002 , n21956 );
nand ( n22006 , n22004 , n22005 );
buf ( n22007 , n6278 );
buf ( n22008 , n22007 );
not ( n22009 , n22008 );
buf ( n22010 , n6279 );
not ( n22011 , n22010 );
not ( n22012 , n22011 );
or ( n22013 , n22009 , n22012 );
not ( n22014 , n22007 );
buf ( n22015 , n22010 );
nand ( n22016 , n22014 , n22015 );
nand ( n22017 , n22013 , n22016 );
and ( n22018 , n22017 , n12046 );
not ( n22019 , n22017 );
not ( n22020 , n12045 );
and ( n22021 , n22019 , n22020 );
nor ( n22022 , n22018 , n22021 );
not ( n22023 , n22022 );
buf ( n22024 , n6280 );
nand ( n22025 , n7258 , n22024 );
buf ( n22026 , n6281 );
buf ( n22027 , n22026 );
and ( n22028 , n22025 , n22027 );
not ( n22029 , n22025 );
not ( n22030 , n22026 );
and ( n22031 , n22029 , n22030 );
nor ( n22032 , n22028 , n22031 );
xor ( n22033 , n22023 , n22032 );
buf ( n22034 , n6282 );
nand ( n22035 , n7107 , n22034 );
buf ( n22036 , n6283 );
buf ( n22037 , n22036 );
and ( n22038 , n22035 , n22037 );
not ( n22039 , n22035 );
not ( n22040 , n22036 );
and ( n22041 , n22039 , n22040 );
nor ( n22042 , n22038 , n22041 );
buf ( n22043 , n22042 );
xnor ( n22044 , n22033 , n22043 );
not ( n22045 , n22044 );
not ( n22046 , n22045 );
xor ( n22047 , n7374 , n22046 );
xnor ( n22048 , n22047 , n18261 );
not ( n22049 , n22048 );
not ( n22050 , n6630 );
not ( n22051 , n10446 );
or ( n22052 , n22050 , n22051 );
nand ( n22053 , n10443 , n6627 );
nand ( n22054 , n22052 , n22053 );
and ( n22055 , n22054 , n20785 );
not ( n22056 , n22054 );
and ( n22057 , n22056 , n20778 );
nor ( n22058 , n22055 , n22057 );
not ( n22059 , n22058 );
nand ( n22060 , n22049 , n22059 );
not ( n22061 , n14640 );
not ( n22062 , n11957 );
or ( n22063 , n22061 , n22062 );
or ( n22064 , n14640 , n11956 );
nand ( n22065 , n22063 , n22064 );
buf ( n22066 , n6284 );
buf ( n22067 , n22066 );
not ( n22068 , n22067 );
buf ( n22069 , n6285 );
not ( n22070 , n22069 );
not ( n22071 , n22070 );
or ( n22072 , n22068 , n22071 );
not ( n22073 , n22066 );
buf ( n22074 , n22069 );
nand ( n22075 , n22073 , n22074 );
nand ( n22076 , n22072 , n22075 );
buf ( n22077 , n6286 );
buf ( n22078 , n22077 );
and ( n22079 , n22076 , n22078 );
not ( n22080 , n22076 );
not ( n22081 , n22077 );
and ( n22082 , n22080 , n22081 );
nor ( n22083 , n22079 , n22082 );
buf ( n22084 , n6287 );
nand ( n22085 , n8954 , n22084 );
buf ( n22086 , n6288 );
buf ( n22087 , n22086 );
and ( n22088 , n22085 , n22087 );
not ( n22089 , n22085 );
not ( n22090 , n22086 );
and ( n22091 , n22089 , n22090 );
nor ( n22092 , n22088 , n22091 );
xor ( n22093 , n22083 , n22092 );
xnor ( n22094 , n22093 , n11528 );
buf ( n22095 , n22094 );
not ( n22096 , n22095 );
not ( n22097 , n22096 );
and ( n22098 , n22065 , n22097 );
not ( n22099 , n22065 );
not ( n22100 , n22094 );
and ( n22101 , n22099 , n22100 );
nor ( n22102 , n22098 , n22101 );
not ( n22103 , n22102 );
and ( n22104 , n22060 , n22103 );
not ( n22105 , n22060 );
and ( n22106 , n22105 , n22102 );
nor ( n22107 , n22104 , n22106 );
not ( n22108 , n22107 );
and ( n22109 , n22006 , n22108 );
not ( n22110 , n22006 );
and ( n22111 , n22110 , n22107 );
nor ( n22112 , n22109 , n22111 );
not ( n22113 , n22112 );
not ( n22114 , n15207 );
not ( n22115 , n20640 );
or ( n22116 , n22114 , n22115 );
or ( n22117 , n20640 , n15207 );
nand ( n22118 , n22116 , n22117 );
not ( n22119 , n22118 );
not ( n22120 , n13254 );
and ( n22121 , n22119 , n22120 );
and ( n22122 , n22118 , n13254 );
nor ( n22123 , n22121 , n22122 );
not ( n22124 , n22123 );
not ( n22125 , n19298 );
not ( n22126 , n13918 );
not ( n22127 , n19290 );
or ( n22128 , n22126 , n22127 );
not ( n22129 , n20836 );
or ( n22130 , n22129 , n13918 );
nand ( n22131 , n22128 , n22130 );
not ( n22132 , n22131 );
or ( n22133 , n22125 , n22132 );
or ( n22134 , n22131 , n19298 );
nand ( n22135 , n22133 , n22134 );
not ( n22136 , n22135 );
nand ( n22137 , n22124 , n22136 );
not ( n22138 , n17882 );
not ( n22139 , n22138 );
not ( n22140 , n22139 );
not ( n22141 , n15261 );
buf ( n22142 , n6289 );
buf ( n22143 , n22142 );
not ( n22144 , n22143 );
buf ( n22145 , n6290 );
not ( n22146 , n22145 );
not ( n22147 , n22146 );
or ( n22148 , n22144 , n22147 );
not ( n22149 , n22142 );
buf ( n22150 , n22145 );
nand ( n22151 , n22149 , n22150 );
nand ( n22152 , n22148 , n22151 );
buf ( n22153 , n6291 );
not ( n22154 , n22153 );
and ( n22155 , n22152 , n22154 );
not ( n22156 , n22152 );
buf ( n22157 , n22153 );
and ( n22158 , n22156 , n22157 );
nor ( n22159 , n22155 , n22158 );
buf ( n22160 , n6292 );
nand ( n22161 , n8364 , n22160 );
buf ( n22162 , n6293 );
buf ( n22163 , n22162 );
and ( n22164 , n22161 , n22163 );
not ( n22165 , n22161 );
not ( n22166 , n22162 );
and ( n22167 , n22165 , n22166 );
nor ( n22168 , n22164 , n22167 );
xor ( n22169 , n22159 , n22168 );
buf ( n22170 , n6294 );
nand ( n22171 , n6502 , n22170 );
buf ( n22172 , n6295 );
buf ( n22173 , n22172 );
and ( n22174 , n22171 , n22173 );
not ( n22175 , n22171 );
not ( n22176 , n22172 );
and ( n22177 , n22175 , n22176 );
nor ( n22178 , n22174 , n22177 );
not ( n22179 , n22178 );
xnor ( n22180 , n22169 , n22179 );
not ( n22181 , n22180 );
or ( n22182 , n22141 , n22181 );
not ( n22183 , n15261 );
not ( n22184 , n22159 );
xor ( n22185 , n22184 , n22178 );
not ( n22186 , n22168 );
xnor ( n22187 , n22185 , n22186 );
nand ( n22188 , n22183 , n22187 );
nand ( n22189 , n22182 , n22188 );
not ( n22190 , n22189 );
or ( n22191 , n22140 , n22190 );
or ( n22192 , n17883 , n22189 );
nand ( n22193 , n22191 , n22192 );
not ( n22194 , n22193 );
and ( n22195 , n22137 , n22194 );
not ( n22196 , n22137 );
and ( n22197 , n22196 , n22193 );
nor ( n22198 , n22195 , n22197 );
not ( n22199 , n21861 );
nand ( n22200 , n21825 , n22199 );
not ( n22201 , n22200 );
not ( n22202 , n20487 );
not ( n22203 , n7580 );
or ( n22204 , n22202 , n22203 );
or ( n22205 , n7580 , n20487 );
nand ( n22206 , n22204 , n22205 );
not ( n22207 , n22206 );
buf ( n22208 , n6296 );
buf ( n22209 , n22208 );
not ( n22210 , n22209 );
buf ( n22211 , n6297 );
not ( n22212 , n22211 );
not ( n22213 , n22212 );
or ( n22214 , n22210 , n22213 );
not ( n22215 , n22208 );
buf ( n22216 , n22211 );
nand ( n22217 , n22215 , n22216 );
nand ( n22218 , n22214 , n22217 );
buf ( n22219 , n6298 );
not ( n22220 , n22219 );
and ( n22221 , n22218 , n22220 );
not ( n22222 , n22218 );
buf ( n22223 , n22219 );
and ( n22224 , n22222 , n22223 );
nor ( n22225 , n22221 , n22224 );
buf ( n22226 , n6299 );
nand ( n22227 , n6927 , n22226 );
buf ( n22228 , n6300 );
not ( n22229 , n22228 );
and ( n22230 , n22227 , n22229 );
not ( n22231 , n22227 );
buf ( n22232 , n22228 );
and ( n22233 , n22231 , n22232 );
nor ( n22234 , n22230 , n22233 );
xor ( n22235 , n22225 , n22234 );
buf ( n22236 , n6301 );
nand ( n22237 , n6770 , n22236 );
buf ( n22238 , n6302 );
buf ( n22239 , n22238 );
and ( n22240 , n22237 , n22239 );
not ( n22241 , n22237 );
not ( n22242 , n22238 );
and ( n22243 , n22241 , n22242 );
nor ( n22244 , n22240 , n22243 );
xor ( n22245 , n22235 , n22244 );
not ( n22246 , n22245 );
buf ( n22247 , n22246 );
not ( n22248 , n22247 );
and ( n22249 , n22207 , n22248 );
and ( n22250 , n22206 , n22247 );
nor ( n22251 , n22249 , n22250 );
not ( n22252 , n22251 );
not ( n22253 , n22252 );
and ( n22254 , n22201 , n22253 );
and ( n22255 , n22200 , n22252 );
nor ( n22256 , n22254 , n22255 );
and ( n22257 , n22198 , n22256 );
not ( n22258 , n22198 );
not ( n22259 , n22256 );
and ( n22260 , n22258 , n22259 );
nor ( n22261 , n22257 , n22260 );
not ( n22262 , n22261 );
not ( n22263 , n22262 );
and ( n22264 , n22113 , n22263 );
and ( n22265 , n22112 , n22262 );
nor ( n22266 , n22264 , n22265 );
not ( n22267 , n22266 );
or ( n22268 , n21881 , n22267 );
not ( n22269 , n21880 );
not ( n22270 , n22262 );
not ( n22271 , n22112 );
or ( n22272 , n22270 , n22271 );
not ( n22273 , n22112 );
nand ( n22274 , n22273 , n22261 );
nand ( n22275 , n22272 , n22274 );
nand ( n22276 , n22269 , n22275 );
nand ( n22277 , n22268 , n22276 );
not ( n22278 , n6574 );
not ( n22279 , n13086 );
not ( n22280 , n22279 );
not ( n22281 , n15052 );
or ( n22282 , n22280 , n22281 );
or ( n22283 , n15052 , n22279 );
nand ( n22284 , n22282 , n22283 );
and ( n22285 , n22284 , n21904 );
not ( n22286 , n22284 );
not ( n22287 , n20274 );
not ( n22288 , n22287 );
and ( n22289 , n22286 , n22288 );
nor ( n22290 , n22285 , n22289 );
not ( n22291 , n22290 );
nand ( n22292 , n22291 , n6664 );
not ( n22293 , n22292 );
or ( n22294 , n22278 , n22293 );
not ( n22295 , n22290 );
nand ( n22296 , n22295 , n6664 );
or ( n22297 , n22296 , n6574 );
nand ( n22298 , n22294 , n22297 );
not ( n22299 , n14445 );
not ( n22300 , n8186 );
or ( n22301 , n22299 , n22300 );
not ( n22302 , n14445 );
nand ( n22303 , n22302 , n8192 );
nand ( n22304 , n22301 , n22303 );
not ( n22305 , n8234 );
and ( n22306 , n22304 , n22305 );
not ( n22307 , n22304 );
and ( n22308 , n22307 , n8233 );
nor ( n22309 , n22306 , n22308 );
not ( n22310 , n9598 );
not ( n22311 , n22310 );
buf ( n22312 , n9929 );
and ( n22313 , n22312 , n21853 );
not ( n22314 , n22312 );
and ( n22315 , n22314 , n21854 );
or ( n22316 , n22313 , n22315 );
not ( n22317 , n22316 );
not ( n22318 , n22317 );
or ( n22319 , n22311 , n22318 );
nand ( n22320 , n22316 , n9598 );
nand ( n22321 , n22319 , n22320 );
nand ( n22322 , n22309 , n22321 );
and ( n22323 , n22322 , n7320 );
not ( n22324 , n22322 );
and ( n22325 , n22324 , n7321 );
nor ( n22326 , n22323 , n22325 );
and ( n22327 , n22298 , n22326 );
not ( n22328 , n22298 );
not ( n22329 , n22326 );
and ( n22330 , n22328 , n22329 );
nor ( n22331 , n22327 , n22330 );
not ( n22332 , n22331 );
not ( n22333 , n8745 );
not ( n22334 , n22333 );
buf ( n22335 , n6303 );
buf ( n22336 , n22335 );
buf ( n22337 , n6304 );
buf ( n22338 , n22337 );
not ( n22339 , n22338 );
buf ( n22340 , n6305 );
not ( n22341 , n22340 );
not ( n22342 , n22341 );
or ( n22343 , n22339 , n22342 );
not ( n22344 , n22337 );
buf ( n22345 , n22340 );
nand ( n22346 , n22344 , n22345 );
nand ( n22347 , n22343 , n22346 );
buf ( n22348 , n22347 );
xor ( n22349 , n22336 , n22348 );
buf ( n22350 , n6306 );
nand ( n22351 , n10372 , n22350 );
buf ( n22352 , n6307 );
not ( n22353 , n22352 );
and ( n22354 , n22351 , n22353 );
not ( n22355 , n22351 );
buf ( n22356 , n22352 );
and ( n22357 , n22355 , n22356 );
nor ( n22358 , n22354 , n22357 );
not ( n22359 , n22358 );
not ( n22360 , n22359 );
buf ( n22361 , n6308 );
nand ( n22362 , n10372 , n22361 );
buf ( n22363 , n6309 );
buf ( n22364 , n22363 );
and ( n22365 , n22362 , n22364 );
not ( n22366 , n22362 );
not ( n22367 , n22363 );
and ( n22368 , n22366 , n22367 );
nor ( n22369 , n22365 , n22368 );
not ( n22370 , n22369 );
not ( n22371 , n22370 );
or ( n22372 , n22360 , n22371 );
nand ( n22373 , n22369 , n22358 );
nand ( n22374 , n22372 , n22373 );
xnor ( n22375 , n22349 , n22374 );
not ( n22376 , n22375 );
or ( n22377 , n22334 , n22376 );
not ( n22378 , n22335 );
xor ( n22379 , n22378 , n22347 );
xor ( n22380 , n22379 , n22374 );
or ( n22381 , n22380 , n22333 );
nand ( n22382 , n22377 , n22381 );
and ( n22383 , n22382 , n10851 );
not ( n22384 , n22382 );
not ( n22385 , n10851 );
and ( n22386 , n22384 , n22385 );
nor ( n22387 , n22383 , n22386 );
not ( n22388 , n10959 );
not ( n22389 , n18322 );
not ( n22390 , n10916 );
not ( n22391 , n22390 );
or ( n22392 , n22389 , n22391 );
not ( n22393 , n18322 );
nand ( n22394 , n22393 , n10916 );
nand ( n22395 , n22392 , n22394 );
not ( n22396 , n22395 );
or ( n22397 , n22388 , n22396 );
or ( n22398 , n22395 , n10959 );
nand ( n22399 , n22397 , n22398 );
nand ( n22400 , n22387 , n22399 );
not ( n22401 , n22400 );
not ( n22402 , n6951 );
and ( n22403 , n22401 , n22402 );
and ( n22404 , n22400 , n6951 );
nor ( n22405 , n22403 , n22404 );
not ( n22406 , n22405 );
or ( n22407 , n22332 , n22406 );
or ( n22408 , n22331 , n22405 );
nand ( n22409 , n22407 , n22408 );
not ( n22410 , n7837 );
not ( n22411 , n13784 );
buf ( n22412 , n19576 );
xor ( n22413 , n22412 , n19586 );
xnor ( n22414 , n22413 , n19593 );
not ( n22415 , n22414 );
not ( n22416 , n22415 );
or ( n22417 , n22411 , n22416 );
not ( n22418 , n13784 );
nand ( n22419 , n22418 , n22414 );
nand ( n22420 , n22417 , n22419 );
and ( n22421 , n22420 , n19608 );
not ( n22422 , n22420 );
and ( n22423 , n22422 , n19605 );
nor ( n22424 , n22421 , n22423 );
buf ( n22425 , n16003 );
not ( n22426 , n22425 );
buf ( n22427 , n6310 );
buf ( n22428 , n22427 );
not ( n22429 , n22428 );
buf ( n22430 , n6311 );
not ( n22431 , n22430 );
not ( n22432 , n22431 );
or ( n22433 , n22429 , n22432 );
not ( n22434 , n22427 );
buf ( n22435 , n22430 );
nand ( n22436 , n22434 , n22435 );
nand ( n22437 , n22433 , n22436 );
buf ( n22438 , n6312 );
not ( n22439 , n22438 );
and ( n22440 , n22437 , n22439 );
not ( n22441 , n22437 );
buf ( n22442 , n22438 );
and ( n22443 , n22441 , n22442 );
nor ( n22444 , n22440 , n22443 );
buf ( n22445 , n6313 );
nand ( n22446 , n7977 , n22445 );
buf ( n22447 , n6314 );
not ( n22448 , n22447 );
and ( n22449 , n22446 , n22448 );
not ( n22450 , n22446 );
buf ( n22451 , n22447 );
and ( n22452 , n22450 , n22451 );
nor ( n22453 , n22449 , n22452 );
xor ( n22454 , n22444 , n22453 );
buf ( n22455 , n6315 );
nand ( n22456 , n8032 , n22455 );
buf ( n22457 , n6316 );
buf ( n22458 , n22457 );
and ( n22459 , n22456 , n22458 );
not ( n22460 , n22456 );
not ( n22461 , n22457 );
and ( n22462 , n22460 , n22461 );
nor ( n22463 , n22459 , n22462 );
xor ( n22464 , n22454 , n22463 );
buf ( n22465 , n22464 );
not ( n22466 , n22465 );
not ( n22467 , n22466 );
or ( n22468 , n22426 , n22467 );
not ( n22469 , n22466 );
not ( n22470 , n22425 );
nand ( n22471 , n22469 , n22470 );
nand ( n22472 , n22468 , n22471 );
buf ( n22473 , n18208 );
and ( n22474 , n22472 , n22473 );
not ( n22475 , n22472 );
buf ( n22476 , n18207 );
and ( n22477 , n22475 , n22476 );
nor ( n22478 , n22474 , n22477 );
nand ( n22479 , n22424 , n22478 );
not ( n22480 , n22479 );
and ( n22481 , n22410 , n22480 );
and ( n22482 , n7837 , n22479 );
nor ( n22483 , n22481 , n22482 );
not ( n22484 , n22483 );
not ( n22485 , n22484 );
buf ( n22486 , n6643 );
and ( n22487 , n22486 , n10443 );
not ( n22488 , n22486 );
and ( n22489 , n22488 , n10446 );
nor ( n22490 , n22487 , n22489 );
not ( n22491 , n20784 );
and ( n22492 , n22490 , n22491 );
not ( n22493 , n22490 );
and ( n22494 , n22493 , n20778 );
nor ( n22495 , n22492 , n22494 );
not ( n22496 , n22495 );
not ( n22497 , n13988 );
not ( n22498 , n20828 );
or ( n22499 , n22497 , n22498 );
or ( n22500 , n21396 , n13988 );
nand ( n22501 , n22499 , n22500 );
and ( n22502 , n22501 , n19290 );
not ( n22503 , n22501 );
and ( n22504 , n22503 , n19293 );
nor ( n22505 , n22502 , n22504 );
not ( n22506 , n22505 );
nand ( n22507 , n22496 , n22506 );
not ( n22508 , n22507 );
not ( n22509 , n7497 );
or ( n22510 , n22508 , n22509 );
or ( n22511 , n7497 , n22507 );
nand ( n22512 , n22510 , n22511 );
not ( n22513 , n22512 );
not ( n22514 , n22513 );
or ( n22515 , n22485 , n22514 );
nand ( n22516 , n22483 , n22512 );
nand ( n22517 , n22515 , n22516 );
and ( n22518 , n22409 , n22517 );
not ( n22519 , n22409 );
not ( n22520 , n22517 );
and ( n22521 , n22519 , n22520 );
nor ( n22522 , n22518 , n22521 );
buf ( n22523 , n22522 );
and ( n22524 , n22277 , n22523 );
not ( n22525 , n22277 );
and ( n22526 , n22409 , n22520 );
not ( n22527 , n22409 );
and ( n22528 , n22527 , n22517 );
nor ( n22529 , n22526 , n22528 );
buf ( n22530 , n22529 );
and ( n22531 , n22525 , n22530 );
nor ( n22532 , n22524 , n22531 );
not ( n22533 , n22532 );
nand ( n22534 , n21822 , n22533 );
xor ( n22535 , n11529 , n11536 );
xnor ( n22536 , n22535 , n11543 );
buf ( n22537 , n22536 );
not ( n22538 , n22537 );
not ( n22539 , n22538 );
not ( n22540 , n22078 );
and ( n22541 , n22539 , n22540 );
not ( n22542 , n22537 );
and ( n22543 , n22542 , n22078 );
nor ( n22544 , n22541 , n22543 );
buf ( n22545 , n11575 );
and ( n22546 , n22544 , n22545 );
not ( n22547 , n22544 );
xor ( n22548 , n11563 , n11573 );
xor ( n22549 , n22548 , n11455 );
buf ( n22550 , n22549 );
and ( n22551 , n22547 , n22550 );
nor ( n22552 , n22546 , n22551 );
not ( n22553 , n10838 );
buf ( n22554 , n21447 );
not ( n22555 , n22554 );
or ( n22556 , n22553 , n22555 );
not ( n22557 , n21699 );
not ( n22558 , n22557 );
nand ( n22559 , n22558 , n10834 );
nand ( n22560 , n22556 , n22559 );
and ( n22561 , n22560 , n21453 );
not ( n22562 , n22560 );
buf ( n22563 , n18710 );
and ( n22564 , n22562 , n22563 );
nor ( n22565 , n22561 , n22564 );
nand ( n22566 , n22552 , n22565 );
not ( n22567 , n11407 );
not ( n22568 , n6792 );
or ( n22569 , n22567 , n22568 );
or ( n22570 , n6791 , n11407 );
nand ( n22571 , n22569 , n22570 );
and ( n22572 , n22571 , n20464 );
not ( n22573 , n22571 );
and ( n22574 , n22573 , n20463 );
nor ( n22575 , n22572 , n22574 );
and ( n22576 , n22566 , n22575 );
not ( n22577 , n22566 );
not ( n22578 , n22575 );
and ( n22579 , n22577 , n22578 );
nor ( n22580 , n22576 , n22579 );
not ( n22581 , n22580 );
and ( n22582 , n10442 , n6656 );
not ( n22583 , n10442 );
and ( n22584 , n22583 , n6657 );
or ( n22585 , n22582 , n22584 );
not ( n22586 , n20783 );
and ( n22587 , n22585 , n22586 );
not ( n22588 , n22585 );
and ( n22589 , n22588 , n20778 );
nor ( n22590 , n22587 , n22589 );
not ( n22591 , n22590 );
not ( n22592 , n22591 );
not ( n22593 , n16408 );
buf ( n22594 , n6317 );
not ( n22595 , n22594 );
and ( n22596 , n22593 , n22595 );
and ( n22597 , n16408 , n22594 );
nor ( n22598 , n22596 , n22597 );
not ( n22599 , n22598 );
not ( n22600 , n16229 );
or ( n22601 , n22599 , n22600 );
or ( n22602 , n16229 , n22598 );
nand ( n22603 , n22601 , n22602 );
not ( n22604 , n11317 );
xor ( n22605 , n17657 , n17661 );
xnor ( n22606 , n22605 , n17671 );
not ( n22607 , n22606 );
or ( n22608 , n22604 , n22607 );
or ( n22609 , n22606 , n11317 );
nand ( n22610 , n22608 , n22609 );
and ( n22611 , n22610 , n17332 );
not ( n22612 , n22610 );
and ( n22613 , n22612 , n17347 );
nor ( n22614 , n22611 , n22613 );
nand ( n22615 , n22603 , n22614 );
not ( n22616 , n22615 );
or ( n22617 , n22592 , n22616 );
or ( n22618 , n22615 , n22591 );
nand ( n22619 , n22617 , n22618 );
not ( n22620 , n22619 );
not ( n22621 , n13368 );
not ( n22622 , n19322 );
not ( n22623 , n22622 );
or ( n22624 , n22621 , n22623 );
not ( n22625 , n13368 );
nand ( n22626 , n22625 , n19322 );
nand ( n22627 , n22624 , n22626 );
buf ( n22628 , n6318 );
buf ( n22629 , n22628 );
not ( n22630 , n22629 );
not ( n22631 , n14226 );
or ( n22632 , n22630 , n22631 );
not ( n22633 , n22628 );
nand ( n22634 , n22633 , n14180 );
nand ( n22635 , n22632 , n22634 );
buf ( n22636 , n6319 );
not ( n22637 , n22636 );
and ( n22638 , n22635 , n22637 );
not ( n22639 , n22635 );
buf ( n22640 , n22636 );
and ( n22641 , n22639 , n22640 );
nor ( n22642 , n22638 , n22641 );
buf ( n22643 , n6320 );
nand ( n22644 , n7698 , n22643 );
buf ( n22645 , n6321 );
xor ( n22646 , n22644 , n22645 );
xor ( n22647 , n22642 , n22646 );
buf ( n22648 , n6322 );
nand ( n22649 , n10383 , n22648 );
buf ( n22650 , n6323 );
not ( n22651 , n22650 );
and ( n22652 , n22649 , n22651 );
not ( n22653 , n22649 );
buf ( n22654 , n22650 );
and ( n22655 , n22653 , n22654 );
nor ( n22656 , n22652 , n22655 );
xnor ( n22657 , n22647 , n22656 );
buf ( n22658 , n22657 );
xor ( n22659 , n22627 , n22658 );
not ( n22660 , n7270 );
buf ( n22661 , n8301 );
not ( n22662 , n22661 );
and ( n22663 , n22660 , n22662 );
and ( n22664 , n7270 , n22661 );
nor ( n22665 , n22663 , n22664 );
and ( n22666 , n22665 , n7315 );
not ( n22667 , n22665 );
and ( n22668 , n22667 , n9001 );
nor ( n22669 , n22666 , n22668 );
nand ( n22670 , n22659 , n22669 );
not ( n22671 , n22670 );
not ( n22672 , n7191 );
not ( n22673 , n19442 );
or ( n22674 , n22672 , n22673 );
not ( n22675 , n7191 );
nand ( n22676 , n22675 , n19446 );
nand ( n22677 , n22674 , n22676 );
and ( n22678 , n22677 , n18863 );
not ( n22679 , n22677 );
not ( n22680 , n18863 );
and ( n22681 , n22679 , n22680 );
nor ( n22682 , n22678 , n22681 );
not ( n22683 , n22682 );
and ( n22684 , n22671 , n22683 );
nand ( n22685 , n22659 , n22669 );
and ( n22686 , n22685 , n22682 );
nor ( n22687 , n22684 , n22686 );
not ( n22688 , n22687 );
or ( n22689 , n22620 , n22688 );
or ( n22690 , n22687 , n22619 );
nand ( n22691 , n22689 , n22690 );
buf ( n22692 , n6324 );
xor ( n22693 , n22692 , n18300 );
not ( n22694 , n12907 );
xnor ( n22695 , n22693 , n22694 );
not ( n22696 , n22695 );
xor ( n22697 , n11072 , n13133 );
xor ( n22698 , n13182 , n13146 );
xnor ( n22699 , n22698 , n13177 );
buf ( n22700 , n22699 );
xnor ( n22701 , n22697 , n22700 );
nand ( n22702 , n22696 , n22701 );
and ( n22703 , n9308 , n21491 );
not ( n22704 , n9308 );
buf ( n22705 , n16658 );
and ( n22706 , n22704 , n22705 );
or ( n22707 , n22703 , n22706 );
not ( n22708 , n16685 );
and ( n22709 , n22707 , n22708 );
not ( n22710 , n22707 );
and ( n22711 , n22710 , n16685 );
nor ( n22712 , n22709 , n22711 );
and ( n22713 , n22702 , n22712 );
not ( n22714 , n22702 );
not ( n22715 , n22712 );
and ( n22716 , n22714 , n22715 );
nor ( n22717 , n22713 , n22716 );
xor ( n22718 , n22691 , n22717 );
not ( n22719 , n22565 );
nand ( n22720 , n22575 , n22719 );
not ( n22721 , n8762 );
buf ( n22722 , n6325 );
nand ( n22723 , n6828 , n22722 );
buf ( n22724 , n6326 );
not ( n22725 , n22724 );
and ( n22726 , n22723 , n22725 );
not ( n22727 , n22723 );
buf ( n22728 , n22724 );
and ( n22729 , n22727 , n22728 );
nor ( n22730 , n22726 , n22729 );
buf ( n22731 , n22730 );
not ( n22732 , n22731 );
not ( n22733 , n18082 );
nor ( n22734 , n22732 , n22733 );
not ( n22735 , n22734 );
not ( n22736 , n22731 );
nand ( n22737 , n22736 , n20428 );
nand ( n22738 , n22735 , n22737 );
not ( n22739 , n22738 );
and ( n22740 , n22721 , n22739 );
not ( n22741 , n8761 );
and ( n22742 , n22741 , n22738 );
nor ( n22743 , n22740 , n22742 );
and ( n22744 , n22720 , n22743 );
not ( n22745 , n22720 );
not ( n22746 , n22743 );
and ( n22747 , n22745 , n22746 );
nor ( n22748 , n22744 , n22747 );
not ( n22749 , n22748 );
not ( n22750 , n15069 );
not ( n22751 , n14508 );
not ( n22752 , n22751 );
or ( n22753 , n22750 , n22752 );
nand ( n22754 , n14508 , n15065 );
nand ( n22755 , n22753 , n22754 );
not ( n22756 , n16898 );
not ( n22757 , n22756 );
and ( n22758 , n22755 , n22757 );
not ( n22759 , n22755 );
and ( n22760 , n22759 , n22756 );
nor ( n22761 , n22758 , n22760 );
not ( n22762 , n13561 );
not ( n22763 , n19243 );
or ( n22764 , n22762 , n22763 );
not ( n22765 , n11228 );
nand ( n22766 , n22765 , n13557 );
nand ( n22767 , n22764 , n22766 );
and ( n22768 , n22767 , n11272 );
not ( n22769 , n22767 );
and ( n22770 , n22769 , n11275 );
nor ( n22771 , n22768 , n22770 );
not ( n22772 , n22771 );
nand ( n22773 , n22761 , n22772 );
not ( n22774 , n22773 );
buf ( n22775 , n10381 );
xor ( n22776 , n22775 , n12149 );
xnor ( n22777 , n22776 , n7829 );
not ( n22778 , n22777 );
and ( n22779 , n22774 , n22778 );
and ( n22780 , n22773 , n22777 );
nor ( n22781 , n22779 , n22780 );
not ( n22782 , n22781 );
or ( n22783 , n22749 , n22782 );
or ( n22784 , n22781 , n22748 );
nand ( n22785 , n22783 , n22784 );
not ( n22786 , n22785 );
and ( n22787 , n22718 , n22786 );
not ( n22788 , n22718 );
and ( n22789 , n22788 , n22785 );
nor ( n22790 , n22787 , n22789 );
not ( n22791 , n22790 );
not ( n22792 , n22791 );
not ( n22793 , n22792 );
or ( n22794 , n22581 , n22793 );
not ( n22795 , n22580 );
nand ( n22796 , n22795 , n22791 );
nand ( n22797 , n22794 , n22796 );
not ( n22798 , n6490 );
not ( n22799 , n15639 );
not ( n22800 , n22799 );
or ( n22801 , n22798 , n22800 );
buf ( n22802 , n15634 );
not ( n22803 , n22802 );
or ( n22804 , n22803 , n6490 );
nand ( n22805 , n22801 , n22804 );
not ( n22806 , n15603 );
not ( n22807 , n22806 );
and ( n22808 , n22805 , n22807 );
not ( n22809 , n22805 );
and ( n22810 , n22809 , n15604 );
nor ( n22811 , n22808 , n22810 );
not ( n22812 , n10120 );
not ( n22813 , n15474 );
or ( n22814 , n22812 , n22813 );
or ( n22815 , n15474 , n10120 );
nand ( n22816 , n22814 , n22815 );
buf ( n22817 , n12707 );
and ( n22818 , n22816 , n22817 );
not ( n22819 , n22816 );
not ( n22820 , n12713 );
not ( n22821 , n22820 );
and ( n22822 , n22819 , n22821 );
nor ( n22823 , n22818 , n22822 );
not ( n22824 , n22823 );
nand ( n22825 , n22811 , n22824 );
not ( n22826 , n22825 );
not ( n22827 , n14656 );
not ( n22828 , n19604 );
or ( n22829 , n22827 , n22828 );
or ( n22830 , n19605 , n14656 );
nand ( n22831 , n22829 , n22830 );
and ( n22832 , n22831 , n11957 );
not ( n22833 , n22831 );
and ( n22834 , n22833 , n11958 );
nor ( n22835 , n22832 , n22834 );
not ( n22836 , n22835 );
not ( n22837 , n22836 );
and ( n22838 , n22826 , n22837 );
and ( n22839 , n22825 , n22836 );
nor ( n22840 , n22838 , n22839 );
not ( n22841 , n22840 );
buf ( n22842 , n22044 );
xor ( n22843 , n7388 , n22842 );
xnor ( n22844 , n22843 , n18261 );
not ( n22845 , n22844 );
not ( n22846 , n21249 );
xor ( n22847 , n21133 , n21143 );
xor ( n22848 , n22847 , n16299 );
not ( n22849 , n22848 );
or ( n22850 , n22846 , n22849 );
or ( n22851 , n21149 , n21249 );
nand ( n22852 , n22850 , n22851 );
and ( n22853 , n22852 , n22180 );
not ( n22854 , n22852 );
and ( n22855 , n22854 , n22187 );
nor ( n22856 , n22853 , n22855 );
not ( n22857 , n22856 );
nand ( n22858 , n22845 , n22857 );
not ( n22859 , n7970 );
not ( n22860 , n14541 );
not ( n22861 , n22860 );
or ( n22862 , n22859 , n22861 );
not ( n22863 , n14541 );
not ( n22864 , n22863 );
nand ( n22865 , n22864 , n7966 );
nand ( n22866 , n22862 , n22865 );
buf ( n22867 , n22751 );
and ( n22868 , n22866 , n22867 );
not ( n22869 , n22866 );
and ( n22870 , n22869 , n14508 );
nor ( n22871 , n22868 , n22870 );
and ( n22872 , n22858 , n22871 );
not ( n22873 , n22858 );
not ( n22874 , n22871 );
and ( n22875 , n22873 , n22874 );
nor ( n22876 , n22872 , n22875 );
not ( n22877 , n22876 );
or ( n22878 , n22841 , n22877 );
or ( n22879 , n22876 , n22840 );
nand ( n22880 , n22878 , n22879 );
not ( n22881 , n22880 );
not ( n22882 , n22881 );
not ( n22883 , n13398 );
not ( n22884 , n16316 );
and ( n22885 , n22883 , n22884 );
and ( n22886 , n13398 , n16316 );
nor ( n22887 , n22885 , n22886 );
not ( n22888 , n7627 );
not ( n22889 , n22888 );
and ( n22890 , n22887 , n22889 );
not ( n22891 , n22887 );
and ( n22892 , n22891 , n19552 );
nor ( n22893 , n22890 , n22892 );
not ( n22894 , n22893 );
buf ( n22895 , n9224 );
not ( n22896 , n22895 );
not ( n22897 , n9033 );
not ( n22898 , n9043 );
or ( n22899 , n22897 , n22898 );
or ( n22900 , n9033 , n9043 );
nand ( n22901 , n22899 , n22900 );
not ( n22902 , n9024 );
and ( n22903 , n22901 , n22902 );
not ( n22904 , n22901 );
and ( n22905 , n22904 , n9024 );
nor ( n22906 , n22903 , n22905 );
not ( n22907 , n22906 );
or ( n22908 , n22896 , n22907 );
not ( n22909 , n22895 );
nand ( n22910 , n22909 , n9045 );
nand ( n22911 , n22908 , n22910 );
not ( n22912 , n22911 );
not ( n22913 , n17717 );
and ( n22914 , n22912 , n22913 );
and ( n22915 , n22911 , n17717 );
nor ( n22916 , n22914 , n22915 );
not ( n22917 , n22916 );
nand ( n22918 , n22894 , n22917 );
not ( n22919 , n22918 );
buf ( n22920 , n6327 );
buf ( n22921 , n22920 );
not ( n22922 , n22921 );
buf ( n22923 , n6328 );
buf ( n22924 , n22923 );
not ( n22925 , n22924 );
not ( n22926 , n20698 );
or ( n22927 , n22925 , n22926 );
not ( n22928 , n22923 );
nand ( n22929 , n22928 , n20693 );
nand ( n22930 , n22927 , n22929 );
xor ( n22931 , n18562 , n22930 );
buf ( n22932 , n6329 );
buf ( n22933 , n6330 );
xor ( n22934 , n22932 , n22933 );
buf ( n22935 , n6331 );
nand ( n22936 , n8223 , n22935 );
xnor ( n22937 , n22934 , n22936 );
xnor ( n22938 , n22931 , n22937 );
not ( n22939 , n22938 );
or ( n22940 , n22922 , n22939 );
or ( n22941 , n22938 , n22921 );
nand ( n22942 , n22940 , n22941 );
buf ( n22943 , n17672 );
xnor ( n22944 , n22942 , n22943 );
not ( n22945 , n22944 );
and ( n22946 , n22919 , n22945 );
not ( n22947 , n22893 );
nand ( n22948 , n22947 , n22917 );
and ( n22949 , n22948 , n22944 );
nor ( n22950 , n22946 , n22949 );
not ( n22951 , n22950 );
not ( n22952 , n22951 );
not ( n22953 , n11104 );
not ( n22954 , n8134 );
and ( n22955 , n22953 , n22954 );
and ( n22956 , n11104 , n8134 );
nor ( n22957 , n22955 , n22956 );
xor ( n22958 , n21260 , n21230 );
xnor ( n22959 , n22958 , n21255 );
and ( n22960 , n22957 , n22959 );
not ( n22961 , n22957 );
and ( n22962 , n22961 , n21268 );
nor ( n22963 , n22960 , n22962 );
not ( n22964 , n19577 );
not ( n22965 , n21622 );
or ( n22966 , n22964 , n22965 );
or ( n22967 , n21622 , n19577 );
nand ( n22968 , n22966 , n22967 );
not ( n22969 , n21632 );
and ( n22970 , n22968 , n22969 );
not ( n22971 , n22968 );
and ( n22972 , n22971 , n21628 );
nor ( n22973 , n22970 , n22972 );
not ( n22974 , n22973 );
nand ( n22975 , n22963 , n22974 );
buf ( n22976 , n6332 );
not ( n22977 , n22976 );
buf ( n22978 , n6333 );
not ( n22979 , n22978 );
buf ( n22980 , n6334 );
buf ( n22981 , n22980 );
nand ( n22982 , n22979 , n22981 );
not ( n22983 , n22980 );
buf ( n22984 , n22978 );
nand ( n22985 , n22983 , n22984 );
and ( n22986 , n22982 , n22985 );
xor ( n22987 , n22977 , n22986 );
buf ( n22988 , n6335 );
buf ( n22989 , n6336 );
xor ( n22990 , n22988 , n22989 );
buf ( n22991 , n6337 );
nand ( n22992 , n7259 , n22991 );
xnor ( n22993 , n22990 , n22992 );
xnor ( n22994 , n22987 , n22993 );
not ( n22995 , n22994 );
not ( n22996 , n14956 );
not ( n22997 , n18821 );
or ( n22998 , n22996 , n22997 );
or ( n22999 , n18821 , n14956 );
nand ( n23000 , n22998 , n22999 );
not ( n23001 , n23000 );
and ( n23002 , n22995 , n23001 );
buf ( n23003 , n22994 );
and ( n23004 , n23003 , n23000 );
nor ( n23005 , n23002 , n23004 );
and ( n23006 , n22975 , n23005 );
not ( n23007 , n22975 );
not ( n23008 , n23005 );
and ( n23009 , n23007 , n23008 );
nor ( n23010 , n23006 , n23009 );
not ( n23011 , n23010 );
not ( n23012 , n23011 );
or ( n23013 , n22952 , n23012 );
nand ( n23014 , n22950 , n23010 );
nand ( n23015 , n23013 , n23014 );
xor ( n23016 , n14813 , n7494 );
xor ( n23017 , n23016 , n10912 );
not ( n23018 , n23017 );
not ( n23019 , n16539 );
not ( n23020 , n17769 );
or ( n23021 , n23019 , n23020 );
nand ( n23022 , n17772 , n16538 );
nand ( n23023 , n23021 , n23022 );
not ( n23024 , n23023 );
not ( n23025 , n17776 );
and ( n23026 , n23024 , n23025 );
and ( n23027 , n17776 , n23023 );
nor ( n23028 , n23026 , n23027 );
not ( n23029 , n23028 );
nand ( n23030 , n23018 , n23029 );
not ( n23031 , n21916 );
not ( n23032 , n8619 );
or ( n23033 , n23031 , n23032 );
not ( n23034 , n8618 );
not ( n23035 , n23034 );
or ( n23036 , n23035 , n21916 );
nand ( n23037 , n23033 , n23036 );
and ( n23038 , n23037 , n8662 );
not ( n23039 , n23037 );
and ( n23040 , n23039 , n8663 );
nor ( n23041 , n23038 , n23040 );
not ( n23042 , n23041 );
and ( n23043 , n23030 , n23042 );
not ( n23044 , n23030 );
and ( n23045 , n23044 , n23041 );
nor ( n23046 , n23043 , n23045 );
and ( n23047 , n23015 , n23046 );
not ( n23048 , n23015 );
not ( n23049 , n23046 );
and ( n23050 , n23048 , n23049 );
nor ( n23051 , n23047 , n23050 );
not ( n23052 , n23051 );
or ( n23053 , n22882 , n23052 );
or ( n23054 , n23051 , n22881 );
nand ( n23055 , n23053 , n23054 );
not ( n23056 , n23055 );
not ( n23057 , n23056 );
not ( n23058 , n23057 );
and ( n23059 , n22797 , n23058 );
not ( n23060 , n22797 );
and ( n23061 , n23060 , n23057 );
nor ( n23062 , n23059 , n23061 );
not ( n23063 , n23062 );
and ( n23064 , n22534 , n23063 );
not ( n23065 , n22534 );
and ( n23066 , n23065 , n23062 );
nor ( n23067 , n23064 , n23066 );
not ( n23068 , n21737 );
buf ( n23069 , n23068 );
or ( n23070 , n23067 , n23069 );
nand ( n23071 , n21746 , n23070 );
buf ( n23072 , n23071 );
buf ( n23073 , n23072 );
not ( n23074 , n12370 );
not ( n23075 , n10541 );
or ( n23076 , n23074 , n23075 );
not ( n23077 , n12370 );
nand ( n23078 , n23077 , n10534 );
nand ( n23079 , n23076 , n23078 );
and ( n23080 , n23079 , n10587 );
not ( n23081 , n23079 );
and ( n23082 , n23081 , n10581 );
nor ( n23083 , n23080 , n23082 );
not ( n23084 , n23083 );
and ( n23085 , n6533 , n15603 );
not ( n23086 , n6533 );
and ( n23087 , n23086 , n15602 );
nor ( n23088 , n23085 , n23087 );
buf ( n23089 , n6338 );
buf ( n23090 , n6339 );
nand ( n23091 , n8537 , n23090 );
buf ( n23092 , n6340 );
buf ( n23093 , n23092 );
and ( n23094 , n23091 , n23093 );
not ( n23095 , n23091 );
not ( n23096 , n23092 );
and ( n23097 , n23095 , n23096 );
nor ( n23098 , n23094 , n23097 );
xor ( n23099 , n23089 , n23098 );
buf ( n23100 , n6341 );
nand ( n23101 , n6647 , n23100 );
buf ( n23102 , n6342 );
not ( n23103 , n23102 );
and ( n23104 , n23101 , n23103 );
not ( n23105 , n23101 );
buf ( n23106 , n23102 );
and ( n23107 , n23105 , n23106 );
nor ( n23108 , n23104 , n23107 );
xnor ( n23109 , n23099 , n23108 );
not ( n23110 , n23109 );
buf ( n23111 , n6343 );
buf ( n23112 , n23111 );
not ( n23113 , n23112 );
buf ( n23114 , n6344 );
not ( n23115 , n23114 );
not ( n23116 , n23115 );
or ( n23117 , n23113 , n23116 );
not ( n23118 , n23111 );
buf ( n23119 , n23114 );
nand ( n23120 , n23118 , n23119 );
nand ( n23121 , n23117 , n23120 );
not ( n23122 , n23121 );
not ( n23123 , n23122 );
and ( n23124 , n23110 , n23123 );
and ( n23125 , n23109 , n23122 );
nor ( n23126 , n23124 , n23125 );
and ( n23127 , n23088 , n23126 );
not ( n23128 , n23088 );
not ( n23129 , n23126 );
and ( n23130 , n23128 , n23129 );
nor ( n23131 , n23127 , n23130 );
nand ( n23132 , n23084 , n23131 );
not ( n23133 , n23132 );
buf ( n23134 , n6345 );
nand ( n23135 , n13581 , n23134 );
buf ( n23136 , n6346 );
not ( n23137 , n23136 );
and ( n23138 , n23135 , n23137 );
not ( n23139 , n23135 );
buf ( n23140 , n23136 );
and ( n23141 , n23139 , n23140 );
nor ( n23142 , n23138 , n23141 );
buf ( n23143 , n23142 );
not ( n23144 , n23143 );
not ( n23145 , n13502 );
or ( n23146 , n23144 , n23145 );
not ( n23147 , n23143 );
not ( n23148 , n13490 );
not ( n23149 , n13500 );
or ( n23150 , n23148 , n23149 );
or ( n23151 , n13490 , n13500 );
nand ( n23152 , n23150 , n23151 );
xnor ( n23153 , n23152 , n13481 );
nand ( n23154 , n23147 , n23153 );
nand ( n23155 , n23146 , n23154 );
and ( n23156 , n23155 , n13516 );
not ( n23157 , n23155 );
and ( n23158 , n23157 , n7224 );
nor ( n23159 , n23156 , n23158 );
not ( n23160 , n23159 );
and ( n23161 , n23133 , n23160 );
not ( n23162 , n23083 );
nand ( n23163 , n23162 , n23131 );
and ( n23164 , n23163 , n23159 );
nor ( n23165 , n23161 , n23164 );
not ( n23166 , n23165 );
not ( n23167 , n23166 );
not ( n23168 , n23159 );
nand ( n23169 , n23168 , n23083 );
not ( n23170 , n18347 );
not ( n23171 , n20496 );
xor ( n23172 , n23171 , n20515 );
not ( n23173 , n20505 );
xnor ( n23174 , n23172 , n23173 );
not ( n23175 , n23174 );
or ( n23176 , n23170 , n23175 );
nand ( n23177 , n20517 , n18350 );
nand ( n23178 , n23176 , n23177 );
not ( n23179 , n23178 );
buf ( n23180 , n20037 );
not ( n23181 , n23180 );
and ( n23182 , n23179 , n23181 );
and ( n23183 , n23178 , n23180 );
nor ( n23184 , n23182 , n23183 );
not ( n23185 , n23184 );
and ( n23186 , n23169 , n23185 );
not ( n23187 , n23169 );
and ( n23188 , n23187 , n23184 );
nor ( n23189 , n23186 , n23188 );
not ( n23190 , n23189 );
not ( n23191 , n23190 );
not ( n23192 , n19091 );
not ( n23193 , n12813 );
not ( n23194 , n12825 );
xor ( n23195 , n23193 , n23194 );
xnor ( n23196 , n23195 , n12831 );
not ( n23197 , n23196 );
or ( n23198 , n23192 , n23197 );
or ( n23199 , n23196 , n19091 );
nand ( n23200 , n23198 , n23199 );
buf ( n23201 , n12809 );
and ( n23202 , n23200 , n23201 );
not ( n23203 , n23200 );
not ( n23204 , n23201 );
and ( n23205 , n23203 , n23204 );
nor ( n23206 , n23202 , n23205 );
buf ( n23207 , n17533 );
not ( n23208 , n23207 );
not ( n23209 , n20336 );
not ( n23210 , n23209 );
or ( n23211 , n23208 , n23210 );
or ( n23212 , n23209 , n23207 );
nand ( n23213 , n23211 , n23212 );
and ( n23214 , n23213 , n8888 );
not ( n23215 , n23213 );
and ( n23216 , n23215 , n18897 );
nor ( n23217 , n23214 , n23216 );
not ( n23218 , n23217 );
nand ( n23219 , n23206 , n23218 );
buf ( n23220 , n7649 );
not ( n23221 , n23220 );
not ( n23222 , n16452 );
or ( n23223 , n23221 , n23222 );
not ( n23224 , n23220 );
nand ( n23225 , n23224 , n16453 );
nand ( n23226 , n23223 , n23225 );
not ( n23227 , n23226 );
not ( n23228 , n16493 );
and ( n23229 , n23227 , n23228 );
and ( n23230 , n23226 , n16493 );
nor ( n23231 , n23229 , n23230 );
buf ( n23232 , n23231 );
xor ( n23233 , n23219 , n23232 );
not ( n23234 , n23233 );
not ( n23235 , n23234 );
or ( n23236 , n23191 , n23235 );
nand ( n23237 , n23233 , n23189 );
nand ( n23238 , n23236 , n23237 );
buf ( n23239 , n20619 );
xor ( n23240 , n22244 , n23239 );
not ( n23241 , n21513 );
and ( n23242 , n21539 , n21184 );
not ( n23243 , n21539 );
not ( n23244 , n21183 );
and ( n23245 , n23243 , n23244 );
nor ( n23246 , n23242 , n23245 );
not ( n23247 , n23246 );
not ( n23248 , n23247 );
or ( n23249 , n23241 , n23248 );
not ( n23250 , n21513 );
nand ( n23251 , n23246 , n23250 );
nand ( n23252 , n23249 , n23251 );
buf ( n23253 , n23252 );
xnor ( n23254 , n23240 , n23253 );
buf ( n23255 , n6347 );
nand ( n23256 , n7912 , n23255 );
buf ( n23257 , n6348 );
not ( n23258 , n23257 );
and ( n23259 , n23256 , n23258 );
not ( n23260 , n23256 );
buf ( n23261 , n23257 );
and ( n23262 , n23260 , n23261 );
nor ( n23263 , n23259 , n23262 );
not ( n23264 , n23263 );
not ( n23265 , n7315 );
or ( n23266 , n23264 , n23265 );
not ( n23267 , n23263 );
nand ( n23268 , n23267 , n7318 );
nand ( n23269 , n23266 , n23268 );
and ( n23270 , n23269 , n11755 );
not ( n23271 , n23269 );
and ( n23272 , n23271 , n16151 );
nor ( n23273 , n23270 , n23272 );
nand ( n23274 , n23254 , n23273 );
not ( n23275 , n23274 );
not ( n23276 , n14729 );
not ( n23277 , n16257 );
or ( n23278 , n23276 , n23277 );
not ( n23279 , n14728 );
nand ( n23280 , n16258 , n23279 );
nand ( n23281 , n23278 , n23280 );
and ( n23282 , n23281 , n19622 );
not ( n23283 , n23281 );
not ( n23284 , n19619 );
not ( n23285 , n23284 );
and ( n23286 , n23283 , n23285 );
nor ( n23287 , n23282 , n23286 );
not ( n23288 , n23287 );
and ( n23289 , n23275 , n23288 );
and ( n23290 , n23274 , n23287 );
nor ( n23291 , n23289 , n23290 );
and ( n23292 , n23238 , n23291 );
not ( n23293 , n23238 );
not ( n23294 , n23291 );
and ( n23295 , n23293 , n23294 );
nor ( n23296 , n23292 , n23295 );
not ( n23297 , n23296 );
not ( n23298 , n17935 );
not ( n23299 , n8663 );
or ( n23300 , n23298 , n23299 );
nand ( n23301 , n10864 , n17932 );
nand ( n23302 , n23300 , n23301 );
buf ( n23303 , n6349 );
buf ( n23304 , n6350 );
buf ( n23305 , n23304 );
not ( n23306 , n23305 );
buf ( n23307 , n6351 );
not ( n23308 , n23307 );
not ( n23309 , n23308 );
or ( n23310 , n23306 , n23309 );
not ( n23311 , n23304 );
buf ( n23312 , n23307 );
nand ( n23313 , n23311 , n23312 );
nand ( n23314 , n23310 , n23313 );
xor ( n23315 , n23303 , n23314 );
buf ( n23316 , n6352 );
buf ( n23317 , n6353 );
xor ( n23318 , n23316 , n23317 );
buf ( n23319 , n6354 );
nand ( n23320 , n10874 , n23319 );
xnor ( n23321 , n23318 , n23320 );
xnor ( n23322 , n23315 , n23321 );
buf ( n23323 , n23322 );
buf ( n23324 , n23323 );
not ( n23325 , n23324 );
and ( n23326 , n23302 , n23325 );
not ( n23327 , n23302 );
and ( n23328 , n23327 , n23324 );
nor ( n23329 , n23326 , n23328 );
not ( n23330 , n23329 );
not ( n23331 , n23330 );
not ( n23332 , n23331 );
buf ( n23333 , n11542 );
not ( n23334 , n23333 );
not ( n23335 , n11539 );
and ( n23336 , n23334 , n23335 );
and ( n23337 , n23333 , n11539 );
nor ( n23338 , n23336 , n23337 );
and ( n23339 , n23338 , n7367 );
not ( n23340 , n23338 );
not ( n23341 , n7370 );
and ( n23342 , n23340 , n23341 );
nor ( n23343 , n23339 , n23342 );
not ( n23344 , n7412 );
and ( n23345 , n23343 , n23344 );
not ( n23346 , n23343 );
and ( n23347 , n23346 , n7412 );
nor ( n23348 , n23345 , n23347 );
not ( n23349 , n23348 );
buf ( n23350 , n16596 );
xor ( n23351 , n19738 , n23350 );
xnor ( n23352 , n23351 , n21803 );
not ( n23353 , n23352 );
nand ( n23354 , n23349 , n23353 );
not ( n23355 , n23354 );
or ( n23356 , n23332 , n23355 );
or ( n23357 , n23354 , n23331 );
nand ( n23358 , n23356 , n23357 );
not ( n23359 , n23358 );
buf ( n23360 , n10743 );
xor ( n23361 , n10154 , n10174 );
buf ( n23362 , n10163 );
xnor ( n23363 , n23361 , n23362 );
buf ( n23364 , n23363 );
xor ( n23365 , n23360 , n23364 );
xnor ( n23366 , n23365 , n13254 );
not ( n23367 , n23366 );
buf ( n23368 , n12808 );
not ( n23369 , n23368 );
not ( n23370 , n23369 );
not ( n23371 , n9374 );
or ( n23372 , n23370 , n23371 );
not ( n23373 , n9374 );
nand ( n23374 , n23373 , n23368 );
nand ( n23375 , n23372 , n23374 );
not ( n23376 , n22802 );
buf ( n23377 , n23376 );
xnor ( n23378 , n23375 , n23377 );
not ( n23379 , n23378 );
nand ( n23380 , n23367 , n23379 );
not ( n23381 , n23380 );
xor ( n23382 , n18688 , n17707 );
not ( n23383 , n7991 );
buf ( n23384 , n23383 );
xnor ( n23385 , n23382 , n23384 );
not ( n23386 , n23385 );
and ( n23387 , n23381 , n23386 );
and ( n23388 , n23380 , n23385 );
nor ( n23389 , n23387 , n23388 );
not ( n23390 , n23389 );
or ( n23391 , n23359 , n23390 );
or ( n23392 , n23389 , n23358 );
nand ( n23393 , n23391 , n23392 );
not ( n23394 , n23393 );
or ( n23395 , n23297 , n23394 );
or ( n23396 , n23393 , n23296 );
nand ( n23397 , n23395 , n23396 );
buf ( n23398 , n23397 );
not ( n23399 , n23398 );
not ( n23400 , n23399 );
or ( n23401 , n23167 , n23400 );
not ( n23402 , n23166 );
nand ( n23403 , n23402 , n23398 );
nand ( n23404 , n23401 , n23403 );
not ( n23405 , n10351 );
not ( n23406 , n9641 );
not ( n23407 , n23406 );
not ( n23408 , n10394 );
not ( n23409 , n23408 );
or ( n23410 , n23407 , n23409 );
or ( n23411 , n10398 , n23406 );
nand ( n23412 , n23410 , n23411 );
not ( n23413 , n23412 );
and ( n23414 , n23405 , n23413 );
and ( n23415 , n10351 , n23412 );
nor ( n23416 , n23414 , n23415 );
not ( n23417 , n23416 );
not ( n23418 , n23417 );
not ( n23419 , n17544 );
not ( n23420 , n23419 );
not ( n23421 , n7772 );
and ( n23422 , n23420 , n23421 );
and ( n23423 , n23419 , n7772 );
nor ( n23424 , n23422 , n23423 );
and ( n23425 , n23424 , n17590 );
not ( n23426 , n23424 );
and ( n23427 , n23426 , n17603 );
nor ( n23428 , n23425 , n23427 );
not ( n23429 , n23428 );
buf ( n23430 , n6355 );
not ( n23431 , n23430 );
not ( n23432 , n18955 );
not ( n23433 , n23432 );
not ( n23434 , n23433 );
or ( n23435 , n23431 , n23434 );
or ( n23436 , n23433 , n23430 );
nand ( n23437 , n23435 , n23436 );
not ( n23438 , n23437 );
not ( n23439 , n19218 );
not ( n23440 , n23439 );
not ( n23441 , n19237 );
or ( n23442 , n23440 , n23441 );
nand ( n23443 , n19236 , n19218 );
nand ( n23444 , n23442 , n23443 );
not ( n23445 , n23444 );
not ( n23446 , n23445 );
or ( n23447 , n23438 , n23446 );
not ( n23448 , n23437 );
buf ( n23449 , n23444 );
nand ( n23450 , n23448 , n23449 );
nand ( n23451 , n23447 , n23450 );
nand ( n23452 , n23429 , n23451 );
not ( n23453 , n23452 );
or ( n23454 , n23418 , n23453 );
or ( n23455 , n23452 , n23417 );
nand ( n23456 , n23454 , n23455 );
not ( n23457 , n23456 );
not ( n23458 , n14577 );
not ( n23459 , n8409 );
and ( n23460 , n23458 , n23459 );
and ( n23461 , n14577 , n8409 );
nor ( n23462 , n23460 , n23461 );
and ( n23463 , n23462 , n14627 );
not ( n23464 , n23462 );
and ( n23465 , n23464 , n14624 );
nor ( n23466 , n23463 , n23465 );
not ( n23467 , n23466 );
not ( n23468 , n11131 );
nand ( n23469 , n23468 , n9785 );
not ( n23470 , n23469 );
nor ( n23471 , n9785 , n11135 );
nor ( n23472 , n23470 , n23471 );
not ( n23473 , n23472 );
not ( n23474 , n9844 );
not ( n23475 , n23474 );
or ( n23476 , n23473 , n23475 );
not ( n23477 , n23472 );
nand ( n23478 , n23477 , n9844 );
nand ( n23479 , n23476 , n23478 );
nand ( n23480 , n23467 , n23479 );
not ( n23481 , n23480 );
not ( n23482 , n10004 );
buf ( n23483 , n6356 );
buf ( n23484 , n23483 );
not ( n23485 , n23484 );
not ( n23486 , n21363 );
not ( n23487 , n23486 );
or ( n23488 , n23485 , n23487 );
not ( n23489 , n23483 );
nand ( n23490 , n23489 , n21364 );
nand ( n23491 , n23488 , n23490 );
buf ( n23492 , n6357 );
not ( n23493 , n23492 );
and ( n23494 , n23491 , n23493 );
not ( n23495 , n23491 );
buf ( n23496 , n23492 );
and ( n23497 , n23495 , n23496 );
nor ( n23498 , n23494 , n23497 );
buf ( n23499 , n6358 );
nand ( n23500 , n8954 , n23499 );
buf ( n23501 , n6359 );
buf ( n23502 , n23501 );
and ( n23503 , n23500 , n23502 );
not ( n23504 , n23500 );
not ( n23505 , n23501 );
and ( n23506 , n23504 , n23505 );
nor ( n23507 , n23503 , n23506 );
xor ( n23508 , n23498 , n23507 );
buf ( n23509 , n6360 );
nand ( n23510 , n8032 , n23509 );
buf ( n23511 , n6361 );
buf ( n23512 , n23511 );
and ( n23513 , n23510 , n23512 );
not ( n23514 , n23510 );
not ( n23515 , n23511 );
and ( n23516 , n23514 , n23515 );
nor ( n23517 , n23513 , n23516 );
xor ( n23518 , n23508 , n23517 );
not ( n23519 , n23518 );
not ( n23520 , n23519 );
not ( n23521 , n23520 );
or ( n23522 , n23482 , n23521 );
buf ( n23523 , n23518 );
or ( n23524 , n23523 , n10004 );
nand ( n23525 , n23522 , n23524 );
xor ( n23526 , n20134 , n20143 );
xnor ( n23527 , n23526 , n20153 );
not ( n23528 , n23527 );
not ( n23529 , n23528 );
not ( n23530 , n23529 );
and ( n23531 , n23525 , n23530 );
not ( n23532 , n23525 );
buf ( n23533 , n23527 );
and ( n23534 , n23532 , n23533 );
nor ( n23535 , n23531 , n23534 );
not ( n23536 , n23535 );
not ( n23537 , n23536 );
and ( n23538 , n23481 , n23537 );
and ( n23539 , n23480 , n23536 );
nor ( n23540 , n23538 , n23539 );
not ( n23541 , n23540 );
or ( n23542 , n23457 , n23541 );
or ( n23543 , n23540 , n23456 );
nand ( n23544 , n23542 , n23543 );
buf ( n23545 , n6362 );
buf ( n23546 , n23545 );
xor ( n23547 , n23546 , n19200 );
not ( n23548 , n20089 );
xnor ( n23549 , n23547 , n23548 );
not ( n23550 , n23549 );
xor ( n23551 , n11703 , n12651 );
buf ( n23552 , n16770 );
xor ( n23553 , n23552 , n16778 );
xor ( n23554 , n23553 , n16794 );
not ( n23555 , n23554 );
xnor ( n23556 , n23551 , n23555 );
not ( n23557 , n23556 );
nand ( n23558 , n23550 , n23557 );
not ( n23559 , n17956 );
not ( n23560 , n10865 );
or ( n23561 , n23559 , n23560 );
or ( n23562 , n10865 , n17956 );
nand ( n23563 , n23561 , n23562 );
and ( n23564 , n23563 , n23325 );
not ( n23565 , n23563 );
and ( n23566 , n23565 , n23324 );
nor ( n23567 , n23564 , n23566 );
not ( n23568 , n23567 );
and ( n23569 , n23558 , n23568 );
not ( n23570 , n23558 );
and ( n23571 , n23570 , n23567 );
nor ( n23572 , n23569 , n23571 );
and ( n23573 , n23544 , n23572 );
not ( n23574 , n23544 );
not ( n23575 , n23572 );
and ( n23576 , n23574 , n23575 );
nor ( n23577 , n23573 , n23576 );
not ( n23578 , n23577 );
not ( n23579 , n23578 );
not ( n23580 , n11926 );
not ( n23581 , n9461 );
not ( n23582 , n23581 );
or ( n23583 , n23580 , n23582 );
or ( n23584 , n9465 , n11926 );
nand ( n23585 , n23583 , n23584 );
not ( n23586 , n22536 );
not ( n23587 , n23586 );
xor ( n23588 , n23585 , n23587 );
not ( n23589 , n23588 );
not ( n23590 , n9253 );
not ( n23591 , n17716 );
or ( n23592 , n23590 , n23591 );
not ( n23593 , n17716 );
nand ( n23594 , n23593 , n9249 );
nand ( n23595 , n23592 , n23594 );
and ( n23596 , n23595 , n17721 );
not ( n23597 , n23595 );
buf ( n23598 , n8140 );
and ( n23599 , n23597 , n23598 );
nor ( n23600 , n23596 , n23599 );
nand ( n23601 , n23589 , n23600 );
not ( n23602 , n23601 );
xor ( n23603 , n14837 , n10912 );
xnor ( n23604 , n23603 , n13718 );
not ( n23605 , n23604 );
not ( n23606 , n23605 );
or ( n23607 , n23602 , n23606 );
or ( n23608 , n23605 , n23601 );
nand ( n23609 , n23607 , n23608 );
not ( n23610 , n23609 );
not ( n23611 , n21227 );
not ( n23612 , n21146 );
or ( n23613 , n23611 , n23612 );
not ( n23614 , n21146 );
nand ( n23615 , n23614 , n21223 );
nand ( n23616 , n23613 , n23615 );
buf ( n23617 , n22180 );
and ( n23618 , n23616 , n23617 );
not ( n23619 , n23616 );
buf ( n23620 , n22187 );
and ( n23621 , n23619 , n23620 );
nor ( n23622 , n23618 , n23621 );
not ( n23623 , n22345 );
not ( n23624 , n15974 );
or ( n23625 , n23623 , n23624 );
nand ( n23626 , n20846 , n22341 );
nand ( n23627 , n23625 , n23626 );
not ( n23628 , n22554 );
and ( n23629 , n23627 , n23628 );
not ( n23630 , n23627 );
and ( n23631 , n23630 , n22554 );
nor ( n23632 , n23629 , n23631 );
and ( n23633 , n23622 , n23632 );
buf ( n23634 , n12530 );
not ( n23635 , n23634 );
not ( n23636 , n10126 );
not ( n23637 , n23636 );
or ( n23638 , n23635 , n23637 );
or ( n23639 , n23636 , n23634 );
nand ( n23640 , n23638 , n23639 );
and ( n23641 , n23640 , n18528 );
not ( n23642 , n23640 );
not ( n23643 , n18528 );
and ( n23644 , n23642 , n23643 );
nor ( n23645 , n23641 , n23644 );
not ( n23646 , n23645 );
not ( n23647 , n23646 );
and ( n23648 , n23633 , n23647 );
not ( n23649 , n23633 );
and ( n23650 , n23649 , n23646 );
nor ( n23651 , n23648 , n23650 );
not ( n23652 , n23651 );
and ( n23653 , n23610 , n23652 );
and ( n23654 , n23609 , n23651 );
nor ( n23655 , n23653 , n23654 );
not ( n23656 , n23655 );
not ( n23657 , n23656 );
and ( n23658 , n23579 , n23657 );
and ( n23659 , n23578 , n23656 );
nor ( n23660 , n23658 , n23659 );
buf ( n23661 , n23660 );
and ( n23662 , n23404 , n23661 );
not ( n23663 , n23404 );
not ( n23664 , n23655 );
not ( n23665 , n23577 );
or ( n23666 , n23664 , n23665 );
not ( n23667 , n23577 );
nand ( n23668 , n23667 , n23656 );
nand ( n23669 , n23666 , n23668 );
not ( n23670 , n23669 );
not ( n23671 , n23670 );
and ( n23672 , n23663 , n23671 );
nor ( n23673 , n23662 , n23672 );
buf ( n23674 , n6363 );
buf ( n23675 , n23674 );
not ( n23676 , n23675 );
buf ( n23677 , n6364 );
not ( n23678 , n23677 );
not ( n23679 , n23678 );
or ( n23680 , n23676 , n23679 );
not ( n23681 , n23674 );
buf ( n23682 , n23677 );
nand ( n23683 , n23681 , n23682 );
nand ( n23684 , n23680 , n23683 );
buf ( n23685 , n6365 );
buf ( n23686 , n23685 );
and ( n23687 , n23684 , n23686 );
not ( n23688 , n23684 );
not ( n23689 , n23685 );
and ( n23690 , n23688 , n23689 );
nor ( n23691 , n23687 , n23690 );
xor ( n23692 , n23691 , n11767 );
xnor ( n23693 , n23692 , n23263 );
buf ( n23694 , n23693 );
xor ( n23695 , n20749 , n23694 );
xnor ( n23696 , n23695 , n8314 );
not ( n23697 , n23696 );
buf ( n23698 , n11082 );
xor ( n23699 , n11817 , n23698 );
xnor ( n23700 , n23699 , n9844 );
not ( n23701 , n13021 );
not ( n23702 , n21992 );
or ( n23703 , n23701 , n23702 );
nand ( n23704 , n14997 , n13017 );
nand ( n23705 , n23703 , n23704 );
and ( n23706 , n23705 , n15047 );
not ( n23707 , n23705 );
and ( n23708 , n23707 , n15055 );
nor ( n23709 , n23706 , n23708 );
not ( n23710 , n23709 );
nand ( n23711 , n23700 , n23710 );
not ( n23712 , n23711 );
or ( n23713 , n23697 , n23712 );
not ( n23714 , n23709 );
nand ( n23715 , n23714 , n23700 );
or ( n23716 , n23715 , n23696 );
nand ( n23717 , n23713 , n23716 );
not ( n23718 , n23717 );
not ( n23719 , n19315 );
not ( n23720 , n15290 );
or ( n23721 , n23719 , n23720 );
not ( n23722 , n19315 );
not ( n23723 , n15290 );
nand ( n23724 , n23722 , n23723 );
nand ( n23725 , n23721 , n23724 );
and ( n23726 , n23725 , n14225 );
not ( n23727 , n23725 );
and ( n23728 , n23727 , n14221 );
nor ( n23729 , n23726 , n23728 );
not ( n23730 , n23729 );
not ( n23731 , n9530 );
not ( n23732 , n13927 );
xor ( n23733 , n17260 , n23732 );
xnor ( n23734 , n23733 , n13934 );
not ( n23735 , n23734 );
or ( n23736 , n23731 , n23735 );
or ( n23737 , n23734 , n9530 );
nand ( n23738 , n23736 , n23737 );
not ( n23739 , n17040 );
and ( n23740 , n23738 , n23739 );
not ( n23741 , n23738 );
and ( n23742 , n23741 , n17044 );
nor ( n23743 , n23740 , n23742 );
nand ( n23744 , n23730 , n23743 );
not ( n23745 , n23744 );
not ( n23746 , n10533 );
not ( n23747 , n15744 );
or ( n23748 , n23746 , n23747 );
or ( n23749 , n15744 , n10533 );
nand ( n23750 , n23748 , n23749 );
nor ( n23751 , n23750 , n10010 );
not ( n23752 , n23751 );
nand ( n23753 , n10011 , n23750 );
nand ( n23754 , n23752 , n23753 );
not ( n23755 , n23754 );
and ( n23756 , n23745 , n23755 );
not ( n23757 , n23729 );
nand ( n23758 , n23757 , n23743 );
and ( n23759 , n23758 , n23754 );
nor ( n23760 , n23756 , n23759 );
not ( n23761 , n23760 );
not ( n23762 , n21750 );
not ( n23763 , n18461 );
or ( n23764 , n23762 , n23763 );
not ( n23765 , n21750 );
nand ( n23766 , n23765 , n15689 );
nand ( n23767 , n23764 , n23766 );
not ( n23768 , n18465 );
and ( n23769 , n23767 , n23768 );
not ( n23770 , n23767 );
and ( n23771 , n23770 , n18465 );
nor ( n23772 , n23769 , n23771 );
buf ( n23773 , n15412 );
not ( n23774 , n23773 );
not ( n23775 , n19746 );
or ( n23776 , n23774 , n23775 );
or ( n23777 , n19746 , n23773 );
nand ( n23778 , n23776 , n23777 );
not ( n23779 , n16983 );
and ( n23780 , n23778 , n23779 );
not ( n23781 , n23778 );
and ( n23782 , n23781 , n16983 );
nor ( n23783 , n23780 , n23782 );
nand ( n23784 , n23772 , n23783 );
buf ( n23785 , n6366 );
nand ( n23786 , n8966 , n23785 );
buf ( n23787 , n6367 );
not ( n23788 , n23787 );
and ( n23789 , n23786 , n23788 );
not ( n23790 , n23786 );
buf ( n23791 , n23787 );
and ( n23792 , n23790 , n23791 );
nor ( n23793 , n23789 , n23792 );
buf ( n23794 , n23793 );
not ( n23795 , n11745 );
xor ( n23796 , n11734 , n23795 );
xnor ( n23797 , n23796 , n11753 );
xor ( n23798 , n23794 , n23797 );
not ( n23799 , n16147 );
not ( n23800 , n23799 );
xnor ( n23801 , n23798 , n23800 );
not ( n23802 , n23801 );
and ( n23803 , n23784 , n23802 );
not ( n23804 , n23784 );
and ( n23805 , n23804 , n23801 );
nor ( n23806 , n23803 , n23805 );
not ( n23807 , n23806 );
and ( n23808 , n23761 , n23807 );
and ( n23809 , n23760 , n23806 );
nor ( n23810 , n23808 , n23809 );
not ( n23811 , n23810 );
or ( n23812 , n23718 , n23811 );
or ( n23813 , n23717 , n23810 );
nand ( n23814 , n23812 , n23813 );
not ( n23815 , n16146 );
not ( n23816 , n18003 );
or ( n23817 , n23815 , n23816 );
not ( n23818 , n16146 );
nand ( n23819 , n23818 , n18004 );
nand ( n23820 , n23817 , n23819 );
not ( n23821 , n13984 );
not ( n23822 , n23821 );
buf ( n23823 , n23822 );
and ( n23824 , n23820 , n23823 );
not ( n23825 , n23820 );
buf ( n23826 , n13991 );
buf ( n23827 , n23826 );
and ( n23828 , n23825 , n23827 );
nor ( n23829 , n23824 , n23828 );
not ( n23830 , n23829 );
not ( n23831 , n23830 );
buf ( n23832 , n22234 );
not ( n23833 , n23832 );
not ( n23834 , n21540 );
or ( n23835 , n23833 , n23834 );
or ( n23836 , n21540 , n23832 );
nand ( n23837 , n23835 , n23836 );
and ( n23838 , n23837 , n23239 );
not ( n23839 , n23837 );
buf ( n23840 , n20625 );
and ( n23841 , n23839 , n23840 );
nor ( n23842 , n23838 , n23841 );
not ( n23843 , n21422 );
not ( n23844 , n18166 );
or ( n23845 , n23843 , n23844 );
or ( n23846 , n18166 , n21422 );
nand ( n23847 , n23845 , n23846 );
and ( n23848 , n23847 , n7992 );
not ( n23849 , n23847 );
and ( n23850 , n23849 , n7993 );
nor ( n23851 , n23848 , n23850 );
nand ( n23852 , n23842 , n23851 );
not ( n23853 , n23852 );
or ( n23854 , n23831 , n23853 );
or ( n23855 , n23852 , n23830 );
nand ( n23856 , n23854 , n23855 );
not ( n23857 , n23856 );
buf ( n23858 , n22045 );
xor ( n23859 , n7409 , n23858 );
xnor ( n23860 , n23859 , n18261 );
not ( n23861 , n14724 );
not ( n23862 , n16257 );
or ( n23863 , n23861 , n23862 );
nand ( n23864 , n16258 , n14720 );
nand ( n23865 , n23863 , n23864 );
and ( n23866 , n23865 , n19622 );
not ( n23867 , n23865 );
and ( n23868 , n23867 , n23285 );
nor ( n23869 , n23866 , n23868 );
nand ( n23870 , n23860 , n23869 );
not ( n23871 , n23870 );
not ( n23872 , n12031 );
and ( n23873 , n12035 , n23872 );
not ( n23874 , n12035 );
and ( n23875 , n23874 , n12032 );
nor ( n23876 , n23873 , n23875 );
not ( n23877 , n23876 );
not ( n23878 , n14311 );
or ( n23879 , n23877 , n23878 );
or ( n23880 , n14311 , n23876 );
nand ( n23881 , n23879 , n23880 );
not ( n23882 , n20901 );
buf ( n23883 , n6368 );
not ( n23884 , n23883 );
not ( n23885 , n23884 );
or ( n23886 , n23882 , n23885 );
not ( n23887 , n20900 );
buf ( n23888 , n23883 );
nand ( n23889 , n23887 , n23888 );
nand ( n23890 , n23886 , n23889 );
buf ( n23891 , n6369 );
buf ( n23892 , n23891 );
and ( n23893 , n23890 , n23892 );
not ( n23894 , n23890 );
not ( n23895 , n23891 );
and ( n23896 , n23894 , n23895 );
nor ( n23897 , n23893 , n23896 );
not ( n23898 , n23897 );
xor ( n23899 , n23898 , n19000 );
buf ( n23900 , n6370 );
nand ( n23901 , n8455 , n23900 );
buf ( n23902 , n6371 );
buf ( n23903 , n23902 );
and ( n23904 , n23901 , n23903 );
not ( n23905 , n23901 );
not ( n23906 , n23902 );
and ( n23907 , n23905 , n23906 );
nor ( n23908 , n23904 , n23907 );
not ( n23909 , n23908 );
xnor ( n23910 , n23899 , n23909 );
not ( n23911 , n23910 );
not ( n23912 , n23911 );
and ( n23913 , n23881 , n23912 );
not ( n23914 , n23881 );
xor ( n23915 , n23897 , n23908 );
xnor ( n23916 , n23915 , n19001 );
buf ( n23917 , n23916 );
and ( n23918 , n23914 , n23917 );
nor ( n23919 , n23913 , n23918 );
not ( n23920 , n23919 );
and ( n23921 , n23871 , n23920 );
and ( n23922 , n23870 , n23919 );
nor ( n23923 , n23921 , n23922 );
not ( n23924 , n23923 );
or ( n23925 , n23857 , n23924 );
or ( n23926 , n23923 , n23856 );
nand ( n23927 , n23925 , n23926 );
and ( n23928 , n23814 , n23927 );
not ( n23929 , n23814 );
not ( n23930 , n23927 );
and ( n23931 , n23929 , n23930 );
nor ( n23932 , n23928 , n23931 );
not ( n23933 , n23932 );
not ( n23934 , n23933 );
not ( n23935 , n8617 );
not ( n23936 , n6982 );
or ( n23937 , n23935 , n23936 );
not ( n23938 , n8617 );
nand ( n23939 , n23938 , n6977 );
nand ( n23940 , n23937 , n23939 );
and ( n23941 , n23940 , n7029 );
not ( n23942 , n23940 );
and ( n23943 , n23942 , n7025 );
nor ( n23944 , n23941 , n23943 );
not ( n23945 , n18460 );
not ( n23946 , n23945 );
buf ( n23947 , n6372 );
buf ( n23948 , n23947 );
not ( n23949 , n23948 );
buf ( n23950 , n6373 );
not ( n23951 , n23950 );
not ( n23952 , n23951 );
or ( n23953 , n23949 , n23952 );
not ( n23954 , n23947 );
buf ( n23955 , n23950 );
nand ( n23956 , n23954 , n23955 );
nand ( n23957 , n23953 , n23956 );
buf ( n23958 , n6374 );
buf ( n23959 , n23958 );
and ( n23960 , n23957 , n23959 );
not ( n23961 , n23957 );
not ( n23962 , n23958 );
and ( n23963 , n23961 , n23962 );
nor ( n23964 , n23960 , n23963 );
buf ( n23965 , n6375 );
nand ( n23966 , n7197 , n23965 );
buf ( n23967 , n6376 );
buf ( n23968 , n23967 );
and ( n23969 , n23966 , n23968 );
not ( n23970 , n23966 );
not ( n23971 , n23967 );
and ( n23972 , n23970 , n23971 );
nor ( n23973 , n23969 , n23972 );
xor ( n23974 , n23964 , n23973 );
buf ( n23975 , n6377 );
nand ( n23976 , n8223 , n23975 );
buf ( n23977 , n6378 );
not ( n23978 , n23977 );
and ( n23979 , n23976 , n23978 );
not ( n23980 , n23976 );
buf ( n23981 , n23977 );
and ( n23982 , n23980 , n23981 );
nor ( n23983 , n23979 , n23982 );
xnor ( n23984 , n23974 , n23983 );
not ( n23985 , n23984 );
or ( n23986 , n23946 , n23985 );
or ( n23987 , n23984 , n23945 );
nand ( n23988 , n23986 , n23987 );
and ( n23989 , n23988 , n10090 );
not ( n23990 , n23988 );
not ( n23991 , n10088 );
not ( n23992 , n23991 );
and ( n23993 , n23990 , n23992 );
nor ( n23994 , n23989 , n23993 );
not ( n23995 , n23994 );
nand ( n23996 , n23944 , n23995 );
not ( n23997 , n23996 );
not ( n23998 , n13259 );
xor ( n23999 , n20386 , n20405 );
not ( n24000 , n20395 );
xnor ( n24001 , n23999 , n24000 );
not ( n24002 , n24001 );
or ( n24003 , n23998 , n24002 );
or ( n24004 , n24001 , n13259 );
nand ( n24005 , n24003 , n24004 );
and ( n24006 , n24005 , n14793 );
not ( n24007 , n24005 );
and ( n24008 , n24007 , n14794 );
nor ( n24009 , n24006 , n24008 );
not ( n24010 , n24009 );
and ( n24011 , n23997 , n24010 );
and ( n24012 , n23996 , n24009 );
nor ( n24013 , n24011 , n24012 );
buf ( n24014 , n24013 );
not ( n24015 , n24014 );
not ( n24016 , n24015 );
buf ( n24017 , n6379 );
buf ( n24018 , n24017 );
not ( n24019 , n24018 );
buf ( n24020 , n6380 );
not ( n24021 , n24020 );
not ( n24022 , n24021 );
or ( n24023 , n24019 , n24022 );
not ( n24024 , n24017 );
buf ( n24025 , n24020 );
nand ( n24026 , n24024 , n24025 );
nand ( n24027 , n24023 , n24026 );
buf ( n24028 , n6381 );
not ( n24029 , n24028 );
and ( n24030 , n24027 , n24029 );
not ( n24031 , n24027 );
buf ( n24032 , n24028 );
and ( n24033 , n24031 , n24032 );
nor ( n24034 , n24030 , n24033 );
buf ( n24035 , n6382 );
nand ( n24036 , n7977 , n24035 );
buf ( n24037 , n6383 );
buf ( n24038 , n24037 );
and ( n24039 , n24036 , n24038 );
not ( n24040 , n24036 );
not ( n24041 , n24037 );
and ( n24042 , n24040 , n24041 );
nor ( n24043 , n24039 , n24042 );
xor ( n24044 , n24034 , n24043 );
buf ( n24045 , n6384 );
nand ( n24046 , n11946 , n24045 );
buf ( n24047 , n6385 );
not ( n24048 , n24047 );
and ( n24049 , n24046 , n24048 );
not ( n24050 , n24046 );
buf ( n24051 , n24047 );
and ( n24052 , n24050 , n24051 );
nor ( n24053 , n24049 , n24052 );
xor ( n24054 , n24044 , n24053 );
buf ( n24055 , n24054 );
not ( n24056 , n24055 );
xor ( n24057 , n10931 , n24056 );
buf ( n24058 , n9277 );
xnor ( n24059 , n24057 , n24058 );
buf ( n24060 , n7011 );
not ( n24061 , n24060 );
buf ( n24062 , n6386 );
buf ( n24063 , n24062 );
not ( n24064 , n24063 );
buf ( n24065 , n6387 );
not ( n24066 , n24065 );
not ( n24067 , n24066 );
or ( n24068 , n24064 , n24067 );
not ( n24069 , n24062 );
buf ( n24070 , n24065 );
nand ( n24071 , n24069 , n24070 );
nand ( n24072 , n24068 , n24071 );
and ( n24073 , n24072 , n16109 );
not ( n24074 , n24072 );
not ( n24075 , n16108 );
and ( n24076 , n24074 , n24075 );
nor ( n24077 , n24073 , n24076 );
xor ( n24078 , n24077 , n23793 );
xnor ( n24079 , n24078 , n18786 );
not ( n24080 , n24079 );
buf ( n24081 , n24080 );
not ( n24082 , n24081 );
or ( n24083 , n24061 , n24082 );
or ( n24084 , n24081 , n24060 );
nand ( n24085 , n24083 , n24084 );
buf ( n24086 , n18154 );
and ( n24087 , n24085 , n24086 );
not ( n24088 , n24085 );
not ( n24089 , n24086 );
and ( n24090 , n24088 , n24089 );
nor ( n24091 , n24087 , n24090 );
not ( n24092 , n24091 );
nand ( n24093 , n24059 , n24092 );
not ( n24094 , n24093 );
buf ( n24095 , n12208 );
not ( n24096 , n24095 );
not ( n24097 , n23239 );
or ( n24098 , n24096 , n24097 );
or ( n24099 , n23239 , n24095 );
nand ( n24100 , n24098 , n24099 );
and ( n24101 , n24100 , n20631 );
not ( n24102 , n24100 );
and ( n24103 , n24102 , n20628 );
nor ( n24104 , n24101 , n24103 );
not ( n24105 , n24104 );
not ( n24106 , n24105 );
and ( n24107 , n24094 , n24106 );
and ( n24108 , n24093 , n24105 );
nor ( n24109 , n24107 , n24108 );
not ( n24110 , n24109 );
not ( n24111 , n24110 );
buf ( n24112 , n11062 );
xor ( n24113 , n24112 , n11074 );
xor ( n24114 , n24113 , n11081 );
buf ( n24115 , n24114 );
xor ( n24116 , n11797 , n24115 );
xnor ( n24117 , n24116 , n9844 );
not ( n24118 , n24117 );
buf ( n24119 , n7986 );
not ( n24120 , n24119 );
not ( n24121 , n22860 );
or ( n24122 , n24120 , n24121 );
not ( n24123 , n24119 );
nand ( n24124 , n24123 , n22864 );
nand ( n24125 , n24122 , n24124 );
and ( n24126 , n24125 , n22867 );
not ( n24127 , n24125 );
and ( n24128 , n24127 , n14508 );
nor ( n24129 , n24126 , n24128 );
not ( n24130 , n24129 );
nand ( n24131 , n24118 , n24130 );
not ( n24132 , n23363 );
not ( n24133 , n24132 );
xor ( n24134 , n10708 , n24133 );
xnor ( n24135 , n24134 , n13254 );
and ( n24136 , n24131 , n24135 );
not ( n24137 , n24131 );
not ( n24138 , n24135 );
and ( n24139 , n24137 , n24138 );
nor ( n24140 , n24136 , n24139 );
not ( n24141 , n24140 );
not ( n24142 , n24141 );
or ( n24143 , n24111 , n24142 );
nand ( n24144 , n24140 , n24109 );
nand ( n24145 , n24143 , n24144 );
not ( n24146 , n11321 );
not ( n24147 , n22606 );
or ( n24148 , n24146 , n24147 );
or ( n24149 , n22606 , n11321 );
nand ( n24150 , n24148 , n24149 );
and ( n24151 , n24150 , n17332 );
not ( n24152 , n24150 );
and ( n24153 , n24152 , n17347 );
nor ( n24154 , n24151 , n24153 );
not ( n24155 , n24154 );
not ( n24156 , n24155 );
not ( n24157 , n20903 );
buf ( n24158 , n14308 );
not ( n24159 , n24158 );
not ( n24160 , n24159 );
not ( n24161 , n12341 );
or ( n24162 , n24160 , n24161 );
nand ( n24163 , n13294 , n24158 );
nand ( n24164 , n24162 , n24163 );
not ( n24165 , n24164 );
and ( n24166 , n24157 , n24165 );
and ( n24167 , n12376 , n24164 );
nor ( n24168 , n24166 , n24167 );
not ( n24169 , n24168 );
nand ( n24170 , n24156 , n24169 );
not ( n24171 , n24170 );
not ( n24172 , n15387 );
not ( n24173 , n19739 );
or ( n24174 , n24172 , n24173 );
not ( n24175 , n15387 );
nand ( n24176 , n24175 , n19746 );
nand ( n24177 , n24174 , n24176 );
and ( n24178 , n24177 , n16984 );
not ( n24179 , n24177 );
and ( n24180 , n24179 , n16983 );
nor ( n24181 , n24178 , n24180 );
not ( n24182 , n24181 );
not ( n24183 , n24182 );
and ( n24184 , n24171 , n24183 );
and ( n24185 , n24170 , n24182 );
nor ( n24186 , n24184 , n24185 );
not ( n24187 , n24186 );
not ( n24188 , n24009 );
not ( n24189 , n23944 );
nand ( n24190 , n24188 , n24189 );
not ( n24191 , n17882 );
not ( n24192 , n15254 );
not ( n24193 , n22180 );
or ( n24194 , n24192 , n24193 );
not ( n24195 , n15254 );
nand ( n24196 , n24195 , n22187 );
nand ( n24197 , n24194 , n24196 );
not ( n24198 , n24197 );
or ( n24199 , n24191 , n24198 );
or ( n24200 , n22139 , n24197 );
nand ( n24201 , n24199 , n24200 );
buf ( n24202 , n24201 );
xnor ( n24203 , n24190 , n24202 );
not ( n24204 , n24203 );
or ( n24205 , n24187 , n24204 );
or ( n24206 , n24203 , n24186 );
nand ( n24207 , n24205 , n24206 );
not ( n24208 , n16212 );
not ( n24209 , n6658 );
not ( n24210 , n24209 );
buf ( n24211 , n12430 );
not ( n24212 , n24211 );
and ( n24213 , n24210 , n24212 );
not ( n24214 , n6659 );
and ( n24215 , n24214 , n24211 );
nor ( n24216 , n24213 , n24215 );
not ( n24217 , n24216 );
or ( n24218 , n24208 , n24217 );
or ( n24219 , n24216 , n16212 );
nand ( n24220 , n24218 , n24219 );
not ( n24221 , n16125 );
not ( n24222 , n18003 );
or ( n24223 , n24221 , n24222 );
or ( n24224 , n18003 , n16125 );
nand ( n24225 , n24223 , n24224 );
and ( n24226 , n24225 , n23827 );
not ( n24227 , n24225 );
and ( n24228 , n24227 , n23823 );
nor ( n24229 , n24226 , n24228 );
not ( n24230 , n24229 );
nand ( n24231 , n24220 , n24230 );
not ( n24232 , n24231 );
xor ( n24233 , n15024 , n11394 );
xnor ( n24234 , n24233 , n23003 );
not ( n24235 , n24234 );
not ( n24236 , n24235 );
and ( n24237 , n24232 , n24236 );
and ( n24238 , n24231 , n24235 );
nor ( n24239 , n24237 , n24238 );
and ( n24240 , n24207 , n24239 );
not ( n24241 , n24207 );
not ( n24242 , n24239 );
and ( n24243 , n24241 , n24242 );
nor ( n24244 , n24240 , n24243 );
xor ( n24245 , n24145 , n24244 );
not ( n24246 , n24245 );
or ( n24247 , n24016 , n24246 );
not ( n24248 , n24244 );
not ( n24249 , n24248 );
not ( n24250 , n24145 );
not ( n24251 , n24250 );
or ( n24252 , n24249 , n24251 );
nand ( n24253 , n24145 , n24244 );
nand ( n24254 , n24252 , n24253 );
nand ( n24255 , n24254 , n24014 );
nand ( n24256 , n24247 , n24255 );
not ( n24257 , n24256 );
or ( n24258 , n23934 , n24257 );
buf ( n24259 , n23932 );
not ( n24260 , n24259 );
or ( n24261 , n24256 , n24260 );
nand ( n24262 , n24258 , n24261 );
not ( n24263 , n24262 );
nand ( n24264 , n23673 , n24263 );
not ( n24265 , n20590 );
not ( n24266 , n7879 );
or ( n24267 , n24265 , n24266 );
or ( n24268 , n7879 , n20590 );
nand ( n24269 , n24267 , n24268 );
not ( n24270 , n12833 );
and ( n24271 , n24269 , n24270 );
not ( n24272 , n24269 );
and ( n24273 , n24272 , n17688 );
nor ( n24274 , n24271 , n24273 );
not ( n24275 , n24274 );
nand ( n24276 , n16199 , n24275 );
not ( n24277 , n24276 );
buf ( n24278 , n7785 );
not ( n24279 , n24278 );
not ( n24280 , n23419 );
not ( n24281 , n24280 );
or ( n24282 , n24279 , n24281 );
not ( n24283 , n17546 );
or ( n24284 , n24283 , n24278 );
nand ( n24285 , n24282 , n24284 );
buf ( n24286 , n17603 );
and ( n24287 , n24285 , n24286 );
not ( n24288 , n24285 );
and ( n24289 , n24288 , n17590 );
nor ( n24290 , n24287 , n24289 );
not ( n24291 , n24290 );
and ( n24292 , n24277 , n24291 );
and ( n24293 , n24276 , n24290 );
nor ( n24294 , n24292 , n24293 );
not ( n24295 , n24294 );
not ( n24296 , n24290 );
nand ( n24297 , n24274 , n24296 );
buf ( n24298 , n16106 );
and ( n24299 , n24297 , n24298 );
not ( n24300 , n24297 );
not ( n24301 , n24298 );
and ( n24302 , n24300 , n24301 );
nor ( n24303 , n24299 , n24302 );
not ( n24304 , n24303 );
not ( n24305 , n24304 );
buf ( n24306 , n8122 );
not ( n24307 , n24306 );
not ( n24308 , n6685 );
or ( n24309 , n24307 , n24308 );
or ( n24310 , n6685 , n24306 );
nand ( n24311 , n24309 , n24310 );
buf ( n24312 , n22959 );
and ( n24313 , n24311 , n24312 );
not ( n24314 , n24311 );
not ( n24315 , n22959 );
and ( n24316 , n24314 , n24315 );
nor ( n24317 , n24313 , n24316 );
not ( n24318 , n19903 );
not ( n24319 , n17611 );
or ( n24320 , n24318 , n24319 );
not ( n24321 , n17611 );
nand ( n24322 , n24321 , n19899 );
nand ( n24323 , n24320 , n24322 );
and ( n24324 , n24323 , n13744 );
not ( n24325 , n24323 );
and ( n24326 , n24325 , n13731 );
nor ( n24327 , n24324 , n24326 );
nand ( n24328 , n24317 , n24327 );
and ( n24329 , n24328 , n16264 );
not ( n24330 , n24328 );
not ( n24331 , n16264 );
and ( n24332 , n24330 , n24331 );
nor ( n24333 , n24329 , n24332 );
not ( n24334 , n24333 );
not ( n24335 , n24334 );
or ( n24336 , n24305 , n24335 );
nand ( n24337 , n24333 , n24303 );
nand ( n24338 , n24336 , n24337 );
not ( n24339 , n24338 );
not ( n24340 , n24339 );
not ( n24341 , n8012 );
buf ( n24342 , n6388 );
nand ( n24343 , n8537 , n24342 );
buf ( n24344 , n6389 );
buf ( n24345 , n24344 );
and ( n24346 , n24343 , n24345 );
not ( n24347 , n24343 );
not ( n24348 , n24344 );
and ( n24349 , n24347 , n24348 );
nor ( n24350 , n24346 , n24349 );
not ( n24351 , n24350 );
buf ( n24352 , n6390 );
nand ( n24353 , n7912 , n24352 );
buf ( n24354 , n6391 );
not ( n24355 , n24354 );
and ( n24356 , n24353 , n24355 );
not ( n24357 , n24353 );
buf ( n24358 , n24354 );
and ( n24359 , n24357 , n24358 );
nor ( n24360 , n24356 , n24359 );
not ( n24361 , n24360 );
or ( n24362 , n24351 , n24361 );
or ( n24363 , n24350 , n24360 );
nand ( n24364 , n24362 , n24363 );
not ( n24365 , n18023 );
buf ( n24366 , n6392 );
not ( n24367 , n24366 );
not ( n24368 , n24367 );
or ( n24369 , n24365 , n24368 );
not ( n24370 , n18022 );
buf ( n24371 , n24366 );
nand ( n24372 , n24370 , n24371 );
nand ( n24373 , n24369 , n24372 );
buf ( n24374 , n6393 );
buf ( n24375 , n24374 );
and ( n24376 , n24373 , n24375 );
not ( n24377 , n24373 );
not ( n24378 , n24374 );
and ( n24379 , n24377 , n24378 );
nor ( n24380 , n24376 , n24379 );
xnor ( n24381 , n24364 , n24380 );
not ( n24382 , n24381 );
or ( n24383 , n24341 , n24382 );
xor ( n24384 , n24380 , n24350 );
xnor ( n24385 , n24384 , n24360 );
nand ( n24386 , n24385 , n8008 );
nand ( n24387 , n24383 , n24386 );
not ( n24388 , n24387 );
not ( n24389 , n22863 );
and ( n24390 , n24388 , n24389 );
and ( n24391 , n24387 , n22860 );
nor ( n24392 , n24390 , n24391 );
not ( n24393 , n24392 );
not ( n24394 , n16905 );
not ( n24395 , n24394 );
not ( n24396 , n18710 );
or ( n24397 , n24395 , n24396 );
or ( n24398 , n18710 , n24394 );
nand ( n24399 , n24397 , n24398 );
and ( n24400 , n24399 , n12342 );
not ( n24401 , n24399 );
and ( n24402 , n24401 , n18714 );
nor ( n24403 , n24400 , n24402 );
nand ( n24404 , n24393 , n24403 );
and ( n24405 , n24404 , n15842 );
not ( n24406 , n24404 );
and ( n24407 , n24406 , n15843 );
nor ( n24408 , n24405 , n24407 );
not ( n24409 , n24408 );
not ( n24410 , n24409 );
not ( n24411 , n18474 );
buf ( n24412 , n6394 );
not ( n24413 , n24412 );
not ( n24414 , n24413 );
or ( n24415 , n24411 , n24414 );
not ( n24416 , n18473 );
buf ( n24417 , n24412 );
nand ( n24418 , n24416 , n24417 );
nand ( n24419 , n24415 , n24418 );
not ( n24420 , n21300 );
and ( n24421 , n24419 , n24420 );
not ( n24422 , n24419 );
and ( n24423 , n24422 , n21301 );
nor ( n24424 , n24421 , n24423 );
buf ( n24425 , n6395 );
nand ( n24426 , n10372 , n24425 );
buf ( n24427 , n6396 );
buf ( n24428 , n24427 );
and ( n24429 , n24426 , n24428 );
not ( n24430 , n24426 );
not ( n24431 , n24427 );
and ( n24432 , n24430 , n24431 );
nor ( n24433 , n24429 , n24432 );
xor ( n24434 , n24424 , n24433 );
xnor ( n24435 , n24434 , n20427 );
buf ( n24436 , n24435 );
not ( n24437 , n24436 );
not ( n24438 , n17872 );
buf ( n24439 , n6397 );
buf ( n24440 , n24439 );
not ( n24441 , n24440 );
not ( n24442 , n7628 );
not ( n24443 , n24442 );
or ( n24444 , n24441 , n24443 );
not ( n24445 , n24439 );
nand ( n24446 , n24445 , n7629 );
nand ( n24447 , n24444 , n24446 );
and ( n24448 , n24447 , n19557 );
not ( n24449 , n24447 );
and ( n24450 , n24449 , n19554 );
nor ( n24451 , n24448 , n24450 );
buf ( n24452 , n6398 );
nand ( n24453 , n8454 , n24452 );
buf ( n24454 , n6399 );
buf ( n24455 , n24454 );
and ( n24456 , n24453 , n24455 );
not ( n24457 , n24453 );
not ( n24458 , n24454 );
and ( n24459 , n24457 , n24458 );
nor ( n24460 , n24456 , n24459 );
xor ( n24461 , n24451 , n24460 );
buf ( n24462 , n6400 );
nand ( n24463 , n6558 , n24462 );
buf ( n24464 , n6401 );
not ( n24465 , n24464 );
and ( n24466 , n24463 , n24465 );
not ( n24467 , n24463 );
buf ( n24468 , n24464 );
and ( n24469 , n24467 , n24468 );
nor ( n24470 , n24466 , n24469 );
xnor ( n24471 , n24461 , n24470 );
buf ( n24472 , n24471 );
not ( n24473 , n24472 );
or ( n24474 , n24438 , n24473 );
not ( n24475 , n24451 );
xor ( n24476 , n24475 , n24460 );
xnor ( n24477 , n24476 , n24470 );
nand ( n24478 , n24477 , n17869 );
nand ( n24479 , n24474 , n24478 );
not ( n24480 , n24479 );
or ( n24481 , n24437 , n24480 );
or ( n24482 , n24479 , n24436 );
nand ( n24483 , n24481 , n24482 );
nand ( n24484 , n15383 , n24483 );
and ( n24485 , n24484 , n15477 );
not ( n24486 , n24484 );
and ( n24487 , n24486 , n15478 );
nor ( n24488 , n24485 , n24487 );
not ( n24489 , n24488 );
not ( n24490 , n24489 );
or ( n24491 , n24410 , n24490 );
nand ( n24492 , n24488 , n24408 );
nand ( n24493 , n24491 , n24492 );
buf ( n24494 , n6402 );
not ( n24495 , n24494 );
buf ( n24496 , n6403 );
buf ( n24497 , n24496 );
and ( n24498 , n24495 , n24497 );
not ( n24499 , n24495 );
not ( n24500 , n24496 );
and ( n24501 , n24499 , n24500 );
nor ( n24502 , n24498 , n24501 );
xor ( n24503 , n11628 , n24502 );
buf ( n24504 , n6404 );
not ( n24505 , n24504 );
buf ( n24506 , n6405 );
nand ( n24507 , n6916 , n24506 );
buf ( n24508 , n6406 );
buf ( n24509 , n24508 );
and ( n24510 , n24507 , n24509 );
not ( n24511 , n24507 );
not ( n24512 , n24508 );
and ( n24513 , n24511 , n24512 );
nor ( n24514 , n24510 , n24513 );
not ( n24515 , n24514 );
or ( n24516 , n24505 , n24515 );
or ( n24517 , n24514 , n24504 );
nand ( n24518 , n24516 , n24517 );
xnor ( n24519 , n24503 , n24518 );
xor ( n24520 , n19170 , n24519 );
buf ( n24521 , n17139 );
and ( n24522 , n24520 , n24521 );
not ( n24523 , n24520 );
buf ( n24524 , n9898 );
and ( n24525 , n24523 , n24524 );
nor ( n24526 , n24522 , n24525 );
not ( n24527 , n24526 );
not ( n24528 , n18103 );
not ( n24529 , n9513 );
or ( n24530 , n24528 , n24529 );
or ( n24531 , n9513 , n18103 );
nand ( n24532 , n24530 , n24531 );
xnor ( n24533 , n24532 , n9562 );
nand ( n24534 , n24527 , n24533 );
not ( n24535 , n24534 );
buf ( n24536 , n15642 );
not ( n24537 , n24536 );
not ( n24538 , n24537 );
and ( n24539 , n24535 , n24538 );
and ( n24540 , n24534 , n24537 );
nor ( n24541 , n24539 , n24540 );
and ( n24542 , n24493 , n24541 );
not ( n24543 , n24493 );
not ( n24544 , n24541 );
and ( n24545 , n24543 , n24544 );
nor ( n24546 , n24542 , n24545 );
not ( n24547 , n24546 );
not ( n24548 , n24547 );
or ( n24549 , n24340 , n24548 );
nand ( n24550 , n24546 , n24338 );
nand ( n24551 , n24549 , n24550 );
not ( n24552 , n24551 );
or ( n24553 , n24295 , n24552 );
or ( n24554 , n24551 , n24294 );
nand ( n24555 , n24553 , n24554 );
not ( n24556 , n24555 );
xor ( n24557 , n19456 , n17614 );
xnor ( n24558 , n24557 , n13547 );
not ( n24559 , n24558 );
buf ( n24560 , n20828 );
xor ( n24561 , n17977 , n24560 );
xor ( n24562 , n24561 , n23324 );
not ( n24563 , n24562 );
nand ( n24564 , n24559 , n24563 );
not ( n24565 , n16687 );
xor ( n24566 , n24564 , n24565 );
not ( n24567 , n24566 );
not ( n24568 , n24567 );
xor ( n24569 , n20755 , n23694 );
not ( n24570 , n8317 );
xnor ( n24571 , n24569 , n24570 );
not ( n24572 , n24571 );
not ( n24573 , n14967 );
not ( n24574 , n18821 );
not ( n24575 , n24574 );
not ( n24576 , n24575 );
or ( n24577 , n24573 , n24576 );
or ( n24578 , n18822 , n14967 );
nand ( n24579 , n24577 , n24578 );
and ( n24580 , n24579 , n23003 );
not ( n24581 , n24579 );
buf ( n24582 , n22976 );
xor ( n24583 , n24582 , n22986 );
xnor ( n24584 , n24583 , n22993 );
and ( n24585 , n24581 , n24584 );
nor ( n24586 , n24580 , n24585 );
not ( n24587 , n24586 );
nand ( n24588 , n24572 , n24587 );
not ( n24589 , n24588 );
not ( n24590 , n16372 );
and ( n24591 , n24589 , n24590 );
and ( n24592 , n24588 , n16372 );
nor ( n24593 , n24591 , n24592 );
not ( n24594 , n24593 );
not ( n24595 , n24594 );
or ( n24596 , n24568 , n24595 );
nand ( n24597 , n24593 , n24566 );
nand ( n24598 , n24596 , n24597 );
buf ( n24599 , n6407 );
not ( n24600 , n24599 );
not ( n24601 , n23916 );
or ( n24602 , n24600 , n24601 );
or ( n24603 , n23916 , n24599 );
nand ( n24604 , n24602 , n24603 );
and ( n24605 , n24604 , n21361 );
not ( n24606 , n24604 );
and ( n24607 , n24606 , n21360 );
nor ( n24608 , n24605 , n24607 );
not ( n24609 , n10063 );
not ( n24610 , n15428 );
or ( n24611 , n24609 , n24610 );
or ( n24612 , n15424 , n10063 );
nand ( n24613 , n24611 , n24612 );
and ( n24614 , n24613 , n15475 );
not ( n24615 , n24613 );
and ( n24616 , n24615 , n15474 );
nor ( n24617 , n24614 , n24616 );
not ( n24618 , n24617 );
nand ( n24619 , n24608 , n24618 );
not ( n24620 , n24619 );
not ( n24621 , n16807 );
and ( n24622 , n24620 , n24621 );
and ( n24623 , n24619 , n16807 );
nor ( n24624 , n24622 , n24623 );
not ( n24625 , n24624 );
not ( n24626 , n14949 );
not ( n24627 , n7502 );
not ( n24628 , n14911 );
or ( n24629 , n24627 , n24628 );
or ( n24630 , n14911 , n7502 );
nand ( n24631 , n24629 , n24630 );
not ( n24632 , n24631 );
or ( n24633 , n24626 , n24632 );
not ( n24634 , n24631 );
nand ( n24635 , n24634 , n14942 );
nand ( n24636 , n24633 , n24635 );
not ( n24637 , n24636 );
not ( n24638 , n8245 );
not ( n24639 , n17332 );
or ( n24640 , n24638 , n24639 );
not ( n24641 , n8245 );
nand ( n24642 , n24641 , n17345 );
nand ( n24643 , n24640 , n24642 );
and ( n24644 , n24643 , n8992 );
not ( n24645 , n24643 );
not ( n24646 , n7270 );
and ( n24647 , n24645 , n24646 );
nor ( n24648 , n24644 , n24647 );
not ( n24649 , n24648 );
nand ( n24650 , n24637 , n24649 );
not ( n24651 , n16920 );
and ( n24652 , n24650 , n24651 );
not ( n24653 , n24650 );
and ( n24654 , n24653 , n16920 );
nor ( n24655 , n24652 , n24654 );
not ( n24656 , n24655 );
or ( n24657 , n24625 , n24656 );
or ( n24658 , n24655 , n24624 );
nand ( n24659 , n24657 , n24658 );
not ( n24660 , n24385 );
not ( n24661 , n24660 );
xor ( n24662 , n18171 , n24661 );
buf ( n24663 , n6408 );
buf ( n24664 , n6409 );
buf ( n24665 , n24664 );
not ( n24666 , n24665 );
buf ( n24667 , n6410 );
not ( n24668 , n24667 );
not ( n24669 , n24668 );
or ( n24670 , n24666 , n24669 );
not ( n24671 , n24664 );
buf ( n24672 , n24667 );
nand ( n24673 , n24671 , n24672 );
nand ( n24674 , n24670 , n24673 );
xor ( n24675 , n24663 , n24674 );
buf ( n24676 , n6411 );
xor ( n24677 , n24676 , n8679 );
xnor ( n24678 , n24677 , n8677 );
xnor ( n24679 , n24675 , n24678 );
not ( n24680 , n24679 );
not ( n24681 , n24680 );
not ( n24682 , n24681 );
xnor ( n24683 , n24662 , n24682 );
not ( n24684 , n24683 );
not ( n24685 , n9113 );
not ( n24686 , n19200 );
or ( n24687 , n24685 , n24686 );
or ( n24688 , n19200 , n9113 );
nand ( n24689 , n24687 , n24688 );
and ( n24690 , n24689 , n21060 );
not ( n24691 , n24689 );
and ( n24692 , n24691 , n21063 );
nor ( n24693 , n24690 , n24692 );
not ( n24694 , n24693 );
nand ( n24695 , n24684 , n24694 );
not ( n24696 , n24695 );
buf ( n24697 , n16499 );
not ( n24698 , n24697 );
and ( n24699 , n24696 , n24698 );
and ( n24700 , n24695 , n24697 );
nor ( n24701 , n24699 , n24700 );
and ( n24702 , n24659 , n24701 );
not ( n24703 , n24659 );
not ( n24704 , n24701 );
and ( n24705 , n24703 , n24704 );
nor ( n24706 , n24702 , n24705 );
and ( n24707 , n24598 , n24706 );
not ( n24708 , n24598 );
not ( n24709 , n24706 );
and ( n24710 , n24708 , n24709 );
nor ( n24711 , n24707 , n24710 );
not ( n24712 , n24711 );
not ( n24713 , n24712 );
not ( n24714 , n24713 );
and ( n24715 , n24556 , n24714 );
and ( n24716 , n24555 , n24713 );
nor ( n24717 , n24715 , n24716 );
nor ( n24718 , n24717 , n20975 );
not ( n24719 , n24718 );
or ( n24720 , n24264 , n24719 );
not ( n24721 , n24717 );
not ( n24722 , n24721 );
not ( n24723 , n23673 );
or ( n24724 , n24722 , n24723 );
nor ( n24725 , n24263 , n17807 );
nand ( n24726 , n24724 , n24725 );
buf ( n24727 , n13353 );
nand ( n24728 , n24727 , n7374 );
nand ( n24729 , n24720 , n24726 , n24728 );
buf ( n24730 , n24729 );
buf ( n24731 , n24730 );
buf ( n24732 , n20975 );
not ( n24733 , n24732 );
not ( n24734 , n21770 );
not ( n24735 , n24734 );
not ( n24736 , n24735 );
not ( n24737 , n18462 );
or ( n24738 , n24736 , n24737 );
or ( n24739 , n18462 , n24735 );
nand ( n24740 , n24738 , n24739 );
and ( n24741 , n24740 , n18465 );
not ( n24742 , n24740 );
and ( n24743 , n24742 , n23768 );
nor ( n24744 , n24741 , n24743 );
not ( n24745 , n24744 );
buf ( n24746 , n7177 );
not ( n24747 , n24746 );
not ( n24748 , n18863 );
or ( n24749 , n24747 , n24748 );
not ( n24750 , n19450 );
or ( n24751 , n24750 , n24746 );
nand ( n24752 , n24749 , n24751 );
xor ( n24753 , n18806 , n18810 );
not ( n24754 , n18820 );
xnor ( n24755 , n24753 , n24754 );
and ( n24756 , n24752 , n24755 );
not ( n24757 , n24752 );
and ( n24758 , n24757 , n18823 );
nor ( n24759 , n24756 , n24758 );
not ( n24760 , n24759 );
nand ( n24761 , n24745 , n24760 );
not ( n24762 , n13656 );
not ( n24763 , n19471 );
or ( n24764 , n24762 , n24763 );
or ( n24765 , n19471 , n13656 );
nand ( n24766 , n24764 , n24765 );
not ( n24767 , n21883 );
not ( n24768 , n24767 );
and ( n24769 , n24766 , n24768 );
not ( n24770 , n24766 );
and ( n24771 , n24770 , n24767 );
nor ( n24772 , n24769 , n24771 );
and ( n24773 , n24761 , n24772 );
not ( n24774 , n24761 );
not ( n24775 , n24772 );
and ( n24776 , n24774 , n24775 );
nor ( n24777 , n24773 , n24776 );
not ( n24778 , n24777 );
not ( n24779 , n18111 );
buf ( n24780 , n6412 );
nand ( n24781 , n6633 , n24780 );
buf ( n24782 , n6413 );
buf ( n24783 , n24782 );
and ( n24784 , n24781 , n24783 );
not ( n24785 , n24781 );
not ( n24786 , n24782 );
and ( n24787 , n24785 , n24786 );
nor ( n24788 , n24784 , n24787 );
buf ( n24789 , n24788 );
not ( n24790 , n24789 );
not ( n24791 , n18154 );
not ( n24792 , n24791 );
or ( n24793 , n24790 , n24792 );
or ( n24794 , n24791 , n24789 );
nand ( n24795 , n24793 , n24794 );
and ( n24796 , n24779 , n24795 );
not ( n24797 , n24779 );
not ( n24798 , n24795 );
and ( n24799 , n24797 , n24798 );
nor ( n24800 , n24796 , n24799 );
not ( n24801 , n8812 );
not ( n24802 , n8836 );
or ( n24803 , n24801 , n24802 );
nand ( n24804 , n24803 , n8840 );
xor ( n24805 , n9439 , n24804 );
xnor ( n24806 , n24805 , n18889 );
nand ( n24807 , n24800 , n24806 );
not ( n24808 , n24807 );
not ( n24809 , n19366 );
not ( n24810 , n24018 );
not ( n24811 , n8135 );
or ( n24812 , n24810 , n24811 );
or ( n24813 , n8135 , n24018 );
nand ( n24814 , n24812 , n24813 );
not ( n24815 , n24814 );
or ( n24816 , n24809 , n24815 );
or ( n24817 , n24814 , n19370 );
nand ( n24818 , n24816 , n24817 );
not ( n24819 , n24818 );
and ( n24820 , n24808 , n24819 );
and ( n24821 , n24807 , n24818 );
nor ( n24822 , n24820 , n24821 );
not ( n24823 , n24822 );
not ( n24824 , n12072 );
not ( n24825 , n7223 );
or ( n24826 , n24824 , n24825 );
not ( n24827 , n12072 );
nand ( n24828 , n24827 , n13515 );
nand ( n24829 , n24826 , n24828 );
and ( n24830 , n24829 , n7189 );
not ( n24831 , n24829 );
not ( n24832 , n7189 );
and ( n24833 , n24831 , n24832 );
nor ( n24834 , n24830 , n24833 );
buf ( n24835 , n19671 );
not ( n24836 , n24835 );
not ( n24837 , n9940 );
or ( n24838 , n24836 , n24837 );
or ( n24839 , n9940 , n24835 );
nand ( n24840 , n24838 , n24839 );
xor ( n24841 , n24840 , n20337 );
nand ( n24842 , n24834 , n24841 );
not ( n24843 , n22938 );
not ( n24844 , n6861 );
not ( n24845 , n14447 );
or ( n24846 , n24844 , n24845 );
nand ( n24847 , n14446 , n6857 );
nand ( n24848 , n24846 , n24847 );
not ( n24849 , n24848 );
and ( n24850 , n24843 , n24849 );
and ( n24851 , n22938 , n24848 );
nor ( n24852 , n24850 , n24851 );
and ( n24853 , n24842 , n24852 );
not ( n24854 , n24842 );
not ( n24855 , n24852 );
and ( n24856 , n24854 , n24855 );
nor ( n24857 , n24853 , n24856 );
not ( n24858 , n24857 );
or ( n24859 , n24823 , n24858 );
or ( n24860 , n24857 , n24822 );
nand ( n24861 , n24859 , n24860 );
not ( n24862 , n13504 );
buf ( n24863 , n6414 );
not ( n24864 , n24863 );
not ( n24865 , n24864 );
or ( n24866 , n24862 , n24865 );
not ( n24867 , n13503 );
buf ( n24868 , n24863 );
nand ( n24869 , n24867 , n24868 );
nand ( n24870 , n24866 , n24869 );
buf ( n24871 , n6415 );
not ( n24872 , n24871 );
and ( n24873 , n24870 , n24872 );
not ( n24874 , n24870 );
buf ( n24875 , n24871 );
and ( n24876 , n24874 , n24875 );
nor ( n24877 , n24873 , n24876 );
buf ( n24878 , n6416 );
nand ( n24879 , n7247 , n24878 );
buf ( n24880 , n6417 );
buf ( n24881 , n24880 );
and ( n24882 , n24879 , n24881 );
not ( n24883 , n24879 );
not ( n24884 , n24880 );
and ( n24885 , n24883 , n24884 );
nor ( n24886 , n24882 , n24885 );
xor ( n24887 , n24877 , n24886 );
xnor ( n24888 , n24887 , n23142 );
not ( n24889 , n24888 );
buf ( n24890 , n24889 );
xor ( n24891 , n18236 , n24890 );
buf ( n24892 , n6418 );
buf ( n24893 , n24892 );
not ( n24894 , n24893 );
buf ( n24895 , n6419 );
not ( n24896 , n24895 );
not ( n24897 , n24896 );
or ( n24898 , n24894 , n24897 );
not ( n24899 , n24892 );
buf ( n24900 , n24895 );
nand ( n24901 , n24899 , n24900 );
nand ( n24902 , n24898 , n24901 );
not ( n24903 , n24902 );
buf ( n24904 , n6420 );
buf ( n24905 , n6421 );
nand ( n24906 , n6770 , n24905 );
buf ( n24907 , n6422 );
buf ( n24908 , n24907 );
and ( n24909 , n24906 , n24908 );
not ( n24910 , n24906 );
not ( n24911 , n24907 );
and ( n24912 , n24910 , n24911 );
nor ( n24913 , n24909 , n24912 );
xor ( n24914 , n24904 , n24913 );
buf ( n24915 , n6423 );
nand ( n24916 , n6515 , n24915 );
buf ( n24917 , n6424 );
not ( n24918 , n24917 );
and ( n24919 , n24916 , n24918 );
not ( n24920 , n24916 );
buf ( n24921 , n24917 );
and ( n24922 , n24920 , n24921 );
nor ( n24923 , n24919 , n24922 );
xnor ( n24924 , n24914 , n24923 );
xor ( n24925 , n24903 , n24924 );
xnor ( n24926 , n24891 , n24925 );
not ( n24927 , n7104 );
not ( n24928 , n19526 );
or ( n24929 , n24927 , n24928 );
or ( n24930 , n19527 , n7104 );
nand ( n24931 , n24929 , n24930 );
not ( n24932 , n24931 );
not ( n24933 , n19480 );
or ( n24934 , n24932 , n24933 );
or ( n24935 , n19480 , n24931 );
nand ( n24936 , n24934 , n24935 );
not ( n24937 , n24936 );
nand ( n24938 , n24926 , n24937 );
not ( n24939 , n24938 );
not ( n24940 , n14761 );
not ( n24941 , n13711 );
or ( n24942 , n24940 , n24941 );
not ( n24943 , n14761 );
nand ( n24944 , n24943 , n7450 );
nand ( n24945 , n24942 , n24944 );
xor ( n24946 , n24945 , n13718 );
not ( n24947 , n24946 );
not ( n24948 , n24947 );
and ( n24949 , n24939 , n24948 );
and ( n24950 , n24938 , n24947 );
nor ( n24951 , n24949 , n24950 );
and ( n24952 , n24861 , n24951 );
not ( n24953 , n24861 );
not ( n24954 , n24951 );
and ( n24955 , n24953 , n24954 );
nor ( n24956 , n24952 , n24955 );
nand ( n24957 , n24772 , n24759 );
not ( n24958 , n24957 );
not ( n24959 , n10099 );
xor ( n24960 , n15449 , n15458 );
xor ( n24961 , n24960 , n15468 );
not ( n24962 , n24961 );
or ( n24963 , n24959 , n24962 );
or ( n24964 , n15469 , n10099 );
nand ( n24965 , n24963 , n24964 );
and ( n24966 , n24965 , n22821 );
not ( n24967 , n24965 );
and ( n24968 , n24967 , n22817 );
nor ( n24969 , n24966 , n24968 );
not ( n24970 , n24969 );
and ( n24971 , n24958 , n24970 );
and ( n24972 , n24957 , n24969 );
nor ( n24973 , n24971 , n24972 );
not ( n24974 , n24973 );
not ( n24975 , n21359 );
and ( n24976 , n23496 , n24975 );
not ( n24977 , n23496 );
and ( n24978 , n24977 , n21361 );
or ( n24979 , n24976 , n24978 );
and ( n24980 , n24979 , n17098 );
not ( n24981 , n24979 );
and ( n24982 , n24981 , n21319 );
nor ( n24983 , n24980 , n24982 );
not ( n24984 , n11748 );
and ( n24985 , n11752 , n24984 );
not ( n24986 , n11752 );
and ( n24987 , n24986 , n11749 );
nor ( n24988 , n24985 , n24987 );
not ( n24989 , n24988 );
not ( n24990 , n20208 );
or ( n24991 , n24989 , n24990 );
not ( n24992 , n20208 );
not ( n24993 , n24988 );
nand ( n24994 , n24992 , n24993 );
nand ( n24995 , n24991 , n24994 );
and ( n24996 , n24995 , n18003 );
not ( n24997 , n24995 );
and ( n24998 , n24997 , n18004 );
nor ( n24999 , n24996 , n24998 );
not ( n25000 , n24999 );
nand ( n25001 , n24983 , n25000 );
not ( n25002 , n7765 );
not ( n25003 , n23419 );
or ( n25004 , n25002 , n25003 );
or ( n25005 , n17546 , n7765 );
nand ( n25006 , n25004 , n25005 );
and ( n25007 , n25006 , n24286 );
not ( n25008 , n25006 );
and ( n25009 , n25008 , n17590 );
nor ( n25010 , n25007 , n25009 );
not ( n25011 , n25010 );
and ( n25012 , n25001 , n25011 );
not ( n25013 , n25001 );
and ( n25014 , n25013 , n25010 );
nor ( n25015 , n25012 , n25014 );
not ( n25016 , n25015 );
or ( n25017 , n24974 , n25016 );
or ( n25018 , n25015 , n24973 );
nand ( n25019 , n25017 , n25018 );
and ( n25020 , n24956 , n25019 );
not ( n25021 , n24956 );
not ( n25022 , n25019 );
and ( n25023 , n25021 , n25022 );
nor ( n25024 , n25020 , n25023 );
not ( n25025 , n25024 );
or ( n25026 , n24778 , n25025 );
not ( n25027 , n24777 );
not ( n25028 , n25024 );
nand ( n25029 , n25027 , n25028 );
nand ( n25030 , n25026 , n25029 );
not ( n25031 , n6698 );
not ( n25032 , n14051 );
or ( n25033 , n25031 , n25032 );
not ( n25034 , n6698 );
nand ( n25035 , n25034 , n14048 );
nand ( n25036 , n25033 , n25035 );
and ( n25037 , n25036 , n14095 );
not ( n25038 , n25036 );
not ( n25039 , n14092 );
buf ( n25040 , n25039 );
not ( n25041 , n25040 );
and ( n25042 , n25038 , n25041 );
nor ( n25043 , n25037 , n25042 );
not ( n25044 , n25043 );
buf ( n25045 , n24043 );
not ( n25046 , n25045 );
not ( n25047 , n8139 );
or ( n25048 , n25046 , n25047 );
or ( n25049 , n8139 , n25045 );
nand ( n25050 , n25048 , n25049 );
and ( n25051 , n25050 , n19366 );
not ( n25052 , n25050 );
and ( n25053 , n25052 , n19371 );
nor ( n25054 , n25051 , n25053 );
nand ( n25055 , n25044 , n25054 );
not ( n25056 , n25055 );
buf ( n25057 , n18851 );
xor ( n25058 , n25057 , n7128 );
xnor ( n25059 , n25058 , n18612 );
not ( n25060 , n25059 );
or ( n25061 , n25056 , n25060 );
or ( n25062 , n25059 , n25055 );
nand ( n25063 , n25061 , n25062 );
not ( n25064 , n25063 );
not ( n25065 , n25064 );
not ( n25066 , n24975 );
buf ( n25067 , n23507 );
not ( n25068 , n25067 );
and ( n25069 , n25066 , n25068 );
and ( n25070 , n21360 , n25067 );
nor ( n25071 , n25069 , n25070 );
not ( n25072 , n25071 );
not ( n25073 , n17101 );
or ( n25074 , n25072 , n25073 );
or ( n25075 , n17101 , n25071 );
nand ( n25076 , n25074 , n25075 );
not ( n25077 , n25076 );
not ( n25078 , n14798 );
not ( n25079 , n25078 );
not ( n25080 , n25079 );
not ( n25081 , n13268 );
not ( n25082 , n24001 );
or ( n25083 , n25081 , n25082 );
buf ( n25084 , n24001 );
or ( n25085 , n25084 , n13268 );
nand ( n25086 , n25083 , n25085 );
not ( n25087 , n25086 );
or ( n25088 , n25080 , n25087 );
or ( n25089 , n25086 , n20415 );
nand ( n25090 , n25088 , n25089 );
nand ( n25091 , n25077 , n25090 );
not ( n25092 , n13490 );
not ( n25093 , n22549 );
or ( n25094 , n25092 , n25093 );
or ( n25095 , n22549 , n13490 );
nand ( n25096 , n25094 , n25095 );
not ( n25097 , n19447 );
and ( n25098 , n25096 , n25097 );
not ( n25099 , n25096 );
not ( n25100 , n19443 );
and ( n25101 , n25099 , n25100 );
nor ( n25102 , n25098 , n25101 );
not ( n25103 , n25102 );
and ( n25104 , n25091 , n25103 );
not ( n25105 , n25091 );
and ( n25106 , n25105 , n25102 );
nor ( n25107 , n25104 , n25106 );
not ( n25108 , n25107 );
not ( n25109 , n25108 );
or ( n25110 , n25065 , n25109 );
nand ( n25111 , n25063 , n25107 );
nand ( n25112 , n25110 , n25111 );
not ( n25113 , n12857 );
not ( n25114 , n6948 );
or ( n25115 , n25113 , n25114 );
not ( n25116 , n12857 );
nand ( n25117 , n25116 , n6892 );
nand ( n25118 , n25115 , n25117 );
not ( n25119 , n22921 );
buf ( n25120 , n6425 );
not ( n25121 , n25120 );
not ( n25122 , n25121 );
or ( n25123 , n25119 , n25122 );
not ( n25124 , n22920 );
buf ( n25125 , n25120 );
nand ( n25126 , n25124 , n25125 );
nand ( n25127 , n25123 , n25126 );
buf ( n25128 , n6426 );
buf ( n25129 , n25128 );
and ( n25130 , n25127 , n25129 );
not ( n25131 , n25127 );
not ( n25132 , n25128 );
and ( n25133 , n25131 , n25132 );
nor ( n25134 , n25130 , n25133 );
buf ( n25135 , n6427 );
nand ( n25136 , n7868 , n25135 );
buf ( n25137 , n6428 );
not ( n25138 , n25137 );
and ( n25139 , n25136 , n25138 );
not ( n25140 , n25136 );
buf ( n25141 , n25137 );
and ( n25142 , n25140 , n25141 );
nor ( n25143 , n25139 , n25142 );
xor ( n25144 , n25134 , n25143 );
buf ( n25145 , n6429 );
nand ( n25146 , n7259 , n25145 );
buf ( n25147 , n6430 );
not ( n25148 , n25147 );
and ( n25149 , n25146 , n25148 );
not ( n25150 , n25146 );
buf ( n25151 , n25147 );
and ( n25152 , n25150 , n25151 );
nor ( n25153 , n25149 , n25152 );
xnor ( n25154 , n25144 , n25153 );
buf ( n25155 , n25154 );
not ( n25156 , n25155 );
and ( n25157 , n25118 , n25156 );
not ( n25158 , n25118 );
buf ( n25159 , n25154 );
and ( n25160 , n25158 , n25159 );
nor ( n25161 , n25157 , n25160 );
not ( n25162 , n25161 );
not ( n25163 , n6801 );
not ( n25164 , n14393 );
or ( n25165 , n25163 , n25164 );
not ( n25166 , n6801 );
xor ( n25167 , n14376 , n14385 );
xor ( n25168 , n25167 , n14392 );
nand ( n25169 , n25166 , n25168 );
nand ( n25170 , n25165 , n25169 );
xor ( n25171 , n25170 , n12594 );
not ( n25172 , n25171 );
nand ( n25173 , n25162 , n25172 );
not ( n25174 , n25173 );
buf ( n25175 , n9501 );
not ( n25176 , n25175 );
not ( n25177 , n25176 );
not ( n25178 , n23822 );
or ( n25179 , n25177 , n25178 );
nand ( n25180 , n23826 , n25175 );
nand ( n25181 , n25179 , n25180 );
and ( n25182 , n25181 , n18579 );
not ( n25183 , n25181 );
not ( n25184 , n18579 );
and ( n25185 , n25183 , n25184 );
nor ( n25186 , n25182 , n25185 );
not ( n25187 , n25186 );
not ( n25188 , n25187 );
not ( n25189 , n25188 );
and ( n25190 , n25174 , n25189 );
and ( n25191 , n25173 , n25188 );
nor ( n25192 , n25190 , n25191 );
and ( n25193 , n25112 , n25192 );
not ( n25194 , n25112 );
not ( n25195 , n25192 );
and ( n25196 , n25194 , n25195 );
nor ( n25197 , n25193 , n25196 );
not ( n25198 , n11775 );
not ( n25199 , n23682 );
not ( n25200 , n7314 );
or ( n25201 , n25199 , n25200 );
buf ( n25202 , n11757 );
nand ( n25203 , n25202 , n23678 );
nand ( n25204 , n25201 , n25203 );
not ( n25205 , n25204 );
not ( n25206 , n25205 );
or ( n25207 , n25198 , n25206 );
nand ( n25208 , n16151 , n25204 );
nand ( n25209 , n25207 , n25208 );
not ( n25210 , n15475 );
not ( n25211 , n10077 );
not ( n25212 , n19541 );
or ( n25213 , n25211 , n25212 );
or ( n25214 , n19541 , n10077 );
nand ( n25215 , n25213 , n25214 );
not ( n25216 , n25215 );
or ( n25217 , n25210 , n25216 );
or ( n25218 , n25215 , n15470 );
nand ( n25219 , n25217 , n25218 );
not ( n25220 , n25219 );
nand ( n25221 , n25209 , n25220 );
not ( n25222 , n7126 );
not ( n25223 , n25222 );
not ( n25224 , n19526 );
or ( n25225 , n25223 , n25224 );
not ( n25226 , n19501 );
xor ( n25227 , n19521 , n25226 );
xnor ( n25228 , n25227 , n19491 );
nand ( n25229 , n25228 , n7126 );
nand ( n25230 , n25225 , n25229 );
not ( n25231 , n25230 );
not ( n25232 , n19480 );
or ( n25233 , n25231 , n25232 );
or ( n25234 , n19480 , n25230 );
nand ( n25235 , n25233 , n25234 );
and ( n25236 , n25221 , n25235 );
not ( n25237 , n25221 );
not ( n25238 , n25235 );
and ( n25239 , n25237 , n25238 );
nor ( n25240 , n25236 , n25239 );
not ( n25241 , n25240 );
buf ( n25242 , n11043 );
not ( n25243 , n25242 );
not ( n25244 , n18668 );
or ( n25245 , n25243 , n25244 );
or ( n25246 , n18668 , n25242 );
nand ( n25247 , n25245 , n25246 );
buf ( n25248 , n7756 );
and ( n25249 , n25247 , n25248 );
not ( n25250 , n25247 );
not ( n25251 , n7752 );
not ( n25252 , n25251 );
not ( n25253 , n7742 );
not ( n25254 , n25253 );
or ( n25255 , n25252 , n25254 );
nand ( n25256 , n7742 , n7752 );
nand ( n25257 , n25255 , n25256 );
buf ( n25258 , n25257 );
and ( n25259 , n25250 , n25258 );
nor ( n25260 , n25249 , n25259 );
not ( n25261 , n14121 );
not ( n25262 , n15518 );
or ( n25263 , n25261 , n25262 );
not ( n25264 , n14121 );
nand ( n25265 , n25264 , n15521 );
nand ( n25266 , n25263 , n25265 );
and ( n25267 , n25266 , n15576 );
not ( n25268 , n25266 );
and ( n25269 , n25268 , n15563 );
nor ( n25270 , n25267 , n25269 );
not ( n25271 , n25270 );
nand ( n25272 , n25260 , n25271 );
not ( n25273 , n25272 );
buf ( n25274 , n6431 );
buf ( n25275 , n25274 );
not ( n25276 , n25275 );
buf ( n25277 , n6432 );
not ( n25278 , n25277 );
not ( n25279 , n25278 );
or ( n25280 , n25276 , n25279 );
not ( n25281 , n25274 );
buf ( n25282 , n25277 );
nand ( n25283 , n25281 , n25282 );
nand ( n25284 , n25280 , n25283 );
buf ( n25285 , n6433 );
buf ( n25286 , n25285 );
and ( n25287 , n25284 , n25286 );
not ( n25288 , n25284 );
not ( n25289 , n25285 );
and ( n25290 , n25288 , n25289 );
nor ( n25291 , n25287 , n25290 );
buf ( n25292 , n6434 );
nand ( n25293 , n7014 , n25292 );
buf ( n25294 , n6435 );
not ( n25295 , n25294 );
and ( n25296 , n25293 , n25295 );
not ( n25297 , n25293 );
buf ( n25298 , n25294 );
and ( n25299 , n25297 , n25298 );
nor ( n25300 , n25296 , n25299 );
xor ( n25301 , n25291 , n25300 );
buf ( n25302 , n6436 );
nand ( n25303 , n6558 , n25302 );
buf ( n25304 , n6437 );
not ( n25305 , n25304 );
and ( n25306 , n25303 , n25305 );
not ( n25307 , n25303 );
buf ( n25308 , n25304 );
and ( n25309 , n25307 , n25308 );
nor ( n25310 , n25306 , n25309 );
xnor ( n25311 , n25301 , n25310 );
buf ( n25312 , n25311 );
not ( n25313 , n25312 );
not ( n25314 , n23317 );
not ( n25315 , n23320 );
or ( n25316 , n25314 , n25315 );
or ( n25317 , n23320 , n23317 );
nand ( n25318 , n25316 , n25317 );
not ( n25319 , n25318 );
not ( n25320 , n18115 );
buf ( n25321 , n6438 );
not ( n25322 , n25321 );
not ( n25323 , n25322 );
or ( n25324 , n25320 , n25323 );
not ( n25325 , n18114 );
buf ( n25326 , n25321 );
nand ( n25327 , n25325 , n25326 );
nand ( n25328 , n25324 , n25327 );
buf ( n25329 , n6439 );
not ( n25330 , n25329 );
and ( n25331 , n25328 , n25330 );
not ( n25332 , n25328 );
buf ( n25333 , n25329 );
and ( n25334 , n25332 , n25333 );
nor ( n25335 , n25331 , n25334 );
xor ( n25336 , n25335 , n24788 );
buf ( n25337 , n6440 );
nand ( n25338 , n8223 , n25337 );
buf ( n25339 , n6441 );
not ( n25340 , n25339 );
and ( n25341 , n25338 , n25340 );
not ( n25342 , n25338 );
buf ( n25343 , n25339 );
and ( n25344 , n25342 , n25343 );
nor ( n25345 , n25341 , n25344 );
xnor ( n25346 , n25336 , n25345 );
not ( n25347 , n25346 );
or ( n25348 , n25319 , n25347 );
or ( n25349 , n25318 , n25346 );
nand ( n25350 , n25348 , n25349 );
not ( n25351 , n25350 );
or ( n25352 , n25313 , n25351 );
or ( n25353 , n25350 , n25312 );
nand ( n25354 , n25352 , n25353 );
not ( n25355 , n25354 );
and ( n25356 , n25273 , n25355 );
and ( n25357 , n25272 , n25354 );
nor ( n25358 , n25356 , n25357 );
not ( n25359 , n25358 );
not ( n25360 , n25359 );
or ( n25361 , n25241 , n25360 );
not ( n25362 , n25240 );
nand ( n25363 , n25362 , n25358 );
nand ( n25364 , n25361 , n25363 );
not ( n25365 , n25364 );
and ( n25366 , n25197 , n25365 );
not ( n25367 , n25197 );
and ( n25368 , n25367 , n25364 );
nor ( n25369 , n25366 , n25368 );
buf ( n25370 , n25369 );
and ( n25371 , n25030 , n25370 );
not ( n25372 , n25030 );
and ( n25373 , n25197 , n25364 );
not ( n25374 , n25197 );
and ( n25375 , n25374 , n25365 );
nor ( n25376 , n25373 , n25375 );
buf ( n25377 , n25376 );
and ( n25378 , n25372 , n25377 );
nor ( n25379 , n25371 , n25378 );
nand ( n25380 , n24733 , n25379 );
not ( n25381 , n7143 );
not ( n25382 , n7671 );
not ( n25383 , n7585 );
nand ( n25384 , n25382 , n25383 );
not ( n25385 , n25384 );
not ( n25386 , n22506 );
and ( n25387 , n25385 , n25386 );
and ( n25388 , n25384 , n22506 );
nor ( n25389 , n25387 , n25388 );
not ( n25390 , n25389 );
not ( n25391 , n25390 );
nand ( n25392 , n7757 , n7934 );
not ( n25393 , n25392 );
not ( n25394 , n22424 );
and ( n25395 , n25393 , n25394 );
and ( n25396 , n25392 , n22424 );
nor ( n25397 , n25395 , n25396 );
not ( n25398 , n25397 );
or ( n25399 , n25391 , n25398 );
not ( n25400 , n25397 );
nand ( n25401 , n25400 , n25389 );
nand ( n25402 , n25399 , n25401 );
not ( n25403 , n25402 );
not ( n25404 , n25403 );
not ( n25405 , n22399 );
nand ( n25406 , n7032 , n6851 );
not ( n25407 , n25406 );
or ( n25408 , n25405 , n25407 );
or ( n25409 , n25406 , n22399 );
nand ( n25410 , n25408 , n25409 );
not ( n25411 , n25410 );
nand ( n25412 , n7138 , n6743 );
not ( n25413 , n25412 );
buf ( n25414 , n22290 );
not ( n25415 , n25414 );
not ( n25416 , n25415 );
and ( n25417 , n25413 , n25416 );
and ( n25418 , n25412 , n25415 );
nor ( n25419 , n25417 , n25418 );
not ( n25420 , n25419 );
or ( n25421 , n25411 , n25420 );
or ( n25422 , n25410 , n25419 );
nand ( n25423 , n25421 , n25422 );
not ( n25424 , n7226 );
nand ( n25425 , n25424 , n7417 );
xnor ( n25426 , n25425 , n22321 );
not ( n25427 , n25426 );
and ( n25428 , n25423 , n25427 );
not ( n25429 , n25423 );
and ( n25430 , n25429 , n25426 );
nor ( n25431 , n25428 , n25430 );
not ( n25432 , n25431 );
not ( n25433 , n25432 );
or ( n25434 , n25404 , n25433 );
not ( n25435 , n25432 );
not ( n25436 , n25403 );
nand ( n25437 , n25435 , n25436 );
nand ( n25438 , n25434 , n25437 );
not ( n25439 , n25438 );
or ( n25440 , n25381 , n25439 );
not ( n25441 , n7143 );
and ( n25442 , n25431 , n25402 );
not ( n25443 , n25431 );
and ( n25444 , n25443 , n25403 );
nor ( n25445 , n25442 , n25444 );
nand ( n25446 , n25441 , n25445 );
nand ( n25447 , n25440 , n25446 );
or ( n25448 , n8050 , n8239 );
not ( n25449 , n12555 );
buf ( n25450 , n6442 );
buf ( n25451 , n25450 );
not ( n25452 , n25451 );
buf ( n25453 , n6443 );
not ( n25454 , n25453 );
not ( n25455 , n25454 );
or ( n25456 , n25452 , n25455 );
not ( n25457 , n25450 );
buf ( n25458 , n25453 );
nand ( n25459 , n25457 , n25458 );
nand ( n25460 , n25456 , n25459 );
buf ( n25461 , n6444 );
buf ( n25462 , n25461 );
and ( n25463 , n25460 , n25462 );
not ( n25464 , n25460 );
not ( n25465 , n25461 );
and ( n25466 , n25464 , n25465 );
nor ( n25467 , n25463 , n25466 );
buf ( n25468 , n6445 );
nand ( n25469 , n6502 , n25468 );
buf ( n25470 , n6446 );
not ( n25471 , n25470 );
and ( n25472 , n25469 , n25471 );
not ( n25473 , n25469 );
buf ( n25474 , n25470 );
and ( n25475 , n25473 , n25474 );
nor ( n25476 , n25472 , n25475 );
xor ( n25477 , n25467 , n25476 );
buf ( n25478 , n6447 );
nand ( n25479 , n8455 , n25478 );
buf ( n25480 , n6448 );
not ( n25481 , n25480 );
and ( n25482 , n25479 , n25481 );
not ( n25483 , n25479 );
buf ( n25484 , n25480 );
and ( n25485 , n25483 , n25484 );
nor ( n25486 , n25482 , n25485 );
xnor ( n25487 , n25477 , n25486 );
not ( n25488 , n25487 );
or ( n25489 , n25449 , n25488 );
or ( n25490 , n25487 , n12555 );
nand ( n25491 , n25489 , n25490 );
xor ( n25492 , n21761 , n18454 );
xnor ( n25493 , n25492 , n24734 );
buf ( n25494 , n25493 );
and ( n25495 , n25491 , n25494 );
not ( n25496 , n25491 );
and ( n25497 , n25496 , n21772 );
nor ( n25498 , n25495 , n25497 );
not ( n25499 , n25498 );
and ( n25500 , n25448 , n25499 );
not ( n25501 , n25448 );
and ( n25502 , n25501 , n25498 );
nor ( n25503 , n25500 , n25502 );
not ( n25504 , n25503 );
not ( n25505 , n25504 );
nand ( n25506 , n8319 , n8445 );
not ( n25507 , n17455 );
not ( n25508 , n14056 );
not ( n25509 , n12993 );
or ( n25510 , n25508 , n25509 );
not ( n25511 , n14056 );
nand ( n25512 , n25511 , n13006 );
nand ( n25513 , n25510 , n25512 );
not ( n25514 , n25513 );
and ( n25515 , n25507 , n25514 );
and ( n25516 , n17455 , n25513 );
nor ( n25517 , n25515 , n25516 );
and ( n25518 , n25506 , n25517 );
not ( n25519 , n25506 );
not ( n25520 , n25517 );
and ( n25521 , n25519 , n25520 );
nor ( n25522 , n25518 , n25521 );
not ( n25523 , n25522 );
not ( n25524 , n25523 );
or ( n25525 , n25505 , n25524 );
nand ( n25526 , n25522 , n25503 );
nand ( n25527 , n25525 , n25526 );
nand ( n25528 , n8553 , n8664 );
xor ( n25529 , n18826 , n7129 );
xor ( n25530 , n25529 , n15361 );
not ( n25531 , n25530 );
and ( n25532 , n25528 , n25531 );
not ( n25533 , n25528 );
and ( n25534 , n25533 , n25530 );
nor ( n25535 , n25532 , n25534 );
and ( n25536 , n25527 , n25535 );
not ( n25537 , n25527 );
not ( n25538 , n25535 );
and ( n25539 , n25537 , n25538 );
nor ( n25540 , n25536 , n25539 );
not ( n25541 , n25540 );
not ( n25542 , n25541 );
and ( n25543 , n14931 , n17085 );
not ( n25544 , n14931 );
not ( n25545 , n17085 );
and ( n25546 , n25544 , n25545 );
or ( n25547 , n25543 , n25546 );
not ( n25548 , n7927 );
not ( n25549 , n25548 );
and ( n25550 , n25547 , n25549 );
not ( n25551 , n25547 );
not ( n25552 , n7923 );
and ( n25553 , n25551 , n25552 );
nor ( n25554 , n25550 , n25553 );
not ( n25555 , n25554 );
not ( n25556 , n25555 );
not ( n25557 , n9003 );
nand ( n25558 , n9069 , n25557 );
not ( n25559 , n25558 );
or ( n25560 , n25556 , n25559 );
not ( n25561 , n9003 );
nand ( n25562 , n25561 , n9069 );
or ( n25563 , n25562 , n25555 );
nand ( n25564 , n25560 , n25563 );
not ( n25565 , n25564 );
not ( n25566 , n8763 );
nand ( n25567 , n25566 , n8919 );
not ( n25568 , n25567 );
xor ( n25569 , n20644 , n20410 );
buf ( n25570 , n23126 );
xor ( n25571 , n25569 , n25570 );
not ( n25572 , n25571 );
not ( n25573 , n25572 );
and ( n25574 , n25568 , n25573 );
not ( n25575 , n8918 );
nand ( n25576 , n25575 , n25566 );
and ( n25577 , n25576 , n25572 );
nor ( n25578 , n25574 , n25577 );
not ( n25579 , n25578 );
or ( n25580 , n25565 , n25579 );
or ( n25581 , n25578 , n25564 );
nand ( n25582 , n25580 , n25581 );
not ( n25583 , n25582 );
not ( n25584 , n25583 );
or ( n25585 , n25542 , n25584 );
nand ( n25586 , n25540 , n25582 );
nand ( n25587 , n25585 , n25586 );
buf ( n25588 , n25587 );
not ( n25589 , n25588 );
and ( n25590 , n25447 , n25589 );
not ( n25591 , n25447 );
and ( n25592 , n25591 , n25588 );
nor ( n25593 , n25590 , n25592 );
not ( n25594 , n17150 );
nand ( n25595 , n25594 , n11110 );
not ( n25596 , n25595 );
not ( n25597 , n17241 );
not ( n25598 , n25597 );
and ( n25599 , n25596 , n25598 );
nand ( n25600 , n25594 , n11110 );
and ( n25601 , n25600 , n25597 );
nor ( n25602 , n25599 , n25601 );
not ( n25603 , n25602 );
not ( n25604 , n17377 );
or ( n25605 , n25603 , n25604 );
not ( n25606 , n25602 );
not ( n25607 , n17372 );
not ( n25608 , n17285 );
and ( n25609 , n25607 , n25608 );
and ( n25610 , n17372 , n17285 );
nor ( n25611 , n25609 , n25610 );
nand ( n25612 , n25606 , n25611 );
nand ( n25613 , n25605 , n25612 );
buf ( n25614 , n17796 );
and ( n25615 , n25613 , n25614 );
not ( n25616 , n25613 );
not ( n25617 , n25614 );
and ( n25618 , n25616 , n25617 );
nor ( n25619 , n25615 , n25618 );
nand ( n25620 , n25593 , n25619 );
or ( n25621 , n25380 , n25620 );
not ( n25622 , n25619 );
not ( n25623 , n25379 );
or ( n25624 , n25622 , n25623 );
buf ( n25625 , n15325 );
nor ( n25626 , n25593 , n25625 );
nand ( n25627 , n25624 , n25626 );
buf ( n25628 , n13353 );
nand ( n25629 , n25628 , n7244 );
nand ( n25630 , n25621 , n25627 , n25629 );
buf ( n25631 , n25630 );
buf ( n25632 , n25631 );
not ( n25633 , n10362 );
not ( n25634 , n11121 );
or ( n25635 , n25633 , n25634 );
or ( n25636 , n11121 , n10362 );
nand ( n25637 , n25635 , n25636 );
and ( n25638 , n25637 , n11155 );
not ( n25639 , n25637 );
and ( n25640 , n25639 , n11156 );
nor ( n25641 , n25638 , n25640 );
not ( n25642 , n25641 );
not ( n25643 , n20080 );
nand ( n25644 , n25642 , n25643 );
and ( n25645 , n25644 , n19998 );
not ( n25646 , n25644 );
not ( n25647 , n19998 );
and ( n25648 , n25646 , n25647 );
nor ( n25649 , n25645 , n25648 );
not ( n25650 , n25649 );
not ( n25651 , n20536 );
or ( n25652 , n25650 , n25651 );
not ( n25653 , n25649 );
nand ( n25654 , n25653 , n20544 );
nand ( n25655 , n25652 , n25654 );
and ( n25656 , n25655 , n20966 );
not ( n25657 , n25655 );
and ( n25658 , n25657 , n20952 );
nor ( n25659 , n25656 , n25658 );
buf ( n25660 , n13345 );
not ( n25661 , n25660 );
nand ( n25662 , n25659 , n25661 );
not ( n25663 , n12180 );
not ( n25664 , n20631 );
or ( n25665 , n25663 , n25664 );
nand ( n25666 , n20628 , n12183 );
nand ( n25667 , n25665 , n25666 );
and ( n25668 , n25667 , n19101 );
not ( n25669 , n25667 );
and ( n25670 , n25669 , n9695 );
nor ( n25671 , n25668 , n25670 );
not ( n25672 , n25671 );
not ( n25673 , n14883 );
not ( n25674 , n17040 );
or ( n25675 , n25673 , n25674 );
nand ( n25676 , n17043 , n14917 );
nand ( n25677 , n25675 , n25676 );
not ( n25678 , n25677 );
not ( n25679 , n17086 );
and ( n25680 , n25678 , n25679 );
not ( n25681 , n17084 );
buf ( n25682 , n25681 );
not ( n25683 , n25682 );
not ( n25684 , n25683 );
and ( n25685 , n25677 , n25684 );
nor ( n25686 , n25680 , n25685 );
not ( n25687 , n25686 );
nand ( n25688 , n25672 , n25687 );
not ( n25689 , n25688 );
xor ( n25690 , n16029 , n14152 );
xnor ( n25691 , n25690 , n14175 );
not ( n25692 , n25691 );
not ( n25693 , n25692 );
or ( n25694 , n25689 , n25693 );
or ( n25695 , n25692 , n25688 );
nand ( n25696 , n25694 , n25695 );
not ( n25697 , n25696 );
not ( n25698 , n14749 );
not ( n25699 , n14727 );
and ( n25700 , n25698 , n25699 );
and ( n25701 , n14749 , n14727 );
nor ( n25702 , n25700 , n25701 );
not ( n25703 , n25702 );
not ( n25704 , n16665 );
not ( n25705 , n16677 );
xor ( n25706 , n25704 , n25705 );
xnor ( n25707 , n25706 , n16680 );
and ( n25708 , n9359 , n25707 );
not ( n25709 , n9359 );
and ( n25710 , n25709 , n16682 );
nor ( n25711 , n25708 , n25710 );
not ( n25712 , n25711 );
and ( n25713 , n25703 , n25712 );
and ( n25714 , n14755 , n25711 );
nor ( n25715 , n25713 , n25714 );
not ( n25716 , n25715 );
not ( n25717 , n25716 );
not ( n25718 , n8568 );
not ( n25719 , n10637 );
not ( n25720 , n13906 );
or ( n25721 , n25719 , n25720 );
nand ( n25722 , n13905 , n10633 );
nand ( n25723 , n25721 , n25722 );
not ( n25724 , n25723 );
and ( n25725 , n25718 , n25724 );
not ( n25726 , n7802 );
and ( n25727 , n25726 , n25723 );
nor ( n25728 , n25725 , n25727 );
not ( n25729 , n15889 );
not ( n25730 , n10036 );
or ( n25731 , n25729 , n25730 );
not ( n25732 , n15889 );
nand ( n25733 , n25732 , n8977 );
nand ( n25734 , n25731 , n25733 );
and ( n25735 , n25734 , n8986 );
not ( n25736 , n25734 );
and ( n25737 , n25736 , n7540 );
nor ( n25738 , n25735 , n25737 );
nand ( n25739 , n25728 , n25738 );
not ( n25740 , n25739 );
or ( n25741 , n25717 , n25740 );
or ( n25742 , n25739 , n25716 );
nand ( n25743 , n25741 , n25742 );
not ( n25744 , n25743 );
and ( n25745 , n14284 , n12341 );
not ( n25746 , n14284 );
and ( n25747 , n25746 , n13294 );
nor ( n25748 , n25745 , n25747 );
xnor ( n25749 , n12376 , n25748 );
not ( n25750 , n19304 );
not ( n25751 , n15291 );
or ( n25752 , n25750 , n25751 );
not ( n25753 , n19304 );
nand ( n25754 , n25753 , n23723 );
nand ( n25755 , n25752 , n25754 );
and ( n25756 , n25755 , n15298 );
not ( n25757 , n25755 );
and ( n25758 , n25757 , n14220 );
nor ( n25759 , n25756 , n25758 );
not ( n25760 , n25759 );
nand ( n25761 , n25749 , n25760 );
not ( n25762 , n25761 );
not ( n25763 , n15533 );
not ( n25764 , n9136 );
not ( n25765 , n25764 );
or ( n25766 , n25763 , n25765 );
not ( n25767 , n9136 );
or ( n25768 , n25767 , n15533 );
nand ( n25769 , n25766 , n25768 );
and ( n25770 , n25769 , n9184 );
not ( n25771 , n25769 );
not ( n25772 , n9181 );
not ( n25773 , n25772 );
and ( n25774 , n25771 , n25773 );
nor ( n25775 , n25770 , n25774 );
not ( n25776 , n25775 );
not ( n25777 , n25776 );
not ( n25778 , n25777 );
and ( n25779 , n25762 , n25778 );
and ( n25780 , n25761 , n25777 );
nor ( n25781 , n25779 , n25780 );
not ( n25782 , n25781 );
or ( n25783 , n25744 , n25782 );
or ( n25784 , n25781 , n25743 );
nand ( n25785 , n25783 , n25784 );
nand ( n25786 , n25691 , n25671 );
not ( n25787 , n10106 );
not ( n25788 , n24961 );
or ( n25789 , n25787 , n25788 );
not ( n25790 , n10106 );
not ( n25791 , n24961 );
nand ( n25792 , n25790 , n25791 );
nand ( n25793 , n25789 , n25792 );
and ( n25794 , n25793 , n22821 );
not ( n25795 , n25793 );
and ( n25796 , n25795 , n22817 );
nor ( n25797 , n25794 , n25796 );
not ( n25798 , n25797 );
and ( n25799 , n25786 , n25798 );
not ( n25800 , n25786 );
and ( n25801 , n25800 , n25797 );
nor ( n25802 , n25799 , n25801 );
not ( n25803 , n25802 );
and ( n25804 , n25785 , n25803 );
not ( n25805 , n25785 );
and ( n25806 , n25805 , n25802 );
nor ( n25807 , n25804 , n25806 );
not ( n25808 , n25807 );
not ( n25809 , n12263 );
buf ( n25810 , n20782 );
not ( n25811 , n25810 );
or ( n25812 , n25809 , n25811 );
or ( n25813 , n22586 , n12263 );
nand ( n25814 , n25812 , n25813 );
buf ( n25815 , n6977 );
and ( n25816 , n25814 , n25815 );
not ( n25817 , n25814 );
and ( n25818 , n25817 , n18730 );
nor ( n25819 , n25816 , n25818 );
not ( n25820 , n7589 );
not ( n25821 , n22658 );
or ( n25822 , n25820 , n25821 );
or ( n25823 , n22658 , n7589 );
nand ( n25824 , n25822 , n25823 );
not ( n25825 , n16453 );
not ( n25826 , n25825 );
not ( n25827 , n25826 );
and ( n25828 , n25824 , n25827 );
not ( n25829 , n25824 );
buf ( n25830 , n21864 );
and ( n25831 , n25829 , n25830 );
nor ( n25832 , n25828 , n25831 );
nand ( n25833 , n25819 , n25832 );
not ( n25834 , n25833 );
not ( n25835 , n9015 );
not ( n25836 , n10227 );
or ( n25837 , n25835 , n25836 );
buf ( n25838 , n12933 );
nand ( n25839 , n25838 , n9011 );
nand ( n25840 , n25837 , n25839 );
not ( n25841 , n12936 );
and ( n25842 , n25840 , n25841 );
not ( n25843 , n25840 );
and ( n25844 , n25843 , n12936 );
nor ( n25845 , n25842 , n25844 );
not ( n25846 , n25845 );
and ( n25847 , n25834 , n25846 );
and ( n25848 , n25833 , n25845 );
nor ( n25849 , n25847 , n25848 );
not ( n25850 , n25849 );
buf ( n25851 , n24381 );
xor ( n25852 , n18182 , n25851 );
not ( n25853 , n24681 );
xnor ( n25854 , n25852 , n25853 );
not ( n25855 , n25854 );
not ( n25856 , n7431 );
buf ( n25857 , n6449 );
buf ( n25858 , n25857 );
not ( n25859 , n25858 );
not ( n25860 , n10750 );
or ( n25861 , n25859 , n25860 );
not ( n25862 , n25857 );
nand ( n25863 , n25862 , n10705 );
nand ( n25864 , n25861 , n25863 );
buf ( n25865 , n6450 );
not ( n25866 , n25865 );
and ( n25867 , n25864 , n25866 );
not ( n25868 , n25864 );
buf ( n25869 , n25865 );
and ( n25870 , n25868 , n25869 );
nor ( n25871 , n25867 , n25870 );
xor ( n25872 , n25871 , n19988 );
buf ( n25873 , n6451 );
nand ( n25874 , n7344 , n25873 );
buf ( n25875 , n6452 );
buf ( n25876 , n25875 );
and ( n25877 , n25874 , n25876 );
not ( n25878 , n25874 );
not ( n25879 , n25875 );
and ( n25880 , n25878 , n25879 );
nor ( n25881 , n25877 , n25880 );
not ( n25882 , n25881 );
xnor ( n25883 , n25872 , n25882 );
buf ( n25884 , n25883 );
not ( n25885 , n25884 );
or ( n25886 , n25856 , n25885 );
not ( n25887 , n25883 );
not ( n25888 , n25887 );
or ( n25889 , n25888 , n7431 );
nand ( n25890 , n25886 , n25889 );
buf ( n25891 , n11614 );
and ( n25892 , n25890 , n25891 );
not ( n25893 , n25890 );
not ( n25894 , n25891 );
and ( n25895 , n25893 , n25894 );
nor ( n25896 , n25892 , n25895 );
nand ( n25897 , n25855 , n25896 );
not ( n25898 , n13822 );
not ( n25899 , n20198 );
or ( n25900 , n25898 , n25899 );
buf ( n25901 , n20202 );
nand ( n25902 , n25901 , n13818 );
nand ( n25903 , n25900 , n25902 );
not ( n25904 , n22414 );
and ( n25905 , n25903 , n25904 );
not ( n25906 , n25903 );
and ( n25907 , n25906 , n22414 );
nor ( n25908 , n25905 , n25907 );
and ( n25909 , n25897 , n25908 );
not ( n25910 , n25897 );
not ( n25911 , n25908 );
and ( n25912 , n25910 , n25911 );
nor ( n25913 , n25909 , n25912 );
not ( n25914 , n25913 );
or ( n25915 , n25850 , n25914 );
or ( n25916 , n25913 , n25849 );
nand ( n25917 , n25915 , n25916 );
not ( n25918 , n25917 );
and ( n25919 , n25808 , n25918 );
not ( n25920 , n25808 );
and ( n25921 , n25920 , n25917 );
nor ( n25922 , n25919 , n25921 );
not ( n25923 , n25922 );
or ( n25924 , n25697 , n25923 );
not ( n25925 , n25696 );
not ( n25926 , n25918 );
not ( n25927 , n25807 );
not ( n25928 , n25927 );
or ( n25929 , n25926 , n25928 );
nand ( n25930 , n25807 , n25917 );
nand ( n25931 , n25929 , n25930 );
nand ( n25932 , n25925 , n25931 );
nand ( n25933 , n25924 , n25932 );
buf ( n25934 , n6453 );
nand ( n25935 , n7563 , n25934 );
buf ( n25936 , n6454 );
buf ( n25937 , n25936 );
and ( n25938 , n25935 , n25937 );
not ( n25939 , n25935 );
not ( n25940 , n25936 );
and ( n25941 , n25939 , n25940 );
nor ( n25942 , n25938 , n25941 );
buf ( n25943 , n25942 );
xor ( n25944 , n25943 , n14624 );
xor ( n25945 , n25944 , n25888 );
buf ( n25946 , n12195 );
not ( n25947 , n25946 );
not ( n25948 , n20628 );
or ( n25949 , n25947 , n25948 );
or ( n25950 , n20628 , n25946 );
nand ( n25951 , n25949 , n25950 );
not ( n25952 , n25951 );
not ( n25953 , n9695 );
and ( n25954 , n25952 , n25953 );
buf ( n25955 , n19102 );
and ( n25956 , n25951 , n25955 );
nor ( n25957 , n25954 , n25956 );
nand ( n25958 , n25945 , n25957 );
not ( n25959 , n8697 );
not ( n25960 , n10849 );
or ( n25961 , n25959 , n25960 );
or ( n25962 , n10849 , n8697 );
nand ( n25963 , n25961 , n25962 );
buf ( n25964 , n16910 );
not ( n25965 , n25964 );
and ( n25966 , n25963 , n25965 );
not ( n25967 , n25963 );
and ( n25968 , n25967 , n25964 );
nor ( n25969 , n25966 , n25968 );
xnor ( n25970 , n25958 , n25969 );
not ( n25971 , n25970 );
buf ( n25972 , n14645 );
and ( n25973 , n14649 , n25972 );
not ( n25974 , n14649 );
and ( n25975 , n25974 , n14646 );
nor ( n25976 , n25973 , n25975 );
xor ( n25977 , n25976 , n11957 );
not ( n25978 , n25977 );
not ( n25979 , n22100 );
and ( n25980 , n25978 , n25979 );
not ( n25981 , n22100 );
not ( n25982 , n25981 );
and ( n25983 , n25977 , n25982 );
nor ( n25984 , n25980 , n25983 );
not ( n25985 , n25984 );
not ( n25986 , n25985 );
buf ( n25987 , n19541 );
xor ( n25988 , n23983 , n25987 );
xnor ( n25989 , n25988 , n20464 );
nand ( n25990 , n25986 , n25989 );
not ( n25991 , n25990 );
not ( n25992 , n11755 );
not ( n25993 , n25992 );
not ( n25994 , n23686 );
not ( n25995 , n7314 );
or ( n25996 , n25994 , n25995 );
not ( n25997 , n23686 );
nand ( n25998 , n25997 , n25202 );
nand ( n25999 , n25996 , n25998 );
not ( n26000 , n25999 );
or ( n26001 , n25993 , n26000 );
or ( n26002 , n25992 , n25999 );
nand ( n26003 , n26001 , n26002 );
not ( n26004 , n26003 );
and ( n26005 , n25991 , n26004 );
not ( n26006 , n25985 );
nand ( n26007 , n26006 , n25989 );
and ( n26008 , n26007 , n26003 );
nor ( n26009 , n26005 , n26008 );
not ( n26010 , n26009 );
or ( n26011 , n25971 , n26010 );
or ( n26012 , n26009 , n25970 );
nand ( n26013 , n26011 , n26012 );
not ( n26014 , n26013 );
buf ( n26015 , n7353 );
not ( n26016 , n26015 );
not ( n26017 , n18237 );
or ( n26018 , n26016 , n26017 );
or ( n26019 , n18237 , n26015 );
nand ( n26020 , n26018 , n26019 );
xnor ( n26021 , n26020 , n18261 );
not ( n26022 , n26021 );
not ( n26023 , n23917 );
not ( n26024 , n12030 );
not ( n26025 , n16913 );
or ( n26026 , n26024 , n26025 );
or ( n26027 , n16913 , n12030 );
nand ( n26028 , n26026 , n26027 );
not ( n26029 , n26028 );
or ( n26030 , n26023 , n26029 );
not ( n26031 , n23916 );
not ( n26032 , n26031 );
or ( n26033 , n26028 , n26032 );
nand ( n26034 , n26030 , n26033 );
nand ( n26035 , n26022 , n26034 );
not ( n26036 , n26035 );
not ( n26037 , n17039 );
not ( n26038 , n14903 );
and ( n26039 , n26037 , n26038 );
and ( n26040 , n17039 , n14903 );
nor ( n26041 , n26039 , n26040 );
and ( n26042 , n26041 , n25682 );
not ( n26043 , n26041 );
and ( n26044 , n26043 , n25545 );
nor ( n26045 , n26042 , n26044 );
not ( n26046 , n26045 );
and ( n26047 , n26036 , n26046 );
and ( n26048 , n26035 , n26045 );
nor ( n26049 , n26047 , n26048 );
not ( n26050 , n26049 );
not ( n26051 , n25815 );
not ( n26052 , n20776 );
not ( n26053 , n12284 );
and ( n26054 , n26052 , n26053 );
not ( n26055 , n12285 );
and ( n26056 , n20776 , n26055 );
nor ( n26057 , n26054 , n26056 );
not ( n26058 , n26057 );
or ( n26059 , n26051 , n26058 );
or ( n26060 , n26057 , n25815 );
nand ( n26061 , n26059 , n26060 );
not ( n26062 , n18377 );
not ( n26063 , n20517 );
or ( n26064 , n26062 , n26063 );
or ( n26065 , n20517 , n18377 );
nand ( n26066 , n26064 , n26065 );
xor ( n26067 , n26066 , n23180 );
nand ( n26068 , n26061 , n26067 );
not ( n26069 , n12787 );
not ( n26070 , n9374 );
or ( n26071 , n26069 , n26070 );
not ( n26072 , n12787 );
nand ( n26073 , n26072 , n9373 );
nand ( n26074 , n26071 , n26073 );
and ( n26075 , n26074 , n22803 );
not ( n26076 , n26074 );
and ( n26077 , n26076 , n22802 );
nor ( n26078 , n26075 , n26077 );
and ( n26079 , n26068 , n26078 );
not ( n26080 , n26068 );
not ( n26081 , n26078 );
and ( n26082 , n26080 , n26081 );
nor ( n26083 , n26079 , n26082 );
not ( n26084 , n26083 );
or ( n26085 , n26050 , n26084 );
or ( n26086 , n26083 , n26049 );
nand ( n26087 , n26085 , n26086 );
not ( n26088 , n25726 );
not ( n26089 , n12650 );
not ( n26090 , n26089 );
not ( n26091 , n19874 );
or ( n26092 , n26090 , n26091 );
or ( n26093 , n19874 , n26089 );
nand ( n26094 , n26092 , n26093 );
not ( n26095 , n26094 );
and ( n26096 , n26088 , n26095 );
and ( n26097 , n8568 , n26094 );
nor ( n26098 , n26096 , n26097 );
not ( n26099 , n26098 );
buf ( n26100 , n20069 );
and ( n26101 , n26100 , n17358 );
not ( n26102 , n26100 );
and ( n26103 , n26102 , n12206 );
nor ( n26104 , n26101 , n26103 );
not ( n26105 , n26104 );
not ( n26106 , n26105 );
not ( n26107 , n17361 );
or ( n26108 , n26106 , n26107 );
nand ( n26109 , n12236 , n26104 );
nand ( n26110 , n26108 , n26109 );
not ( n26111 , n26110 );
nand ( n26112 , n26099 , n26111 );
not ( n26113 , n26112 );
buf ( n26114 , n17864 );
xor ( n26115 , n26114 , n24471 );
xnor ( n26116 , n26115 , n24435 );
not ( n26117 , n26116 );
and ( n26118 , n26113 , n26117 );
and ( n26119 , n26112 , n26116 );
nor ( n26120 , n26118 , n26119 );
and ( n26121 , n26087 , n26120 );
not ( n26122 , n26087 );
not ( n26123 , n26120 );
and ( n26124 , n26122 , n26123 );
nor ( n26125 , n26121 , n26124 );
not ( n26126 , n26125 );
or ( n26127 , n26014 , n26126 );
or ( n26128 , n26013 , n26125 );
nand ( n26129 , n26127 , n26128 );
buf ( n26130 , n26129 );
not ( n26131 , n26130 );
not ( n26132 , n26131 );
not ( n26133 , n26132 );
and ( n26134 , n25933 , n26133 );
not ( n26135 , n25933 );
not ( n26136 , n26130 );
not ( n26137 , n26136 );
and ( n26138 , n26135 , n26137 );
nor ( n26139 , n26134 , n26138 );
not ( n26140 , n21587 );
not ( n26141 , n6843 );
not ( n26142 , n26141 );
not ( n26143 , n25168 );
or ( n26144 , n26142 , n26143 );
nand ( n26145 , n14393 , n6843 );
nand ( n26146 , n26144 , n26145 );
not ( n26147 , n26146 );
or ( n26148 , n26140 , n26147 );
or ( n26149 , n26146 , n12594 );
nand ( n26150 , n26148 , n26149 );
not ( n26151 , n26150 );
not ( n26152 , n22656 );
not ( n26153 , n14224 );
or ( n26154 , n26152 , n26153 );
not ( n26155 , n22656 );
nand ( n26156 , n26155 , n14220 );
nand ( n26157 , n26154 , n26156 );
and ( n26158 , n26157 , n14268 );
not ( n26159 , n26157 );
and ( n26160 , n26159 , n14272 );
nor ( n26161 , n26158 , n26160 );
not ( n26162 , n26161 );
nand ( n26163 , n26151 , n26162 );
xor ( n26164 , n19454 , n13537 );
xnor ( n26165 , n26164 , n17614 );
buf ( n26166 , n26165 );
xor ( n26167 , n26163 , n26166 );
not ( n26168 , n26167 );
not ( n26169 , n26168 );
not ( n26170 , n14993 );
not ( n26171 , n12102 );
not ( n26172 , n21983 );
or ( n26173 , n26171 , n26172 );
nand ( n26174 , n21988 , n12105 );
nand ( n26175 , n26173 , n26174 );
not ( n26176 , n26175 );
or ( n26177 , n26170 , n26176 );
or ( n26178 , n26175 , n14993 );
nand ( n26179 , n26177 , n26178 );
not ( n26180 , n26179 );
not ( n26181 , n17083 );
not ( n26182 , n18378 );
or ( n26183 , n26181 , n26182 );
or ( n26184 , n18372 , n17083 );
nand ( n26185 , n26183 , n26184 );
buf ( n26186 , n19773 );
and ( n26187 , n26185 , n26186 );
not ( n26188 , n26185 );
and ( n26189 , n26188 , n10271 );
or ( n26190 , n26187 , n26189 );
nand ( n26191 , n26180 , n26190 );
not ( n26192 , n26191 );
not ( n26193 , n17824 );
not ( n26194 , n24435 );
or ( n26195 , n26193 , n26194 );
or ( n26196 , n24435 , n17824 );
nand ( n26197 , n26195 , n26196 );
buf ( n26198 , n6455 );
buf ( n26199 , n26198 );
not ( n26200 , n26199 );
not ( n26201 , n18041 );
not ( n26202 , n26201 );
or ( n26203 , n26200 , n26202 );
not ( n26204 , n26198 );
nand ( n26205 , n26204 , n18042 );
nand ( n26206 , n26203 , n26205 );
buf ( n26207 , n6456 );
buf ( n26208 , n26207 );
and ( n26209 , n26206 , n26208 );
not ( n26210 , n26206 );
not ( n26211 , n26207 );
and ( n26212 , n26210 , n26211 );
nor ( n26213 , n26209 , n26212 );
buf ( n26214 , n6457 );
nand ( n26215 , n6871 , n26214 );
buf ( n26216 , n6458 );
buf ( n26217 , n26216 );
and ( n26218 , n26215 , n26217 );
not ( n26219 , n26215 );
not ( n26220 , n26216 );
and ( n26221 , n26219 , n26220 );
nor ( n26222 , n26218 , n26221 );
xor ( n26223 , n26213 , n26222 );
xnor ( n26224 , n26223 , n22730 );
buf ( n26225 , n26224 );
not ( n26226 , n26225 );
and ( n26227 , n26197 , n26226 );
not ( n26228 , n26197 );
and ( n26229 , n26228 , n26225 );
nor ( n26230 , n26227 , n26229 );
not ( n26231 , n26230 );
not ( n26232 , n26231 );
and ( n26233 , n26192 , n26232 );
and ( n26234 , n26191 , n26231 );
nor ( n26235 , n26233 , n26234 );
not ( n26236 , n26235 );
nand ( n26237 , n26165 , n26150 );
not ( n26238 , n18730 );
not ( n26239 , n12256 );
not ( n26240 , n20782 );
or ( n26241 , n26239 , n26240 );
nand ( n26242 , n20776 , n12252 );
nand ( n26243 , n26241 , n26242 );
not ( n26244 , n26243 );
or ( n26245 , n26238 , n26244 );
not ( n26246 , n26243 );
nand ( n26247 , n26246 , n25815 );
nand ( n26248 , n26245 , n26247 );
not ( n26249 , n26248 );
and ( n26250 , n26237 , n26249 );
not ( n26251 , n26237 );
and ( n26252 , n26251 , n26248 );
nor ( n26253 , n26250 , n26252 );
not ( n26254 , n26253 );
or ( n26255 , n26236 , n26254 );
or ( n26256 , n26253 , n26235 );
nand ( n26257 , n26255 , n26256 );
not ( n26258 , n15662 );
not ( n26259 , n23973 );
xor ( n26260 , n23964 , n26259 );
xnor ( n26261 , n26260 , n23983 );
buf ( n26262 , n26261 );
not ( n26263 , n26262 );
or ( n26264 , n26258 , n26263 );
buf ( n26265 , n23984 );
buf ( n26266 , n26265 );
nand ( n26267 , n26266 , n15659 );
nand ( n26268 , n26264 , n26267 );
buf ( n26269 , n23991 );
not ( n26270 , n26269 );
and ( n26271 , n26268 , n26270 );
not ( n26272 , n26268 );
and ( n26273 , n26272 , n26269 );
nor ( n26274 , n26271 , n26273 );
not ( n26275 , n26274 );
not ( n26276 , n7136 );
not ( n26277 , n24754 );
not ( n26278 , n7127 );
not ( n26279 , n26278 );
or ( n26280 , n26277 , n26279 );
not ( n26281 , n24754 );
nand ( n26282 , n26281 , n7128 );
nand ( n26283 , n26280 , n26282 );
not ( n26284 , n26283 );
and ( n26285 , n26276 , n26284 );
and ( n26286 , n7136 , n26283 );
nor ( n26287 , n26285 , n26286 );
not ( n26288 , n26287 );
nand ( n26289 , n26275 , n26288 );
not ( n26290 , n8097 );
not ( n26291 , n11108 );
or ( n26292 , n26290 , n26291 );
or ( n26293 , n6741 , n8097 );
nand ( n26294 , n26292 , n26293 );
and ( n26295 , n26294 , n24315 );
not ( n26296 , n26294 );
and ( n26297 , n26296 , n24312 );
nor ( n26298 , n26295 , n26297 );
buf ( n26299 , n26298 );
xnor ( n26300 , n26289 , n26299 );
xnor ( n26301 , n26257 , n26300 );
buf ( n26302 , n24494 );
not ( n26303 , n26302 );
buf ( n26304 , n11672 );
not ( n26305 , n26304 );
or ( n26306 , n26303 , n26305 );
nand ( n26307 , n20232 , n24495 );
nand ( n26308 , n26306 , n26307 );
xor ( n26309 , n11719 , n20107 );
buf ( n26310 , n11697 );
xnor ( n26311 , n26309 , n26310 );
buf ( n26312 , n26311 );
buf ( n26313 , n26312 );
and ( n26314 , n26308 , n26313 );
not ( n26315 , n26308 );
buf ( n26316 , n11727 );
and ( n26317 , n26315 , n26316 );
nor ( n26318 , n26314 , n26317 );
not ( n26319 , n26318 );
xor ( n26320 , n25129 , n17676 );
buf ( n26321 , n22938 );
xnor ( n26322 , n26320 , n26321 );
not ( n26323 , n26322 );
not ( n26324 , n12590 );
not ( n26325 , n25487 );
not ( n26326 , n26325 );
or ( n26327 , n26324 , n26326 );
or ( n26328 , n26325 , n12590 );
nand ( n26329 , n26327 , n26328 );
and ( n26330 , n26329 , n25494 );
not ( n26331 , n26329 );
buf ( n26332 , n21772 );
and ( n26333 , n26331 , n26332 );
nor ( n26334 , n26330 , n26333 );
not ( n26335 , n26334 );
nand ( n26336 , n26323 , n26335 );
not ( n26337 , n26336 );
or ( n26338 , n26319 , n26337 );
not ( n26339 , n26335 );
not ( n26340 , n26339 );
nand ( n26341 , n26340 , n26323 );
or ( n26342 , n26341 , n26318 );
nand ( n26343 , n26338 , n26342 );
not ( n26344 , n26343 );
not ( n26345 , n11246 );
not ( n26346 , n20576 );
or ( n26347 , n26345 , n26346 );
nand ( n26348 , n20575 , n11249 );
nand ( n26349 , n26347 , n26348 );
not ( n26350 , n26349 );
not ( n26351 , n14692 );
and ( n26352 , n26350 , n26351 );
and ( n26353 , n14692 , n26349 );
nor ( n26354 , n26352 , n26353 );
buf ( n26355 , n15872 );
not ( n26356 , n15868 );
and ( n26357 , n26355 , n26356 );
not ( n26358 , n26355 );
and ( n26359 , n26358 , n15869 );
or ( n26360 , n26357 , n26359 );
not ( n26361 , n26360 );
not ( n26362 , n8986 );
or ( n26363 , n26361 , n26362 );
or ( n26364 , n8986 , n26360 );
nand ( n26365 , n26363 , n26364 );
and ( n26366 , n26365 , n7583 );
not ( n26367 , n26365 );
and ( n26368 , n26367 , n7580 );
nor ( n26369 , n26366 , n26368 );
nand ( n26370 , n26354 , n26369 );
not ( n26371 , n26370 );
not ( n26372 , n13615 );
buf ( n26373 , n21883 );
not ( n26374 , n26373 );
or ( n26375 , n26372 , n26374 );
nand ( n26376 , n24767 , n13611 );
nand ( n26377 , n26375 , n26376 );
not ( n26378 , n21892 );
not ( n26379 , n26378 );
xor ( n26380 , n26377 , n26379 );
not ( n26381 , n26380 );
and ( n26382 , n26371 , n26381 );
and ( n26383 , n26370 , n26380 );
nor ( n26384 , n26382 , n26383 );
not ( n26385 , n26384 );
and ( n26386 , n26344 , n26385 );
and ( n26387 , n26343 , n26384 );
nor ( n26388 , n26386 , n26387 );
and ( n26389 , n26301 , n26388 );
not ( n26390 , n26301 );
not ( n26391 , n26388 );
and ( n26392 , n26390 , n26391 );
nor ( n26393 , n26389 , n26392 );
not ( n26394 , n26393 );
or ( n26395 , n26169 , n26394 );
not ( n26396 , n26168 );
and ( n26397 , n26301 , n26391 );
not ( n26398 , n26301 );
and ( n26399 , n26398 , n26388 );
nor ( n26400 , n26397 , n26399 );
nand ( n26401 , n26396 , n26400 );
nand ( n26402 , n26395 , n26401 );
not ( n26403 , n16814 );
buf ( n26404 , n15905 );
not ( n26405 , n26404 );
not ( n26406 , n26405 );
or ( n26407 , n26403 , n26406 );
not ( n26408 , n26404 );
or ( n26409 , n26408 , n16814 );
nand ( n26410 , n26407 , n26409 );
not ( n26411 , n26410 );
not ( n26412 , n20520 );
not ( n26413 , n26412 );
and ( n26414 , n26411 , n26413 );
and ( n26415 , n26410 , n20522 );
nor ( n26416 , n26414 , n26415 );
not ( n26417 , n26416 );
not ( n26418 , n16083 );
not ( n26419 , n14152 );
or ( n26420 , n26418 , n26419 );
or ( n26421 , n14152 , n16083 );
nand ( n26422 , n26420 , n26421 );
and ( n26423 , n26422 , n20232 );
not ( n26424 , n26422 );
buf ( n26425 , n26304 );
and ( n26426 , n26424 , n26425 );
nor ( n26427 , n26423 , n26426 );
not ( n26428 , n26427 );
nand ( n26429 , n26417 , n26428 );
not ( n26430 , n26429 );
not ( n26431 , n15684 );
not ( n26432 , n26262 );
or ( n26433 , n26431 , n26432 );
not ( n26434 , n15684 );
nand ( n26435 , n26434 , n26265 );
nand ( n26436 , n26433 , n26435 );
and ( n26437 , n26436 , n26270 );
not ( n26438 , n26436 );
and ( n26439 , n26438 , n26269 );
nor ( n26440 , n26437 , n26439 );
not ( n26441 , n26440 );
and ( n26442 , n26430 , n26441 );
and ( n26443 , n26429 , n26440 );
nor ( n26444 , n26442 , n26443 );
not ( n26445 , n26444 );
not ( n26446 , n26445 );
not ( n26447 , n13718 );
not ( n26448 , n7450 );
buf ( n26449 , n14781 );
nor ( n26450 , n26448 , n26449 );
not ( n26451 , n26450 );
not ( n26452 , n7450 );
nand ( n26453 , n26449 , n26452 );
nand ( n26454 , n26451 , n26453 );
not ( n26455 , n26454 );
or ( n26456 , n26447 , n26455 );
or ( n26457 , n26454 , n7495 );
nand ( n26458 , n26456 , n26457 );
not ( n26459 , n26458 );
not ( n26460 , n17515 );
not ( n26461 , n20338 );
or ( n26462 , n26460 , n26461 );
nand ( n26463 , n20341 , n17511 );
nand ( n26464 , n26462 , n26463 );
and ( n26465 , n26464 , n20344 );
not ( n26466 , n26464 );
and ( n26467 , n26466 , n20345 );
nor ( n26468 , n26465 , n26467 );
not ( n26469 , n26468 );
nand ( n26470 , n26459 , n26469 );
buf ( n26471 , n14936 );
and ( n26472 , n14940 , n26471 );
not ( n26473 , n14940 );
and ( n26474 , n26473 , n14937 );
nor ( n26475 , n26472 , n26474 );
not ( n26476 , n26475 );
not ( n26477 , n25545 );
or ( n26478 , n26476 , n26477 );
or ( n26479 , n25683 , n26475 );
nand ( n26480 , n26478 , n26479 );
and ( n26481 , n26480 , n25552 );
not ( n26482 , n26480 );
and ( n26483 , n26482 , n25549 );
nor ( n26484 , n26481 , n26483 );
not ( n26485 , n26484 );
and ( n26486 , n26470 , n26485 );
not ( n26487 , n26470 );
and ( n26488 , n26487 , n26484 );
nor ( n26489 , n26486 , n26488 );
not ( n26490 , n26489 );
not ( n26491 , n26490 );
or ( n26492 , n26446 , n26491 );
nand ( n26493 , n26489 , n26444 );
nand ( n26494 , n26492 , n26493 );
not ( n26495 , n16458 );
not ( n26496 , n7596 );
xor ( n26497 , n22642 , n22646 );
xnor ( n26498 , n26497 , n22656 );
not ( n26499 , n26498 );
or ( n26500 , n26496 , n26499 );
or ( n26501 , n26498 , n7596 );
nand ( n26502 , n26500 , n26501 );
not ( n26503 , n26502 );
or ( n26504 , n26495 , n26503 );
or ( n26505 , n26502 , n25825 );
nand ( n26506 , n26504 , n26505 );
buf ( n26507 , n17849 );
not ( n26508 , n26507 );
not ( n26509 , n24433 );
xor ( n26510 , n24424 , n26509 );
xnor ( n26511 , n26510 , n20427 );
not ( n26512 , n26511 );
or ( n26513 , n26508 , n26512 );
or ( n26514 , n26511 , n26507 );
nand ( n26515 , n26513 , n26514 );
and ( n26516 , n26515 , n26226 );
not ( n26517 , n26515 );
not ( n26518 , n26224 );
not ( n26519 , n26518 );
and ( n26520 , n26517 , n26519 );
nor ( n26521 , n26516 , n26520 );
nand ( n26522 , n26506 , n26521 );
not ( n26523 , n25476 );
not ( n26524 , n20300 );
or ( n26525 , n26523 , n26524 );
or ( n26526 , n20300 , n25476 );
nand ( n26527 , n26525 , n26526 );
and ( n26528 , n26527 , n18462 );
not ( n26529 , n26527 );
buf ( n26530 , n18461 );
and ( n26531 , n26529 , n26530 );
nor ( n26532 , n26528 , n26531 );
not ( n26533 , n26532 );
and ( n26534 , n26522 , n26533 );
not ( n26535 , n26522 );
and ( n26536 , n26535 , n26532 );
nor ( n26537 , n26534 , n26536 );
not ( n26538 , n14691 );
buf ( n26539 , n11260 );
not ( n26540 , n26539 );
not ( n26541 , n14683 );
or ( n26542 , n26540 , n26541 );
or ( n26543 , n14683 , n26539 );
nand ( n26544 , n26542 , n26543 );
not ( n26545 , n26544 );
not ( n26546 , n26545 );
or ( n26547 , n26538 , n26546 );
nand ( n26548 , n14692 , n26544 );
nand ( n26549 , n26547 , n26548 );
not ( n26550 , n26549 );
not ( n26551 , n23598 );
not ( n26552 , n9246 );
not ( n26553 , n17717 );
or ( n26554 , n26552 , n26553 );
not ( n26555 , n23593 );
or ( n26556 , n26555 , n9246 );
nand ( n26557 , n26554 , n26556 );
not ( n26558 , n26557 );
or ( n26559 , n26551 , n26558 );
or ( n26560 , n26557 , n17724 );
nand ( n26561 , n26559 , n26560 );
nand ( n26562 , n26550 , n26561 );
not ( n26563 , n26562 );
buf ( n26564 , n6459 );
buf ( n26565 , n26564 );
not ( n26566 , n26565 );
buf ( n26567 , n6460 );
not ( n26568 , n26567 );
not ( n26569 , n26568 );
or ( n26570 , n26566 , n26569 );
not ( n26571 , n26564 );
buf ( n26572 , n26567 );
nand ( n26573 , n26571 , n26572 );
nand ( n26574 , n26570 , n26573 );
buf ( n26575 , n6461 );
not ( n26576 , n26575 );
and ( n26577 , n26574 , n26576 );
not ( n26578 , n26574 );
buf ( n26579 , n26575 );
and ( n26580 , n26578 , n26579 );
nor ( n26581 , n26577 , n26580 );
buf ( n26582 , n6462 );
nand ( n26583 , n8966 , n26582 );
buf ( n26584 , n6463 );
buf ( n26585 , n26584 );
and ( n26586 , n26583 , n26585 );
not ( n26587 , n26583 );
not ( n26588 , n26584 );
and ( n26589 , n26587 , n26588 );
nor ( n26590 , n26586 , n26589 );
xor ( n26591 , n26581 , n26590 );
xor ( n26592 , n26591 , n20242 );
buf ( n26593 , n26592 );
not ( n26594 , n26593 );
buf ( n26595 , n14348 );
not ( n26596 , n26595 );
not ( n26597 , n26596 );
not ( n26598 , n13087 );
or ( n26599 , n26597 , n26598 );
xor ( n26600 , n13066 , n13085 );
buf ( n26601 , n13075 );
xnor ( n26602 , n26600 , n26601 );
nand ( n26603 , n26602 , n26595 );
nand ( n26604 , n26599 , n26603 );
not ( n26605 , n26604 );
or ( n26606 , n26594 , n26605 );
or ( n26607 , n26604 , n26593 );
nand ( n26608 , n26606 , n26607 );
not ( n26609 , n26608 );
and ( n26610 , n26563 , n26609 );
and ( n26611 , n26562 , n26608 );
nor ( n26612 , n26610 , n26611 );
or ( n26613 , n26537 , n26612 );
nand ( n26614 , n26612 , n26537 );
nand ( n26615 , n26613 , n26614 );
not ( n26616 , n12512 );
not ( n26617 , n10096 );
not ( n26618 , n10108 );
xor ( n26619 , n26617 , n26618 );
xnor ( n26620 , n26619 , n10124 );
not ( n26621 , n26620 );
or ( n26622 , n26616 , n26621 );
or ( n26623 , n26620 , n12512 );
nand ( n26624 , n26622 , n26623 );
not ( n26625 , n26624 );
not ( n26626 , n18498 );
not ( n26627 , n18520 );
or ( n26628 , n26626 , n26627 );
nand ( n26629 , n26628 , n18524 );
not ( n26630 , n26629 );
not ( n26631 , n26630 );
and ( n26632 , n26625 , n26631 );
and ( n26633 , n26624 , n26630 );
nor ( n26634 , n26632 , n26633 );
not ( n26635 , n26634 );
not ( n26636 , n8619 );
not ( n26637 , n12459 );
xor ( n26638 , n12265 , n12284 );
not ( n26639 , n12274 );
xnor ( n26640 , n26638 , n26639 );
not ( n26641 , n26640 );
or ( n26642 , n26637 , n26641 );
or ( n26643 , n12286 , n12459 );
nand ( n26644 , n26642 , n26643 );
not ( n26645 , n26644 );
or ( n26646 , n26636 , n26645 );
or ( n26647 , n26644 , n8620 );
nand ( n26648 , n26646 , n26647 );
not ( n26649 , n26648 );
nand ( n26650 , n26635 , n26649 );
not ( n26651 , n26650 );
not ( n26652 , n12236 );
buf ( n26653 , n20036 );
not ( n26654 , n22245 );
and ( n26655 , n26653 , n26654 );
not ( n26656 , n26653 );
and ( n26657 , n26656 , n22245 );
nor ( n26658 , n26655 , n26657 );
not ( n26659 , n26658 );
and ( n26660 , n26652 , n26659 );
and ( n26661 , n12236 , n26658 );
nor ( n26662 , n26660 , n26661 );
not ( n26663 , n26662 );
not ( n26664 , n26663 );
and ( n26665 , n26651 , n26664 );
and ( n26666 , n26650 , n26663 );
nor ( n26667 , n26665 , n26666 );
and ( n26668 , n26615 , n26667 );
not ( n26669 , n26615 );
not ( n26670 , n26667 );
and ( n26671 , n26669 , n26670 );
nor ( n26672 , n26668 , n26671 );
and ( n26673 , n26494 , n26672 );
not ( n26674 , n26494 );
not ( n26675 , n26672 );
and ( n26676 , n26674 , n26675 );
nor ( n26677 , n26673 , n26676 );
not ( n26678 , n26677 );
not ( n26679 , n26678 );
and ( n26680 , n26402 , n26679 );
not ( n26681 , n26402 );
not ( n26682 , n26494 );
not ( n26683 , n26672 );
or ( n26684 , n26682 , n26683 );
not ( n26685 , n26494 );
nand ( n26686 , n26685 , n26675 );
nand ( n26687 , n26684 , n26686 );
buf ( n26688 , n26687 );
and ( n26689 , n26681 , n26688 );
nor ( n26690 , n26680 , n26689 );
nand ( n26691 , n26139 , n26690 );
or ( n26692 , n25662 , n26691 );
not ( n26693 , n25659 );
not ( n26694 , n26690 );
or ( n26695 , n26693 , n26694 );
buf ( n26696 , n13349 );
nor ( n26697 , n26139 , n26696 );
nand ( n26698 , n26695 , n26697 );
buf ( n26699 , n13353 );
nand ( n26700 , n26699 , n7431 );
nand ( n26701 , n26692 , n26698 , n26700 );
buf ( n26702 , n26701 );
buf ( n26703 , n26702 );
xor ( n26704 , n10920 , n24055 );
xnor ( n26705 , n26704 , n24058 );
not ( n26706 , n26705 );
not ( n26707 , n12569 );
not ( n26708 , n26325 );
not ( n26709 , n26708 );
or ( n26710 , n26707 , n26709 );
buf ( n26711 , n25487 );
not ( n26712 , n26711 );
nand ( n26713 , n26712 , n12566 );
nand ( n26714 , n26710 , n26713 );
and ( n26715 , n26714 , n25494 );
not ( n26716 , n26714 );
and ( n26717 , n26716 , n26332 );
nor ( n26718 , n26715 , n26717 );
not ( n26719 , n26718 );
nand ( n26720 , n26706 , n26719 );
not ( n26721 , n26720 );
not ( n26722 , n10227 );
not ( n26723 , n9053 );
not ( n26724 , n23363 );
or ( n26725 , n26723 , n26724 );
not ( n26726 , n9053 );
nand ( n26727 , n26726 , n10175 );
nand ( n26728 , n26725 , n26727 );
not ( n26729 , n26728 );
or ( n26730 , n26722 , n26729 );
or ( n26731 , n26728 , n10227 );
nand ( n26732 , n26730 , n26731 );
buf ( n26733 , n26732 );
not ( n26734 , n26733 );
and ( n26735 , n26721 , n26734 );
and ( n26736 , n26720 , n26733 );
nor ( n26737 , n26735 , n26736 );
not ( n26738 , n26737 );
not ( n26739 , n17298 );
not ( n26740 , n12441 );
or ( n26741 , n26739 , n26740 );
or ( n26742 , n12441 , n17298 );
nand ( n26743 , n26741 , n26742 );
xor ( n26744 , n12462 , n26743 );
not ( n26745 , n19335 );
not ( n26746 , n21230 );
or ( n26747 , n26745 , n26746 );
nand ( n26748 , n21229 , n19331 );
nand ( n26749 , n26747 , n26748 );
and ( n26750 , n26749 , n21265 );
not ( n26751 , n26749 );
and ( n26752 , n26751 , n21262 );
or ( n26753 , n26750 , n26752 );
and ( n26754 , n26753 , n15291 );
not ( n26755 , n26753 );
and ( n26756 , n26755 , n21217 );
nor ( n26757 , n26754 , n26756 );
nand ( n26758 , n26744 , n26757 );
not ( n26759 , n26758 );
not ( n26760 , n22889 );
buf ( n26761 , n16327 );
not ( n26762 , n26761 );
not ( n26763 , n17908 );
or ( n26764 , n26762 , n26763 );
or ( n26765 , n17908 , n26761 );
nand ( n26766 , n26764 , n26765 );
not ( n26767 , n26766 );
or ( n26768 , n26760 , n26767 );
or ( n26769 , n26766 , n22889 );
nand ( n26770 , n26768 , n26769 );
not ( n26771 , n26770 );
and ( n26772 , n26759 , n26771 );
and ( n26773 , n26758 , n26770 );
nor ( n26774 , n26772 , n26773 );
not ( n26775 , n26774 );
not ( n26776 , n23955 );
not ( n26777 , n20937 );
or ( n26778 , n26776 , n26777 );
not ( n26779 , n23955 );
nand ( n26780 , n26779 , n20462 );
nand ( n26781 , n26778 , n26780 );
not ( n26782 , n25987 );
and ( n26783 , n26781 , n26782 );
not ( n26784 , n26781 );
and ( n26785 , n26784 , n15429 );
nor ( n26786 , n26783 , n26785 );
not ( n26787 , n22629 );
not ( n26788 , n14219 );
or ( n26789 , n26787 , n26788 );
not ( n26790 , n14220 );
or ( n26791 , n26790 , n22629 );
nand ( n26792 , n26789 , n26791 );
and ( n26793 , n26792 , n14268 );
not ( n26794 , n26792 );
and ( n26795 , n26794 , n14272 );
nor ( n26796 , n26793 , n26795 );
not ( n26797 , n26796 );
nand ( n26798 , n26786 , n26797 );
not ( n26799 , n6601 );
not ( n26800 , n8547 );
or ( n26801 , n26799 , n26800 );
or ( n26802 , n8547 , n6601 );
nand ( n26803 , n26801 , n26802 );
and ( n26804 , n26803 , n15849 );
not ( n26805 , n26803 );
and ( n26806 , n26805 , n10443 );
nor ( n26807 , n26804 , n26806 );
buf ( n26808 , n26807 );
and ( n26809 , n26798 , n26808 );
not ( n26810 , n26798 );
not ( n26811 , n26808 );
and ( n26812 , n26810 , n26811 );
nor ( n26813 , n26809 , n26812 );
not ( n26814 , n26813 );
or ( n26815 , n26775 , n26814 );
or ( n26816 , n26813 , n26774 );
nand ( n26817 , n26815 , n26816 );
not ( n26818 , n26733 );
nand ( n26819 , n26818 , n26705 );
not ( n26820 , n26819 );
not ( n26821 , n22415 );
not ( n26822 , n13835 );
not ( n26823 , n20202 );
or ( n26824 , n26822 , n26823 );
or ( n26825 , n20199 , n13835 );
nand ( n26826 , n26824 , n26825 );
not ( n26827 , n26826 );
and ( n26828 , n26821 , n26827 );
not ( n26829 , n22415 );
not ( n26830 , n26829 );
and ( n26831 , n26830 , n26826 );
nor ( n26832 , n26828 , n26831 );
not ( n26833 , n26832 );
not ( n26834 , n26833 );
and ( n26835 , n26820 , n26834 );
and ( n26836 , n26819 , n26833 );
nor ( n26837 , n26835 , n26836 );
and ( n26838 , n26817 , n26837 );
not ( n26839 , n26817 );
not ( n26840 , n26837 );
and ( n26841 , n26839 , n26840 );
nor ( n26842 , n26838 , n26841 );
not ( n26843 , n26842 );
buf ( n26844 , n9793 );
not ( n26845 , n26844 );
not ( n26846 , n20557 );
not ( n26847 , n26846 );
or ( n26848 , n26845 , n26847 );
or ( n26849 , n20553 , n26844 );
nand ( n26850 , n26848 , n26849 );
not ( n26851 , n22700 );
and ( n26852 , n26850 , n26851 );
not ( n26853 , n26850 );
buf ( n26854 , n22700 );
and ( n26855 , n26853 , n26854 );
nor ( n26856 , n26852 , n26855 );
not ( n26857 , n9884 );
not ( n26858 , n11727 );
or ( n26859 , n26857 , n26858 );
nand ( n26860 , n26312 , n9880 );
nand ( n26861 , n26859 , n26860 );
and ( n26862 , n26861 , n21854 );
not ( n26863 , n26861 );
and ( n26864 , n26863 , n21857 );
nor ( n26865 , n26862 , n26864 );
nand ( n26866 , n26856 , n26865 );
and ( n26867 , n8437 , n16716 );
not ( n26868 , n8437 );
and ( n26869 , n26868 , n16763 );
or ( n26870 , n26867 , n26869 );
not ( n26871 , n14624 );
and ( n26872 , n26870 , n26871 );
not ( n26873 , n26870 );
not ( n26874 , n14624 );
not ( n26875 , n26874 );
and ( n26876 , n26873 , n26875 );
nor ( n26877 , n26872 , n26876 );
not ( n26878 , n26877 );
and ( n26879 , n26866 , n26878 );
not ( n26880 , n26866 );
and ( n26881 , n26880 , n26877 );
nor ( n26882 , n26879 , n26881 );
not ( n26883 , n26882 );
not ( n26884 , n25326 );
not ( n26885 , n24086 );
or ( n26886 , n26884 , n26885 );
not ( n26887 , n24791 );
not ( n26888 , n26887 );
nand ( n26889 , n26888 , n25322 );
nand ( n26890 , n26886 , n26889 );
xnor ( n26891 , n26890 , n18112 );
not ( n26892 , n26891 );
buf ( n26893 , n6464 );
buf ( n26894 , n26893 );
xor ( n26895 , n26894 , n19200 );
xnor ( n26896 , n26895 , n23548 );
nand ( n26897 , n26892 , n26896 );
not ( n26898 , n26897 );
buf ( n26899 , n6465 );
buf ( n26900 , n26899 );
not ( n26901 , n26900 );
buf ( n26902 , n6466 );
not ( n26903 , n26902 );
not ( n26904 , n26903 );
or ( n26905 , n26901 , n26904 );
not ( n26906 , n26899 );
buf ( n26907 , n26902 );
nand ( n26908 , n26906 , n26907 );
nand ( n26909 , n26905 , n26908 );
buf ( n26910 , n6467 );
not ( n26911 , n26910 );
and ( n26912 , n26909 , n26911 );
not ( n26913 , n26909 );
buf ( n26914 , n26910 );
and ( n26915 , n26913 , n26914 );
nor ( n26916 , n26912 , n26915 );
buf ( n26917 , n6468 );
nand ( n26918 , n7912 , n26917 );
buf ( n26919 , n6469 );
buf ( n26920 , n26919 );
and ( n26921 , n26918 , n26920 );
not ( n26922 , n26918 );
not ( n26923 , n26919 );
and ( n26924 , n26922 , n26923 );
nor ( n26925 , n26921 , n26924 );
xor ( n26926 , n26916 , n26925 );
buf ( n26927 , n6470 );
nand ( n26928 , n8455 , n26927 );
buf ( n26929 , n6471 );
buf ( n26930 , n26929 );
and ( n26931 , n26928 , n26930 );
not ( n26932 , n26928 );
not ( n26933 , n26929 );
and ( n26934 , n26932 , n26933 );
nor ( n26935 , n26931 , n26934 );
xor ( n26936 , n26926 , n26935 );
not ( n26937 , n26936 );
xor ( n26938 , n17766 , n26937 );
xnor ( n26939 , n26938 , n26630 );
not ( n26940 , n26939 );
and ( n26941 , n26898 , n26940 );
not ( n26942 , n26891 );
nand ( n26943 , n26942 , n26896 );
and ( n26944 , n26943 , n26939 );
nor ( n26945 , n26941 , n26944 );
not ( n26946 , n26945 );
or ( n26947 , n26883 , n26946 );
or ( n26948 , n26945 , n26882 );
nand ( n26949 , n26947 , n26948 );
not ( n26950 , n26949 );
or ( n26951 , n26843 , n26950 );
not ( n26952 , n26949 );
not ( n26953 , n26842 );
nand ( n26954 , n26952 , n26953 );
nand ( n26955 , n26951 , n26954 );
not ( n26956 , n26955 );
or ( n26957 , n26738 , n26956 );
not ( n26958 , n26737 );
not ( n26959 , n26952 );
not ( n26960 , n26953 );
and ( n26961 , n26959 , n26960 );
and ( n26962 , n26952 , n26953 );
nor ( n26963 , n26961 , n26962 );
nand ( n26964 , n26958 , n26963 );
nand ( n26965 , n26957 , n26964 );
buf ( n26966 , n26393 );
and ( n26967 , n26965 , n26966 );
not ( n26968 , n26965 );
buf ( n26969 , n26400 );
and ( n26970 , n26968 , n26969 );
nor ( n26971 , n26967 , n26970 );
not ( n26972 , n26971 );
not ( n26973 , n23398 );
not ( n26974 , n26973 );
not ( n26975 , n10011 );
not ( n26976 , n10498 );
not ( n26977 , n15748 );
or ( n26978 , n26976 , n26977 );
or ( n26979 , n15748 , n10498 );
nand ( n26980 , n26978 , n26979 );
not ( n26981 , n26980 );
and ( n26982 , n26975 , n26981 );
and ( n26983 , n10011 , n26980 );
nor ( n26984 , n26982 , n26983 );
not ( n26985 , n26984 );
not ( n26986 , n26985 );
not ( n26987 , n26116 );
nand ( n26988 , n26987 , n26110 );
not ( n26989 , n26988 );
or ( n26990 , n26986 , n26989 );
or ( n26991 , n26988 , n26985 );
nand ( n26992 , n26990 , n26991 );
not ( n26993 , n26992 );
not ( n26994 , n17508 );
not ( n26995 , n20337 );
or ( n26996 , n26994 , n26995 );
not ( n26997 , n17508 );
nand ( n26998 , n26997 , n23209 );
nand ( n26999 , n26996 , n26998 );
not ( n27000 , n18897 );
and ( n27001 , n26999 , n27000 );
not ( n27002 , n26999 );
and ( n27003 , n27002 , n18897 );
nor ( n27004 , n27001 , n27003 );
nand ( n27005 , n27004 , n26045 );
not ( n27006 , n27005 );
not ( n27007 , n7756 );
and ( n27008 , n11025 , n9730 );
not ( n27009 , n11025 );
and ( n27010 , n27009 , n18667 );
nor ( n27011 , n27008 , n27010 );
not ( n27012 , n27011 );
not ( n27013 , n27012 );
or ( n27014 , n27007 , n27013 );
nand ( n27015 , n27011 , n25257 );
nand ( n27016 , n27014 , n27015 );
not ( n27017 , n27016 );
or ( n27018 , n27006 , n27017 );
or ( n27019 , n27016 , n27005 );
nand ( n27020 , n27018 , n27019 );
not ( n27021 , n27020 );
not ( n27022 , n27021 );
nand ( n27023 , n26984 , n26116 );
not ( n27024 , n27023 );
not ( n27025 , n19652 );
not ( n27026 , n17139 );
or ( n27027 , n27025 , n27026 );
nand ( n27028 , n9898 , n19648 );
nand ( n27029 , n27027 , n27028 );
not ( n27030 , n27029 );
not ( n27031 , n9942 );
and ( n27032 , n27030 , n27031 );
and ( n27033 , n27029 , n9942 );
nor ( n27034 , n27032 , n27033 );
not ( n27035 , n27034 );
not ( n27036 , n27035 );
and ( n27037 , n27024 , n27036 );
and ( n27038 , n27023 , n27035 );
nor ( n27039 , n27037 , n27038 );
not ( n27040 , n27039 );
not ( n27041 , n27040 );
or ( n27042 , n27022 , n27041 );
nand ( n27043 , n27039 , n27020 );
nand ( n27044 , n27042 , n27043 );
not ( n27045 , n15481 );
buf ( n27046 , n6472 );
not ( n27047 , n26894 );
not ( n27048 , n23545 );
not ( n27049 , n27048 );
or ( n27050 , n27047 , n27049 );
not ( n27051 , n26893 );
nand ( n27052 , n27051 , n23546 );
nand ( n27053 , n27050 , n27052 );
xor ( n27054 , n27046 , n27053 );
not ( n27055 , n19132 );
buf ( n27056 , n6473 );
nand ( n27057 , n6557 , n27056 );
buf ( n27058 , n6474 );
buf ( n27059 , n27058 );
and ( n27060 , n27057 , n27059 );
not ( n27061 , n27057 );
not ( n27062 , n27058 );
and ( n27063 , n27061 , n27062 );
nor ( n27064 , n27060 , n27063 );
not ( n27065 , n27064 );
not ( n27066 , n27065 );
or ( n27067 , n27055 , n27066 );
nand ( n27068 , n27064 , n19116 );
nand ( n27069 , n27067 , n27068 );
xnor ( n27070 , n27054 , n27069 );
buf ( n27071 , n27070 );
not ( n27072 , n27071 );
or ( n27073 , n27045 , n27072 );
or ( n27074 , n27071 , n15481 );
nand ( n27075 , n27073 , n27074 );
and ( n27076 , n27075 , n25767 );
not ( n27077 , n27075 );
and ( n27078 , n27077 , n9136 );
nor ( n27079 , n27076 , n27078 );
nand ( n27080 , n27079 , n26081 );
not ( n27081 , n27080 );
xor ( n27082 , n16519 , n16538 );
not ( n27083 , n16528 );
xor ( n27084 , n27082 , n27083 );
not ( n27085 , n27084 );
not ( n27086 , n27085 );
not ( n27087 , n15772 );
and ( n27088 , n27086 , n27087 );
and ( n27089 , n16541 , n15772 );
nor ( n27090 , n27088 , n27089 );
and ( n27091 , n27090 , n16058 );
not ( n27092 , n27090 );
not ( n27093 , n16057 );
not ( n27094 , n27093 );
buf ( n27095 , n27094 );
and ( n27096 , n27092 , n27095 );
nor ( n27097 , n27091 , n27096 );
buf ( n27098 , n27097 );
not ( n27099 , n27098 );
and ( n27100 , n27081 , n27099 );
and ( n27101 , n27080 , n27098 );
nor ( n27102 , n27100 , n27101 );
not ( n27103 , n27102 );
and ( n27104 , n27044 , n27103 );
not ( n27105 , n27044 );
and ( n27106 , n27105 , n27102 );
nor ( n27107 , n27104 , n27106 );
not ( n27108 , n14230 );
buf ( n27109 , n17860 );
not ( n27110 , n27109 );
or ( n27111 , n27108 , n27110 );
or ( n27112 , n17862 , n14230 );
nand ( n27113 , n27111 , n27112 );
not ( n27114 , n27113 );
not ( n27115 , n22465 );
not ( n27116 , n27115 );
and ( n27117 , n27114 , n27116 );
not ( n27118 , n22464 );
buf ( n27119 , n27118 );
and ( n27120 , n27113 , n27119 );
nor ( n27121 , n27117 , n27120 );
nand ( n27122 , n26003 , n27121 );
not ( n27123 , n27122 );
not ( n27124 , n14018 );
not ( n27125 , n10958 );
or ( n27126 , n27124 , n27125 );
or ( n27127 , n10958 , n14018 );
nand ( n27128 , n27126 , n27127 );
and ( n27129 , n27128 , n13007 );
not ( n27130 , n27128 );
and ( n27131 , n27130 , n12994 );
nor ( n27132 , n27129 , n27131 );
not ( n27133 , n27132 );
and ( n27134 , n27123 , n27133 );
and ( n27135 , n27122 , n27132 );
nor ( n27136 , n27134 , n27135 );
not ( n27137 , n27136 );
not ( n27138 , n27137 );
not ( n27139 , n21598 );
not ( n27140 , n19833 );
or ( n27141 , n27139 , n27140 );
or ( n27142 , n19833 , n21598 );
nand ( n27143 , n27141 , n27142 );
not ( n27144 , n8786 );
and ( n27145 , n27143 , n27144 );
not ( n27146 , n27143 );
and ( n27147 , n27146 , n8786 );
nor ( n27148 , n27145 , n27147 );
not ( n27149 , n27148 );
not ( n27150 , n27149 );
not ( n27151 , n9056 );
not ( n27152 , n23363 );
or ( n27153 , n27151 , n27152 );
buf ( n27154 , n10175 );
nand ( n27155 , n27154 , n9051 );
nand ( n27156 , n27153 , n27155 );
and ( n27157 , n27156 , n10228 );
not ( n27158 , n27156 );
and ( n27159 , n27158 , n25838 );
nor ( n27160 , n27157 , n27159 );
nand ( n27161 , n25969 , n27160 );
not ( n27162 , n27161 );
or ( n27163 , n27150 , n27162 );
or ( n27164 , n27161 , n27149 );
nand ( n27165 , n27163 , n27164 );
not ( n27166 , n27165 );
not ( n27167 , n27166 );
or ( n27168 , n27138 , n27167 );
nand ( n27169 , n27165 , n27136 );
nand ( n27170 , n27168 , n27169 );
not ( n27171 , n27170 );
and ( n27172 , n27107 , n27171 );
not ( n27173 , n27107 );
and ( n27174 , n27173 , n27170 );
nor ( n27175 , n27172 , n27174 );
not ( n27176 , n27175 );
or ( n27177 , n26993 , n27176 );
not ( n27178 , n27175 );
not ( n27179 , n26992 );
nand ( n27180 , n27178 , n27179 );
nand ( n27181 , n27177 , n27180 );
not ( n27182 , n27181 );
and ( n27183 , n26974 , n27182 );
not ( n27184 , n23398 );
and ( n27185 , n27184 , n27181 );
nor ( n27186 , n27183 , n27185 );
nand ( n27187 , n26972 , n27186 );
not ( n27188 , n24155 );
not ( n27189 , n16352 );
not ( n27190 , n17904 );
or ( n27191 , n27189 , n27190 );
or ( n27192 , n17904 , n16352 );
nand ( n27193 , n27191 , n27192 );
and ( n27194 , n27193 , n17908 );
not ( n27195 , n27193 );
and ( n27196 , n27195 , n13399 );
nor ( n27197 , n27194 , n27196 );
nand ( n27198 , n24168 , n27197 );
not ( n27199 , n27198 );
or ( n27200 , n27188 , n27199 );
or ( n27201 , n27198 , n24155 );
nand ( n27202 , n27200 , n27201 );
not ( n27203 , n27202 );
not ( n27204 , n24245 );
or ( n27205 , n27203 , n27204 );
not ( n27206 , n27202 );
nand ( n27207 , n27206 , n24254 );
nand ( n27208 , n27205 , n27207 );
and ( n27209 , n27208 , n24259 );
not ( n27210 , n27208 );
and ( n27211 , n27210 , n23933 );
nor ( n27212 , n27209 , n27211 );
not ( n27213 , n27212 );
buf ( n27214 , n13345 );
nor ( n27215 , n27213 , n27214 );
not ( n27216 , n27215 );
or ( n27217 , n27187 , n27216 );
nand ( n27218 , n27212 , n27186 );
not ( n27219 , n20976 );
nand ( n27220 , n27218 , n26971 , n27219 );
nand ( n27221 , n17813 , n20455 );
nand ( n27222 , n27217 , n27220 , n27221 );
buf ( n27223 , n27222 );
buf ( n27224 , n27223 );
not ( n27225 , n8866 );
xor ( n27226 , n27225 , n8885 );
xnor ( n27227 , n27226 , n8875 );
and ( n27228 , n17588 , n27227 );
not ( n27229 , n17588 );
and ( n27230 , n27229 , n8888 );
nor ( n27231 , n27228 , n27230 );
buf ( n27232 , n8913 );
not ( n27233 , n27232 );
and ( n27234 , n27231 , n27233 );
not ( n27235 , n27231 );
and ( n27236 , n27235 , n27232 );
nor ( n27237 , n27234 , n27236 );
not ( n27238 , n27237 );
not ( n27239 , n10110 );
not ( n27240 , n24961 );
or ( n27241 , n27239 , n27240 );
not ( n27242 , n10110 );
nand ( n27243 , n27242 , n25791 );
nand ( n27244 , n27241 , n27243 );
and ( n27245 , n27244 , n12713 );
not ( n27246 , n27244 );
and ( n27247 , n27246 , n22817 );
nor ( n27248 , n27245 , n27247 );
nand ( n27249 , n27238 , n27248 );
not ( n27250 , n27249 );
not ( n27251 , n14244 );
not ( n27252 , n17860 );
not ( n27253 , n27252 );
not ( n27254 , n27253 );
or ( n27255 , n27251 , n27254 );
not ( n27256 , n14244 );
nand ( n27257 , n27256 , n17861 );
nand ( n27258 , n27255 , n27257 );
and ( n27259 , n27258 , n27119 );
not ( n27260 , n27258 );
not ( n27261 , n27115 );
and ( n27262 , n27260 , n27261 );
nor ( n27263 , n27259 , n27262 );
not ( n27264 , n27263 );
not ( n27265 , n27264 );
and ( n27266 , n27250 , n27265 );
and ( n27267 , n27249 , n27264 );
nor ( n27268 , n27266 , n27267 );
not ( n27269 , n27268 );
nand ( n27270 , n27237 , n27263 );
not ( n27271 , n27270 );
not ( n27272 , n21506 );
not ( n27273 , n7922 );
not ( n27274 , n27273 );
or ( n27275 , n27272 , n27274 );
or ( n27276 , n27273 , n21506 );
nand ( n27277 , n27275 , n27276 );
and ( n27278 , n27277 , n7879 );
not ( n27279 , n27277 );
and ( n27280 , n27279 , n21189 );
nor ( n27281 , n27278 , n27280 );
not ( n27282 , n27281 );
not ( n27283 , n27282 );
and ( n27284 , n27271 , n27283 );
and ( n27285 , n27270 , n27282 );
nor ( n27286 , n27284 , n27285 );
not ( n27287 , n27286 );
buf ( n27288 , n8711 );
not ( n27289 , n27288 );
not ( n27290 , n10850 );
or ( n27291 , n27289 , n27290 );
or ( n27292 , n10850 , n27288 );
nand ( n27293 , n27291 , n27292 );
and ( n27294 , n27293 , n10826 );
not ( n27295 , n27293 );
and ( n27296 , n27295 , n25964 );
nor ( n27297 , n27294 , n27296 );
buf ( n27298 , n13030 );
not ( n27299 , n27298 );
not ( n27300 , n21991 );
or ( n27301 , n27299 , n27300 );
or ( n27302 , n21991 , n27298 );
nand ( n27303 , n27301 , n27302 );
and ( n27304 , n27303 , n15046 );
not ( n27305 , n27303 );
and ( n27306 , n27305 , n15053 );
nor ( n27307 , n27304 , n27306 );
nand ( n27308 , n27297 , n27307 );
not ( n27309 , n17767 );
not ( n27310 , n16503 );
and ( n27311 , n27309 , n27310 );
and ( n27312 , n17767 , n16503 );
nor ( n27313 , n27311 , n27312 );
xor ( n27314 , n14175 , n27313 );
and ( n27315 , n27308 , n27314 );
not ( n27316 , n27308 );
not ( n27317 , n27314 );
and ( n27318 , n27316 , n27317 );
nor ( n27319 , n27315 , n27318 );
not ( n27320 , n27319 );
or ( n27321 , n27287 , n27320 );
or ( n27322 , n27319 , n27286 );
nand ( n27323 , n27321 , n27322 );
buf ( n27324 , n26222 );
not ( n27325 , n27324 );
not ( n27326 , n27325 );
not ( n27327 , n18082 );
or ( n27328 , n27326 , n27327 );
nand ( n27329 , n22733 , n27324 );
nand ( n27330 , n27328 , n27329 );
not ( n27331 , n27330 );
not ( n27332 , n8762 );
or ( n27333 , n27331 , n27332 );
or ( n27334 , n22741 , n27330 );
nand ( n27335 , n27333 , n27334 );
not ( n27336 , n15073 );
not ( n27337 , n15701 );
or ( n27338 , n27336 , n27337 );
or ( n27339 , n14509 , n15073 );
nand ( n27340 , n27338 , n27339 );
not ( n27341 , n27340 );
not ( n27342 , n16898 );
and ( n27343 , n27341 , n27342 );
and ( n27344 , n27340 , n22757 );
nor ( n27345 , n27343 , n27344 );
nand ( n27346 , n27335 , n27345 );
not ( n27347 , n10036 );
not ( n27348 , n27347 );
xor ( n27349 , n25275 , n27348 );
xnor ( n27350 , n27349 , n18112 );
and ( n27351 , n27346 , n27350 );
not ( n27352 , n27346 );
not ( n27353 , n27350 );
and ( n27354 , n27352 , n27353 );
nor ( n27355 , n27351 , n27354 );
xor ( n27356 , n27323 , n27355 );
not ( n27357 , n27356 );
not ( n27358 , n10823 );
not ( n27359 , n18705 );
or ( n27360 , n27358 , n27359 );
not ( n27361 , n10823 );
nand ( n27362 , n27361 , n22563 );
nand ( n27363 , n27360 , n27362 );
buf ( n27364 , n12342 );
and ( n27365 , n27363 , n27364 );
not ( n27366 , n27363 );
and ( n27367 , n27366 , n18714 );
nor ( n27368 , n27365 , n27367 );
not ( n27369 , n27368 );
xor ( n27370 , n23959 , n15428 );
xnor ( n27371 , n27370 , n20464 );
nand ( n27372 , n27369 , n27371 );
not ( n27373 , n27372 );
not ( n27374 , n8766 );
not ( n27375 , n11272 );
or ( n27376 , n27374 , n27375 );
or ( n27377 , n11272 , n8766 );
nand ( n27378 , n27376 , n27377 );
not ( n27379 , n17419 );
not ( n27380 , n27379 );
and ( n27381 , n27378 , n27380 );
not ( n27382 , n27378 );
buf ( n27383 , n17190 );
and ( n27384 , n27382 , n27383 );
nor ( n27385 , n27381 , n27384 );
not ( n27386 , n27385 );
and ( n27387 , n27373 , n27386 );
not ( n27388 , n27368 );
nand ( n27389 , n27371 , n27388 );
and ( n27390 , n27389 , n27385 );
nor ( n27391 , n27387 , n27390 );
not ( n27392 , n27391 );
and ( n27393 , n9595 , n9592 );
not ( n27394 , n9595 );
buf ( n27395 , n9591 );
and ( n27396 , n27394 , n27395 );
nor ( n27397 , n27393 , n27396 );
xor ( n27398 , n27397 , n23408 );
xnor ( n27399 , n27398 , n10679 );
not ( n27400 , n8065 );
not ( n27401 , n6729 );
or ( n27402 , n27400 , n27401 );
or ( n27403 , n6731 , n8065 );
nand ( n27404 , n27402 , n27403 );
not ( n27405 , n27404 );
not ( n27406 , n11108 );
and ( n27407 , n27405 , n27406 );
not ( n27408 , n6685 );
and ( n27409 , n27404 , n27408 );
nor ( n27410 , n27407 , n27409 );
nand ( n27411 , n27399 , n27410 );
not ( n27412 , n14362 );
buf ( n27413 , n26602 );
not ( n27414 , n27413 );
or ( n27415 , n27412 , n27414 );
or ( n27416 , n27413 , n14362 );
nand ( n27417 , n27415 , n27416 );
not ( n27418 , n26592 );
not ( n27419 , n27418 );
and ( n27420 , n27417 , n27419 );
not ( n27421 , n27417 );
xor ( n27422 , n26581 , n20242 );
buf ( n27423 , n26590 );
xnor ( n27424 , n27422 , n27423 );
not ( n27425 , n27424 );
not ( n27426 , n27425 );
and ( n27427 , n27421 , n27426 );
nor ( n27428 , n27420 , n27427 );
and ( n27429 , n27411 , n27428 );
not ( n27430 , n27411 );
not ( n27431 , n27428 );
and ( n27432 , n27430 , n27431 );
nor ( n27433 , n27429 , n27432 );
not ( n27434 , n27433 );
or ( n27435 , n27392 , n27434 );
or ( n27436 , n27433 , n27391 );
nand ( n27437 , n27435 , n27436 );
not ( n27438 , n27437 );
not ( n27439 , n27438 );
or ( n27440 , n27357 , n27439 );
not ( n27441 , n27356 );
nand ( n27442 , n27441 , n27437 );
nand ( n27443 , n27440 , n27442 );
not ( n27444 , n27443 );
or ( n27445 , n27269 , n27444 );
or ( n27446 , n27443 , n27268 );
nand ( n27447 , n27445 , n27446 );
not ( n27448 , n27447 );
buf ( n27449 , n21523 );
not ( n27450 , n27449 );
not ( n27451 , n7926 );
or ( n27452 , n27450 , n27451 );
or ( n27453 , n7926 , n27449 );
nand ( n27454 , n27452 , n27453 );
and ( n27455 , n27454 , n21189 );
not ( n27456 , n27454 );
and ( n27457 , n27456 , n7879 );
nor ( n27458 , n27455 , n27457 );
not ( n27459 , n18343 );
not ( n27460 , n23174 );
or ( n27461 , n27459 , n27460 );
or ( n27462 , n23174 , n18343 );
nand ( n27463 , n27461 , n27462 );
buf ( n27464 , n20038 );
not ( n27465 , n27464 );
and ( n27466 , n27463 , n27465 );
not ( n27467 , n27463 );
not ( n27468 , n20038 );
not ( n27469 , n27468 );
and ( n27470 , n27467 , n27469 );
nor ( n27471 , n27466 , n27470 );
nor ( n27472 , n27458 , n27471 );
xor ( n27473 , n18703 , n17707 );
xnor ( n27474 , n27473 , n23384 );
not ( n27475 , n27474 );
and ( n27476 , n27472 , n27475 );
not ( n27477 , n27472 );
and ( n27478 , n27477 , n27474 );
nor ( n27479 , n27476 , n27478 );
not ( n27480 , n27479 );
not ( n27481 , n27480 );
not ( n27482 , n10550 );
not ( n27483 , n10010 );
or ( n27484 , n27482 , n27483 );
or ( n27485 , n10010 , n10550 );
nand ( n27486 , n27484 , n27485 );
and ( n27487 , n27486 , n13457 );
not ( n27488 , n27486 );
and ( n27489 , n27488 , n9990 );
nor ( n27490 , n27487 , n27489 );
not ( n27491 , n27490 );
not ( n27492 , n15786 );
not ( n27493 , n16541 );
or ( n27494 , n27492 , n27493 );
not ( n27495 , n15786 );
nand ( n27496 , n27495 , n16540 );
nand ( n27497 , n27494 , n27496 );
and ( n27498 , n27497 , n16058 );
not ( n27499 , n27497 );
and ( n27500 , n27499 , n27095 );
nor ( n27501 , n27498 , n27500 );
nand ( n27502 , n27491 , n27501 );
not ( n27503 , n27502 );
not ( n27504 , n16178 );
buf ( n27505 , n19470 );
xor ( n27506 , n27504 , n27505 );
xnor ( n27507 , n27506 , n10351 );
not ( n27508 , n27507 );
or ( n27509 , n27503 , n27508 );
nand ( n27510 , n27491 , n27501 );
or ( n27511 , n27507 , n27510 );
nand ( n27512 , n27509 , n27511 );
not ( n27513 , n27512 );
not ( n27514 , n27513 );
or ( n27515 , n27481 , n27514 );
nand ( n27516 , n27512 , n27479 );
nand ( n27517 , n27515 , n27516 );
not ( n27518 , n27517 );
buf ( n27519 , n15097 );
not ( n27520 , n27519 );
not ( n27521 , n14507 );
or ( n27522 , n27520 , n27521 );
or ( n27523 , n14507 , n27519 );
nand ( n27524 , n27522 , n27523 );
and ( n27525 , n27524 , n22756 );
not ( n27526 , n27524 );
and ( n27527 , n27526 , n15745 );
nor ( n27528 , n27525 , n27527 );
not ( n27529 , n27528 );
buf ( n27530 , n13590 );
not ( n27531 , n27530 );
not ( n27532 , n19243 );
or ( n27533 , n27531 , n27532 );
or ( n27534 , n19243 , n27530 );
nand ( n27535 , n27533 , n27534 );
and ( n27536 , n27535 , n11272 );
not ( n27537 , n27535 );
and ( n27538 , n27537 , n11275 );
nor ( n27539 , n27536 , n27538 );
not ( n27540 , n9598 );
not ( n27541 , n9911 );
not ( n27542 , n21854 );
or ( n27543 , n27541 , n27542 );
or ( n27544 , n21854 , n9911 );
nand ( n27545 , n27543 , n27544 );
not ( n27546 , n27545 );
or ( n27547 , n27540 , n27546 );
or ( n27548 , n9598 , n27545 );
nand ( n27549 , n27547 , n27548 );
nand ( n27550 , n27539 , n27549 );
not ( n27551 , n27550 );
or ( n27552 , n27529 , n27551 );
or ( n27553 , n27550 , n27528 );
nand ( n27554 , n27552 , n27553 );
not ( n27555 , n27554 );
not ( n27556 , n11105 );
not ( n27557 , n8089 );
not ( n27558 , n6730 );
or ( n27559 , n27557 , n27558 );
not ( n27560 , n8090 );
or ( n27561 , n6734 , n27560 );
nand ( n27562 , n27559 , n27561 );
not ( n27563 , n27562 );
and ( n27564 , n27556 , n27563 );
and ( n27565 , n6741 , n27562 );
nor ( n27566 , n27564 , n27565 );
not ( n27567 , n25311 );
not ( n27568 , n27567 );
not ( n27569 , n27568 );
not ( n27570 , n23305 );
xor ( n27571 , n25335 , n24788 );
xnor ( n27572 , n27571 , n25345 );
not ( n27573 , n27572 );
or ( n27574 , n27570 , n27573 );
or ( n27575 , n27572 , n23305 );
nand ( n27576 , n27574 , n27575 );
not ( n27577 , n27576 );
or ( n27578 , n27569 , n27577 );
or ( n27579 , n27576 , n25312 );
nand ( n27580 , n27578 , n27579 );
nand ( n27581 , n27566 , n27580 );
not ( n27582 , n27581 );
not ( n27583 , n22370 );
not ( n27584 , n15974 );
or ( n27585 , n27583 , n27584 );
not ( n27586 , n22370 );
nand ( n27587 , n27586 , n20845 );
nand ( n27588 , n27585 , n27587 );
not ( n27589 , n27588 );
not ( n27590 , n22557 );
and ( n27591 , n27589 , n27590 );
not ( n27592 , n21444 );
and ( n27593 , n27588 , n27592 );
nor ( n27594 , n27591 , n27593 );
not ( n27595 , n27594 );
not ( n27596 , n27595 );
and ( n27597 , n27582 , n27596 );
and ( n27598 , n27581 , n27595 );
nor ( n27599 , n27597 , n27598 );
not ( n27600 , n27599 );
or ( n27601 , n27555 , n27600 );
or ( n27602 , n27599 , n27554 );
nand ( n27603 , n27601 , n27602 );
not ( n27604 , n7268 );
not ( n27605 , n12466 );
or ( n27606 , n27604 , n27605 );
not ( n27607 , n7268 );
nand ( n27608 , n27607 , n12462 );
nand ( n27609 , n27606 , n27608 );
not ( n27610 , n21949 );
buf ( n27611 , n27610 );
xor ( n27612 , n27609 , n27611 );
not ( n27613 , n11509 );
not ( n27614 , n11554 );
not ( n27615 , n7410 );
not ( n27616 , n27615 );
or ( n27617 , n27614 , n27616 );
or ( n27618 , n27615 , n11554 );
nand ( n27619 , n27617 , n27618 );
not ( n27620 , n27619 );
or ( n27621 , n27613 , n27620 );
or ( n27622 , n27619 , n11509 );
nand ( n27623 , n27621 , n27622 );
nand ( n27624 , n27612 , n27623 );
not ( n27625 , n27624 );
not ( n27626 , n7823 );
not ( n27627 , n7826 );
or ( n27628 , n27626 , n27627 );
or ( n27629 , n7826 , n7823 );
nand ( n27630 , n27628 , n27629 );
not ( n27631 , n27630 );
not ( n27632 , n17589 );
or ( n27633 , n27631 , n27632 );
not ( n27634 , n27630 );
nand ( n27635 , n27634 , n17602 );
nand ( n27636 , n27633 , n27635 );
and ( n27637 , n27636 , n10695 );
not ( n27638 , n27636 );
and ( n27639 , n27638 , n9788 );
nor ( n27640 , n27637 , n27639 );
buf ( n27641 , n27640 );
not ( n27642 , n27641 );
and ( n27643 , n27625 , n27642 );
and ( n27644 , n27624 , n27641 );
nor ( n27645 , n27643 , n27644 );
and ( n27646 , n27603 , n27645 );
not ( n27647 , n27603 );
not ( n27648 , n27645 );
and ( n27649 , n27647 , n27648 );
nor ( n27650 , n27646 , n27649 );
not ( n27651 , n27650 );
and ( n27652 , n27518 , n27651 );
and ( n27653 , n27517 , n27650 );
nor ( n27654 , n27652 , n27653 );
buf ( n27655 , n27654 );
not ( n27656 , n27655 );
and ( n27657 , n27448 , n27656 );
and ( n27658 , n27447 , n27655 );
nor ( n27659 , n27657 , n27658 );
buf ( n27660 , n21737 );
nand ( n27661 , n27659 , n27660 );
not ( n27662 , n11235 );
not ( n27663 , n20571 );
or ( n27664 , n27662 , n27663 );
or ( n27665 , n20576 , n11235 );
nand ( n27666 , n27664 , n27665 );
and ( n27667 , n27666 , n14691 );
not ( n27668 , n27666 );
and ( n27669 , n27668 , n14692 );
nor ( n27670 , n27667 , n27669 );
nand ( n27671 , n23366 , n27670 );
and ( n27672 , n27671 , n23378 );
not ( n27673 , n27671 );
and ( n27674 , n27673 , n23379 );
or ( n27675 , n27672 , n27674 );
not ( n27676 , n27675 );
not ( n27677 , n23399 );
or ( n27678 , n27676 , n27677 );
not ( n27679 , n27675 );
nand ( n27680 , n27679 , n23398 );
nand ( n27681 , n27678 , n27680 );
and ( n27682 , n27681 , n23671 );
not ( n27683 , n27681 );
and ( n27684 , n27683 , n23661 );
nor ( n27685 , n27682 , n27684 );
xor ( n27686 , n20171 , n21622 );
not ( n27687 , n15159 );
not ( n27688 , n15183 );
or ( n27689 , n27687 , n27688 );
nand ( n27690 , n27689 , n15186 );
xnor ( n27691 , n27686 , n27690 );
not ( n27692 , n27691 );
and ( n27693 , n26639 , n20782 );
not ( n27694 , n26639 );
and ( n27695 , n27694 , n20776 );
nor ( n27696 , n27693 , n27695 );
not ( n27697 , n27696 );
and ( n27698 , n25815 , n27697 );
not ( n27699 , n25815 );
and ( n27700 , n27699 , n27696 );
nor ( n27701 , n27698 , n27700 );
not ( n27702 , n8907 );
not ( n27703 , n16193 );
or ( n27704 , n27702 , n27703 );
not ( n27705 , n8906 );
nand ( n27706 , n16167 , n27705 );
nand ( n27707 , n27704 , n27706 );
not ( n27708 , n27707 );
not ( n27709 , n16190 );
or ( n27710 , n27708 , n27709 );
or ( n27711 , n16190 , n27707 );
nand ( n27712 , n27710 , n27711 );
and ( n27713 , n27712 , n13676 );
not ( n27714 , n27712 );
and ( n27715 , n27714 , n13690 );
nor ( n27716 , n27713 , n27715 );
not ( n27717 , n27716 );
nor ( n27718 , n27701 , n27717 );
not ( n27719 , n27718 );
and ( n27720 , n27692 , n27719 );
and ( n27721 , n27691 , n27718 );
nor ( n27722 , n27720 , n27721 );
not ( n27723 , n27722 );
not ( n27724 , n17189 );
not ( n27725 , n14651 );
or ( n27726 , n27724 , n27725 );
or ( n27727 , n14651 , n17189 );
nand ( n27728 , n27726 , n27727 );
and ( n27729 , n27728 , n24925 );
not ( n27730 , n27728 );
not ( n27731 , n24902 );
not ( n27732 , n24924 );
not ( n27733 , n27732 );
or ( n27734 , n27731 , n27733 );
nand ( n27735 , n24924 , n24903 );
nand ( n27736 , n27734 , n27735 );
and ( n27737 , n27730 , n27736 );
nor ( n27738 , n27729 , n27737 );
not ( n27739 , n13225 );
not ( n27740 , n14792 );
or ( n27741 , n27739 , n27740 );
or ( n27742 , n14792 , n13225 );
nand ( n27743 , n27741 , n27742 );
and ( n27744 , n27743 , n14845 );
not ( n27745 , n27743 );
and ( n27746 , n27745 , n14838 );
nor ( n27747 , n27744 , n27746 );
not ( n27748 , n27747 );
nand ( n27749 , n27738 , n27748 );
xor ( n27750 , n27046 , n19200 );
xnor ( n27751 , n27750 , n20089 );
and ( n27752 , n27749 , n27751 );
not ( n27753 , n27749 );
not ( n27754 , n27751 );
and ( n27755 , n27753 , n27754 );
nor ( n27756 , n27752 , n27755 );
not ( n27757 , n27756 );
or ( n27758 , n27723 , n27757 );
or ( n27759 , n27722 , n27756 );
nand ( n27760 , n27758 , n27759 );
not ( n27761 , n13579 );
not ( n27762 , n27761 );
not ( n27763 , n19243 );
or ( n27764 , n27762 , n27763 );
nand ( n27765 , n22765 , n13579 );
nand ( n27766 , n27764 , n27765 );
and ( n27767 , n27766 , n11275 );
not ( n27768 , n27766 );
and ( n27769 , n27768 , n11272 );
nor ( n27770 , n27767 , n27769 );
not ( n27771 , n27770 );
buf ( n27772 , n21440 );
not ( n27773 , n27772 );
not ( n27774 , n27773 );
not ( n27775 , n8046 );
or ( n27776 , n27774 , n27775 );
nand ( n27777 , n8047 , n27772 );
nand ( n27778 , n27776 , n27777 );
not ( n27779 , n27778 );
not ( n27780 , n7993 );
and ( n27781 , n27779 , n27780 );
and ( n27782 , n23384 , n27778 );
nor ( n27783 , n27781 , n27782 );
not ( n27784 , n27783 );
nand ( n27785 , n27771 , n27784 );
not ( n27786 , n27785 );
not ( n27787 , n11561 );
not ( n27788 , n27615 );
or ( n27789 , n27787 , n27788 );
not ( n27790 , n27615 );
nand ( n27791 , n27790 , n11558 );
nand ( n27792 , n27789 , n27791 );
xnor ( n27793 , n27792 , n11503 );
not ( n27794 , n27793 );
not ( n27795 , n27794 );
and ( n27796 , n27786 , n27795 );
and ( n27797 , n27785 , n27794 );
nor ( n27798 , n27796 , n27797 );
xor ( n27799 , n27760 , n27798 );
not ( n27800 , n26593 );
not ( n27801 , n14358 );
not ( n27802 , n13087 );
or ( n27803 , n27801 , n27802 );
not ( n27804 , n14358 );
nand ( n27805 , n27804 , n26602 );
nand ( n27806 , n27803 , n27805 );
not ( n27807 , n27806 );
or ( n27808 , n27800 , n27807 );
or ( n27809 , n27806 , n27419 );
nand ( n27810 , n27808 , n27809 );
not ( n27811 , n13502 );
not ( n27812 , n24913 );
not ( n27813 , n27812 );
not ( n27814 , n22100 );
or ( n27815 , n27813 , n27814 );
nand ( n27816 , n22095 , n24913 );
nand ( n27817 , n27815 , n27816 );
not ( n27818 , n27817 );
or ( n27819 , n27811 , n27818 );
not ( n27820 , n13502 );
not ( n27821 , n27820 );
or ( n27822 , n27817 , n27821 );
nand ( n27823 , n27819 , n27822 );
not ( n27824 , n27823 );
nand ( n27825 , n27810 , n27824 );
not ( n27826 , n27825 );
not ( n27827 , n20320 );
not ( n27828 , n9598 );
or ( n27829 , n27827 , n27828 );
or ( n27830 , n9598 , n20320 );
nand ( n27831 , n27829 , n27830 );
and ( n27832 , n27831 , n9650 );
not ( n27833 , n27831 );
and ( n27834 , n27833 , n9644 );
nor ( n27835 , n27832 , n27834 );
not ( n27836 , n27835 );
not ( n27837 , n27836 );
and ( n27838 , n27826 , n27837 );
and ( n27839 , n27825 , n27836 );
nor ( n27840 , n27838 , n27839 );
not ( n27841 , n27840 );
not ( n27842 , n27841 );
not ( n27843 , n8992 );
and ( n27844 , n8262 , n8258 );
not ( n27845 , n8262 );
not ( n27846 , n8257 );
and ( n27847 , n27845 , n27846 );
nor ( n27848 , n27844 , n27847 );
nor ( n27849 , n17345 , n27848 );
not ( n27850 , n27849 );
nand ( n27851 , n17345 , n27848 );
nand ( n27852 , n27850 , n27851 );
not ( n27853 , n27852 );
or ( n27854 , n27843 , n27853 );
or ( n27855 , n27852 , n7270 );
nand ( n27856 , n27854 , n27855 );
not ( n27857 , n27856 );
not ( n27858 , n7921 );
not ( n27859 , n19773 );
or ( n27860 , n27858 , n27859 );
not ( n27861 , n7921 );
nand ( n27862 , n27861 , n10270 );
nand ( n27863 , n27860 , n27862 );
and ( n27864 , n27863 , n10314 );
not ( n27865 , n27863 );
and ( n27866 , n27865 , n10311 );
nor ( n27867 , n27864 , n27866 );
nand ( n27868 , n27857 , n27867 );
not ( n27869 , n14527 );
not ( n27870 , n18028 );
or ( n27871 , n27869 , n27870 );
not ( n27872 , n14527 );
nand ( n27873 , n27872 , n12010 );
nand ( n27874 , n27871 , n27873 );
not ( n27875 , n27874 );
not ( n27876 , n12037 );
and ( n27877 , n27875 , n27876 );
and ( n27878 , n12037 , n27874 );
nor ( n27879 , n27877 , n27878 );
and ( n27880 , n27868 , n27879 );
not ( n27881 , n27868 );
not ( n27882 , n27879 );
and ( n27883 , n27881 , n27882 );
nor ( n27884 , n27880 , n27883 );
not ( n27885 , n27884 );
not ( n27886 , n27885 );
or ( n27887 , n27842 , n27886 );
nand ( n27888 , n27884 , n27840 );
nand ( n27889 , n27887 , n27888 );
and ( n27890 , n27799 , n27889 );
not ( n27891 , n27799 );
not ( n27892 , n27889 );
and ( n27893 , n27891 , n27892 );
nor ( n27894 , n27890 , n27893 );
buf ( n27895 , n27894 );
not ( n27896 , n27895 );
buf ( n27897 , n10337 );
not ( n27898 , n27897 );
not ( n27899 , n10346 );
not ( n27900 , n16158 );
and ( n27901 , n27899 , n27900 );
and ( n27902 , n10346 , n16158 );
nor ( n27903 , n27901 , n27902 );
not ( n27904 , n27903 );
and ( n27905 , n27898 , n27904 );
and ( n27906 , n27897 , n27903 );
nor ( n27907 , n27905 , n27906 );
not ( n27908 , n19471 );
and ( n27909 , n27907 , n27908 );
not ( n27910 , n27907 );
and ( n27911 , n27910 , n19471 );
nor ( n27912 , n27909 , n27911 );
not ( n27913 , n27912 );
not ( n27914 , n27913 );
buf ( n27915 , n9418 );
not ( n27916 , n27915 );
not ( n27917 , n8785 );
or ( n27918 , n27916 , n27917 );
or ( n27919 , n8785 , n27915 );
nand ( n27920 , n27918 , n27919 );
xor ( n27921 , n27920 , n8841 );
not ( n27922 , n14155 );
not ( n27923 , n26936 );
or ( n27924 , n27922 , n27923 );
or ( n27925 , n26936 , n14155 );
nand ( n27926 , n27924 , n27925 );
and ( n27927 , n27926 , n15521 );
not ( n27928 , n27926 );
and ( n27929 , n27928 , n15518 );
nor ( n27930 , n27927 , n27929 );
not ( n27931 , n27930 );
nand ( n27932 , n27921 , n27931 );
not ( n27933 , n27932 );
or ( n27934 , n27914 , n27933 );
nand ( n27935 , n27921 , n27931 );
or ( n27936 , n27935 , n27913 );
nand ( n27937 , n27934 , n27936 );
not ( n27938 , n27937 );
not ( n27939 , n18930 );
not ( n27940 , n13457 );
or ( n27941 , n27939 , n27940 );
or ( n27942 , n13457 , n18930 );
nand ( n27943 , n27941 , n27942 );
and ( n27944 , n27943 , n20866 );
not ( n27945 , n27943 );
buf ( n27946 , n13838 );
and ( n27947 , n27945 , n27946 );
nor ( n27948 , n27944 , n27947 );
not ( n27949 , n27948 );
not ( n27950 , n13239 );
not ( n27951 , n14797 );
or ( n27952 , n27950 , n27951 );
not ( n27953 , n14792 );
or ( n27954 , n27953 , n13239 );
nand ( n27955 , n27952 , n27954 );
and ( n27956 , n27955 , n14847 );
not ( n27957 , n27955 );
and ( n27958 , n27957 , n14840 );
nor ( n27959 , n27956 , n27958 );
nand ( n27960 , n27949 , n27959 );
not ( n27961 , n7381 );
not ( n27962 , n18260 );
or ( n27963 , n27961 , n27962 );
or ( n27964 , n18260 , n7381 );
nand ( n27965 , n27963 , n27964 );
and ( n27966 , n27965 , n22046 );
not ( n27967 , n27965 );
not ( n27968 , n22842 );
and ( n27969 , n27967 , n27968 );
nor ( n27970 , n27966 , n27969 );
not ( n27971 , n27970 );
and ( n27972 , n27960 , n27971 );
not ( n27973 , n27960 );
and ( n27974 , n27973 , n27970 );
nor ( n27975 , n27972 , n27974 );
not ( n27976 , n27975 );
nand ( n27977 , n27912 , n27930 );
not ( n27978 , n27977 );
not ( n27979 , n20651 );
not ( n27980 , n23122 );
or ( n27981 , n27979 , n27980 );
nand ( n27982 , n23121 , n20647 );
nand ( n27983 , n27981 , n27982 );
not ( n27984 , n27983 );
not ( n27985 , n23109 );
not ( n27986 , n27985 );
or ( n27987 , n27984 , n27986 );
or ( n27988 , n27985 , n27983 );
nand ( n27989 , n27987 , n27988 );
and ( n27990 , n27989 , n20410 );
not ( n27991 , n27989 );
not ( n27992 , n24001 );
not ( n27993 , n27992 );
and ( n27994 , n27991 , n27993 );
nor ( n27995 , n27990 , n27994 );
not ( n27996 , n27995 );
and ( n27997 , n27978 , n27996 );
and ( n27998 , n27977 , n27995 );
nor ( n27999 , n27997 , n27998 );
not ( n28000 , n27999 );
and ( n28001 , n27976 , n28000 );
and ( n28002 , n27975 , n27999 );
nor ( n28003 , n28001 , n28002 );
not ( n28004 , n28003 );
not ( n28005 , n28004 );
not ( n28006 , n11018 );
not ( n28007 , n9731 );
or ( n28008 , n28006 , n28007 );
or ( n28009 , n9731 , n11018 );
nand ( n28010 , n28008 , n28009 );
and ( n28011 , n28010 , n25248 );
not ( n28012 , n28010 );
and ( n28013 , n28012 , n25258 );
nor ( n28014 , n28011 , n28013 );
not ( n28015 , n24904 );
not ( n28016 , n22100 );
or ( n28017 , n28015 , n28016 );
or ( n28018 , n22096 , n24904 );
nand ( n28019 , n28017 , n28018 );
not ( n28020 , n28019 );
not ( n28021 , n27821 );
and ( n28022 , n28020 , n28021 );
and ( n28023 , n28019 , n27821 );
nor ( n28024 , n28022 , n28023 );
not ( n28025 , n28024 );
nand ( n28026 , n28014 , n28025 );
not ( n28027 , n12823 );
not ( n28028 , n9322 );
or ( n28029 , n28027 , n28028 );
or ( n28030 , n9322 , n12823 );
nand ( n28031 , n28029 , n28030 );
buf ( n28032 , n9374 );
and ( n28033 , n28031 , n28032 );
not ( n28034 , n28031 );
not ( n28035 , n28032 );
and ( n28036 , n28034 , n28035 );
nor ( n28037 , n28033 , n28036 );
and ( n28038 , n28026 , n28037 );
not ( n28039 , n28026 );
not ( n28040 , n28037 );
and ( n28041 , n28039 , n28040 );
nor ( n28042 , n28038 , n28041 );
not ( n28043 , n28042 );
not ( n28044 , n28043 );
or ( n28045 , n28005 , n28044 );
nand ( n28046 , n28003 , n28042 );
nand ( n28047 , n28045 , n28046 );
not ( n28048 , n21429 );
not ( n28049 , n18166 );
or ( n28050 , n28048 , n28049 );
or ( n28051 , n18166 , n21429 );
nand ( n28052 , n28050 , n28051 );
not ( n28053 , n28052 );
not ( n28054 , n7993 );
and ( n28055 , n28053 , n28054 );
and ( n28056 , n28052 , n23384 );
nor ( n28057 , n28055 , n28056 );
not ( n28058 , n28057 );
not ( n28059 , n16071 );
not ( n28060 , n18015 );
or ( n28061 , n28059 , n28060 );
or ( n28062 , n18015 , n16071 );
nand ( n28063 , n28061 , n28062 );
and ( n28064 , n28063 , n26425 );
not ( n28065 , n28063 );
and ( n28066 , n28065 , n20232 );
nor ( n28067 , n28064 , n28066 );
nand ( n28068 , n28058 , n28067 );
not ( n28069 , n28068 );
not ( n28070 , n15655 );
not ( n28071 , n26262 );
or ( n28072 , n28070 , n28071 );
nand ( n28073 , n26265 , n15651 );
nand ( n28074 , n28072 , n28073 );
and ( n28075 , n28074 , n26270 );
not ( n28076 , n28074 );
and ( n28077 , n28076 , n26269 );
nor ( n28078 , n28075 , n28077 );
not ( n28079 , n28078 );
and ( n28080 , n28069 , n28079 );
and ( n28081 , n28068 , n28078 );
nor ( n28082 , n28080 , n28081 );
not ( n28083 , n28082 );
xor ( n28084 , n13880 , n17546 );
buf ( n28085 , n19689 );
xnor ( n28086 , n28084 , n28085 );
not ( n28087 , n28086 );
not ( n28088 , n14383 );
not ( n28089 , n26593 );
or ( n28090 , n28088 , n28089 );
or ( n28091 , n26593 , n14383 );
nand ( n28092 , n28090 , n28091 );
and ( n28093 , n28092 , n26708 );
not ( n28094 , n28092 );
and ( n28095 , n28094 , n26712 );
nor ( n28096 , n28093 , n28095 );
nand ( n28097 , n28087 , n28096 );
not ( n28098 , n26321 );
not ( n28099 , n6854 );
not ( n28100 , n14447 );
or ( n28101 , n28099 , n28100 );
or ( n28102 , n14449 , n6854 );
nand ( n28103 , n28101 , n28102 );
not ( n28104 , n28103 );
or ( n28105 , n28098 , n28104 );
or ( n28106 , n28103 , n26321 );
nand ( n28107 , n28105 , n28106 );
not ( n28108 , n28107 );
and ( n28109 , n28097 , n28108 );
not ( n28110 , n28097 );
and ( n28111 , n28110 , n28107 );
nor ( n28112 , n28109 , n28111 );
not ( n28113 , n28112 );
or ( n28114 , n28083 , n28113 );
not ( n28115 , n28082 );
not ( n28116 , n28112 );
nand ( n28117 , n28115 , n28116 );
nand ( n28118 , n28114 , n28117 );
and ( n28119 , n28047 , n28118 );
not ( n28120 , n28047 );
not ( n28121 , n28118 );
and ( n28122 , n28120 , n28121 );
nor ( n28123 , n28119 , n28122 );
not ( n28124 , n28123 );
not ( n28125 , n28124 );
or ( n28126 , n27938 , n28125 );
not ( n28127 , n27937 );
and ( n28128 , n28047 , n28118 );
not ( n28129 , n28047 );
and ( n28130 , n28129 , n28121 );
nor ( n28131 , n28128 , n28130 );
nand ( n28132 , n28127 , n28131 );
nand ( n28133 , n28126 , n28132 );
not ( n28134 , n28133 );
or ( n28135 , n27896 , n28134 );
or ( n28136 , n28133 , n27895 );
nand ( n28137 , n28135 , n28136 );
not ( n28138 , n28137 );
nand ( n28139 , n27685 , n28138 );
or ( n28140 , n27661 , n28139 );
not ( n28141 , n27685 );
not ( n28142 , n27659 );
or ( n28143 , n28141 , n28142 );
buf ( n28144 , n15324 );
nor ( n28145 , n28138 , n28144 );
nand ( n28146 , n28143 , n28145 );
buf ( n28147 , n13353 );
nand ( n28148 , n28147 , n7566 );
nand ( n28149 , n28140 , n28146 , n28148 );
buf ( n28150 , n28149 );
buf ( n28151 , n28150 );
endmodule

