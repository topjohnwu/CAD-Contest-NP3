//
// Conformal-LEC Version 16.10-d160 ( 04-Jul-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 ;
output n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 ;

wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , 
     n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , 
     n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , 
     n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , 
     n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , 
     n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , 
     n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , 
     n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , 
     n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , 
     n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , 
     n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , 
     n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , 
     n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , 
     n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , 
     n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , 
     n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , 
     n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , 
     n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , 
     n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , 
     n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , 
     n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , 
     n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , 
     n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , 
     n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , 
     n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , 
     n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , 
     n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , 
     n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , 
     n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , 
     n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , 
     n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 ;
buf ( n62 , n320 );
buf ( n66 , n325 );
buf ( n63 , n334 );
buf ( n67 , n338 );
buf ( n60 , n343 );
buf ( n59 , n359 );
buf ( n58 , n371 );
buf ( n65 , n390 );
buf ( n64 , n408 );
buf ( n61 , n443 );
buf ( n185 , n44 );
buf ( n186 , n24 );
buf ( n187 , n43 );
buf ( n188 , n37 );
buf ( n189 , n3 );
buf ( n190 , n36 );
buf ( n191 , n25 );
buf ( n192 , n8 );
buf ( n193 , n34 );
buf ( n194 , n56 );
buf ( n195 , n48 );
buf ( n196 , n13 );
buf ( n197 , n1 );
buf ( n198 , n19 );
buf ( n199 , n50 );
buf ( n200 , n5 );
buf ( n201 , n6 );
buf ( n202 , n9 );
buf ( n203 , n4 );
buf ( n204 , n27 );
buf ( n205 , n38 );
buf ( n206 , n14 );
buf ( n207 , n22 );
buf ( n208 , n35 );
buf ( n209 , n41 );
buf ( n210 , n45 );
buf ( n211 , n26 );
buf ( n212 , n33 );
buf ( n213 , n15 );
buf ( n214 , n49 );
buf ( n215 , n16 );
buf ( n216 , n0 );
buf ( n217 , n21 );
buf ( n218 , n42 );
buf ( n219 , n18 );
buf ( n220 , n29 );
buf ( n221 , n23 );
buf ( n222 , n40 );
buf ( n223 , n57 );
buf ( n224 , n28 );
buf ( n225 , n51 );
buf ( n226 , n2 );
buf ( n227 , n46 );
buf ( n228 , n12 );
buf ( n229 , n31 );
buf ( n230 , n55 );
buf ( n231 , n54 );
buf ( n232 , n52 );
buf ( n233 , n39 );
buf ( n234 , n20 );
buf ( n235 , n32 );
buf ( n236 , n10 );
buf ( n237 , n7 );
buf ( n238 , n11 );
buf ( n239 , n30 );
buf ( n240 , n17 );
buf ( n241 , n47 );
buf ( n242 , n53 );
nor ( n243 , n210 , n211 , n212 , n213 );
not ( n244 , n243 );
and ( n245 , n244 , n185 );
not ( n246 , n220 );
not ( n247 , n215 );
not ( n248 , n185 );
not ( n249 , n208 );
and ( n250 , n188 , n189 , n190 , n191 );
and ( n251 , n187 , n250 );
not ( n252 , n188 );
and ( n253 , n252 , n189 , n190 , n191 );
and ( n254 , n192 , n253 );
not ( n255 , n189 );
and ( n256 , n188 , n255 , n190 , n191 );
and ( n257 , n193 , n256 );
and ( n258 , n252 , n255 , n190 , n191 );
and ( n259 , n194 , n258 );
not ( n260 , n190 );
and ( n261 , n188 , n189 , n260 , n191 );
and ( n262 , n195 , n261 );
and ( n263 , n252 , n189 , n260 , n191 );
and ( n264 , n196 , n263 );
and ( n265 , n188 , n255 , n260 , n191 );
and ( n266 , n197 , n265 );
and ( n267 , n252 , n255 , n260 , n191 );
and ( n268 , n198 , n267 );
nor ( n269 , n252 , n255 , n260 , n191 );
and ( n270 , n199 , n269 );
nor ( n271 , n188 , n255 , n260 , n191 );
and ( n272 , n200 , n271 );
nor ( n273 , n252 , n189 , n260 , n191 );
and ( n274 , n201 , n273 );
nor ( n275 , n188 , n189 , n260 , n191 );
and ( n276 , n202 , n275 );
nor ( n277 , n252 , n255 , n190 , n191 );
and ( n278 , n203 , n277 );
nor ( n279 , n188 , n255 , n190 , n191 );
and ( n280 , n204 , n279 );
nor ( n281 , n252 , n189 , n190 , n191 );
and ( n282 , n205 , n281 );
nor ( n283 , n188 , n189 , n190 , n191 );
and ( n284 , n206 , n283 );
or ( n285 , n251 , n254 , n257 , n259 , n262 , n264 , n266 , n268 , n270 , n272 , n274 , n276 , n278 , n280 , n282 , n284 );
and ( n286 , n249 , n285 );
and ( n287 , n207 , n208 );
or ( n288 , n286 , n287 );
xor ( n289 , n248 , n288 );
xor ( n290 , n186 , n289 );
and ( n291 , n210 , n211 , n212 , n213 );
not ( n292 , n291 );
and ( n293 , n292 , n209 );
and ( n294 , n248 , n291 );
or ( n295 , n293 , n294 );
xor ( n296 , n290 , n295 );
and ( n297 , n247 , n296 );
and ( n298 , n214 , n215 );
or ( n299 , n297 , n298 );
and ( n300 , n246 , n299 );
not ( n301 , n215 );
xor ( n302 , n185 , n217 );
xor ( n303 , n216 , n302 );
not ( n304 , n291 );
and ( n305 , n304 , n218 );
and ( n306 , n185 , n291 );
or ( n307 , n305 , n306 );
xor ( n308 , n303 , n307 );
and ( n309 , n301 , n308 );
and ( n310 , n219 , n215 );
or ( n311 , n309 , n310 );
not ( n312 , n311 );
and ( n313 , n312 , n220 );
or ( n314 , n300 , n313 );
and ( n315 , n314 , n243 );
or ( n316 , n245 , n315 );
not ( n317 , n221 );
and ( n318 , n316 , n317 );
buf ( n319 , n318 );
buf ( n320 , n319 );
not ( n321 , n221 );
and ( n322 , n321 , n299 );
or ( n323 , n322 , 1'b0 );
buf ( n324 , n323 );
buf ( n325 , n324 );
and ( n326 , n186 , n289 );
and ( n327 , n186 , n295 );
or ( n328 , n326 , n327 );
and ( n329 , n289 , n295 );
or ( n330 , n328 , n329 );
not ( n331 , n221 );
and ( n332 , n330 , n331 );
buf ( n333 , n332 );
buf ( n334 , n333 );
not ( n335 , n221 );
and ( n336 , n288 , n335 );
buf ( n337 , n336 );
buf ( n338 , n337 );
not ( n339 , n221 );
and ( n340 , n339 , n311 );
or ( n341 , n340 , 1'b0 );
buf ( n342 , n341 );
buf ( n343 , n342 );
not ( n344 , n221 );
not ( n345 , n243 );
and ( n346 , n345 , n222 );
buf ( n347 , n273 );
buf ( n348 , n275 );
buf ( n349 , n277 );
buf ( n350 , n279 );
buf ( n351 , n281 );
buf ( n352 , n283 );
or ( n353 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , n347 , n348 , n349 , n350 , n351 , n352 , 1'b0 );
and ( n354 , n353 , n243 );
or ( n355 , n346 , n354 );
and ( n356 , n344 , n355 );
or ( n357 , n356 , 1'b0 );
buf ( n358 , n357 );
buf ( n359 , n358 );
not ( n360 , n221 );
not ( n361 , n243 );
and ( n362 , n361 , n223 );
buf ( n363 , n283 );
buf ( n364 , n256 );
or ( n365 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , n363 , n364 );
and ( n366 , n365 , n243 );
or ( n367 , n362 , n366 );
and ( n368 , n360 , n367 );
or ( n369 , n368 , 1'b0 );
buf ( n370 , n369 );
buf ( n371 , n370 );
not ( n372 , n221 );
not ( n373 , n243 );
and ( n374 , n373 , n224 );
buf ( n375 , n265 );
buf ( n376 , n267 );
buf ( n377 , n269 );
buf ( n378 , n271 );
buf ( n379 , n273 );
buf ( n380 , n275 );
buf ( n381 , n277 );
buf ( n382 , n281 );
buf ( n383 , n283 );
or ( n384 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , 1'b0 , n382 , n383 , 1'b0 );
and ( n385 , n384 , n243 );
or ( n386 , n374 , n385 );
and ( n387 , n372 , n386 );
or ( n388 , n387 , 1'b0 );
buf ( n389 , n388 );
buf ( n390 , n389 );
not ( n391 , n221 );
not ( n392 , n243 );
and ( n393 , n392 , n225 );
buf ( n394 , n269 );
buf ( n395 , n271 );
buf ( n396 , n273 );
buf ( n397 , n275 );
buf ( n398 , n277 );
buf ( n399 , n279 );
buf ( n400 , n281 );
buf ( n401 , n283 );
or ( n402 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , 1'b0 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , 1'b0 );
and ( n403 , n402 , n243 );
or ( n404 , n393 , n403 );
and ( n405 , n391 , n404 );
or ( n406 , n405 , 1'b0 );
buf ( n407 , n406 );
buf ( n408 , n407 );
not ( n409 , n208 );
and ( n410 , n226 , n250 );
and ( n411 , n227 , n253 );
and ( n412 , n228 , n256 );
and ( n413 , n229 , n258 );
and ( n414 , n230 , n261 );
and ( n415 , n231 , n263 );
and ( n416 , n232 , n265 );
and ( n417 , n233 , n267 );
and ( n418 , n234 , n269 );
and ( n419 , n235 , n271 );
and ( n420 , n236 , n273 );
and ( n421 , n237 , n275 );
and ( n422 , n238 , n277 );
and ( n423 , n239 , n279 );
and ( n424 , n240 , n281 );
and ( n425 , n186 , n283 );
or ( n426 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 );
and ( n427 , n409 , n426 );
and ( n428 , n241 , n208 );
or ( n429 , n427 , n428 );
xor ( n430 , n185 , n429 );
and ( n431 , n206 , n430 );
not ( n432 , n291 );
and ( n433 , n432 , n242 );
and ( n434 , n185 , n291 );
or ( n435 , n433 , n434 );
and ( n436 , n206 , n435 );
or ( n437 , n431 , n436 );
and ( n438 , n430 , n435 );
or ( n439 , n437 , n438 );
not ( n440 , n221 );
and ( n441 , n439 , n440 );
buf ( n442 , n441 );
buf ( n443 , n442 );
endmodule

