//
// Conformal-LEC Version 15.20-d227 ( 10-Mar-2016) ( 64 bit executable)
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 ;
output n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;

wire n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , 
     n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , 
     n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , 
     n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , 
     n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , 
     n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , 
     n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , 
     n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , 
     n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , 
     n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , 
     n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , 
     n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , 
     n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , 
     n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , 
     n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , 
     n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , 
     n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , 
     n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , 
     n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , 
     n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , 
     n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , 
     n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , 
     n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , 
     n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , 
     n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , 
     n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , 
     n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , 
     n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , 
     n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , 
     n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , 
     n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , 
     n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , 
     n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , 
     n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , 
     n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , 
     n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , 
     n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , 
     n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , 
     n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , 
     n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , 
     n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , 
     n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , 
     n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , 
     n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , 
     n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , 
     n513 , n514 , n515 , n516 , n517 , n518 , n519 ;
buf ( n17 , n474 );
buf ( n28 , n477 );
buf ( n20 , n480 );
buf ( n26 , n483 );
buf ( n30 , n486 );
buf ( n25 , n489 );
buf ( n19 , n492 );
buf ( n16 , n495 );
buf ( n18 , n498 );
buf ( n21 , n501 );
buf ( n22 , n504 );
buf ( n31 , n507 );
buf ( n24 , n510 );
buf ( n29 , n513 );
buf ( n27 , n516 );
buf ( n23 , n519 );
buf ( n66 , n14 );
buf ( n67 , n11 );
buf ( n68 , n13 );
buf ( n69 , n10 );
buf ( n70 , n3 );
buf ( n71 , n12 );
buf ( n72 , n5 );
buf ( n73 , n8 );
buf ( n74 , n0 );
buf ( n75 , n7 );
buf ( n76 , n15 );
buf ( n77 , n2 );
buf ( n78 , n9 );
buf ( n79 , n4 );
buf ( n80 , n6 );
buf ( n81 , n1 );
buf ( n82 , n66 );
buf ( n83 , n74 );
and ( n84 , n82 , n83 );
buf ( n85 , n69 );
not ( n86 , n85 );
not ( n87 , n83 );
and ( n88 , n87 , n85 );
nor ( n89 , n86 , n88 );
buf ( n90 , n68 );
buf ( n91 , n75 );
and ( n92 , n90 , n91 );
and ( n93 , n89 , n92 );
buf ( n94 , n67 );
buf ( n95 , n76 );
and ( n96 , n94 , n95 );
and ( n97 , n92 , n96 );
and ( n98 , n89 , n96 );
or ( n99 , n93 , n97 , n98 );
not ( n100 , n90 );
and ( n101 , n87 , n90 );
nor ( n102 , n100 , n101 );
and ( n103 , n99 , n102 );
and ( n104 , n94 , n91 );
and ( n105 , n102 , n104 );
and ( n106 , n99 , n104 );
or ( n107 , n103 , n105 , n106 );
not ( n108 , n94 );
and ( n109 , n87 , n94 );
nor ( n110 , n108 , n109 );
and ( n111 , n107 , n110 );
not ( n112 , n82 );
and ( n113 , n112 , n91 );
not ( n114 , n91 );
nor ( n115 , n113 , n114 );
and ( n116 , n110 , n115 );
and ( n117 , n107 , n115 );
or ( n118 , n111 , n116 , n117 );
and ( n119 , n84 , n118 );
xor ( n120 , n84 , n118 );
xor ( n121 , n107 , n110 );
xor ( n122 , n121 , n115 );
buf ( n123 , n70 );
not ( n124 , n123 );
and ( n125 , n87 , n123 );
nor ( n126 , n124 , n125 );
and ( n127 , n85 , n91 );
and ( n128 , n126 , n127 );
buf ( n129 , n78 );
and ( n130 , n112 , n129 );
not ( n131 , n129 );
nor ( n132 , n130 , n131 );
and ( n133 , n127 , n132 );
and ( n134 , n126 , n132 );
or ( n135 , n128 , n133 , n134 );
and ( n136 , n85 , n95 );
buf ( n137 , n77 );
and ( n138 , n90 , n137 );
and ( n139 , n136 , n138 );
and ( n140 , n94 , n129 );
and ( n141 , n138 , n140 );
and ( n142 , n136 , n140 );
or ( n143 , n139 , n141 , n142 );
and ( n144 , n90 , n95 );
and ( n145 , n143 , n144 );
and ( n146 , n94 , n137 );
and ( n147 , n144 , n146 );
and ( n148 , n143 , n146 );
or ( n149 , n145 , n147 , n148 );
and ( n150 , n135 , n149 );
xor ( n151 , n89 , n92 );
xor ( n152 , n151 , n96 );
and ( n153 , n149 , n152 );
and ( n154 , n135 , n152 );
or ( n155 , n150 , n153 , n154 );
and ( n156 , n112 , n95 );
not ( n157 , n95 );
nor ( n158 , n156 , n157 );
and ( n159 , n155 , n158 );
xor ( n160 , n99 , n102 );
xor ( n161 , n160 , n104 );
and ( n162 , n158 , n161 );
and ( n163 , n155 , n161 );
or ( n164 , n159 , n162 , n163 );
and ( n165 , n122 , n164 );
xor ( n166 , n122 , n164 );
xor ( n167 , n155 , n158 );
xor ( n168 , n167 , n161 );
and ( n169 , n85 , n137 );
and ( n170 , n90 , n129 );
and ( n171 , n169 , n170 );
buf ( n172 , n79 );
and ( n173 , n94 , n172 );
and ( n174 , n170 , n173 );
and ( n175 , n169 , n173 );
or ( n176 , n171 , n174 , n175 );
buf ( n177 , n71 );
and ( n178 , n177 , n91 );
and ( n179 , n123 , n95 );
and ( n180 , n178 , n179 );
and ( n181 , n176 , n180 );
xor ( n182 , n136 , n138 );
xor ( n183 , n182 , n140 );
and ( n184 , n180 , n183 );
and ( n185 , n176 , n183 );
or ( n186 , n181 , n184 , n185 );
xor ( n187 , n126 , n127 );
xor ( n188 , n187 , n132 );
and ( n189 , n186 , n188 );
xor ( n190 , n143 , n144 );
xor ( n191 , n190 , n146 );
and ( n192 , n188 , n191 );
and ( n193 , n186 , n191 );
or ( n194 , n189 , n192 , n193 );
and ( n195 , n112 , n137 );
not ( n196 , n137 );
nor ( n197 , n195 , n196 );
and ( n198 , n194 , n197 );
xor ( n199 , n135 , n149 );
xor ( n200 , n199 , n152 );
and ( n201 , n197 , n200 );
and ( n202 , n194 , n200 );
or ( n203 , n198 , n201 , n202 );
and ( n204 , n168 , n203 );
xor ( n205 , n168 , n203 );
xor ( n206 , n194 , n197 );
xor ( n207 , n206 , n200 );
not ( n208 , n177 );
and ( n209 , n87 , n177 );
nor ( n210 , n208 , n209 );
and ( n211 , n123 , n91 );
and ( n212 , n210 , n211 );
and ( n213 , n112 , n172 );
not ( n214 , n172 );
nor ( n215 , n213 , n214 );
and ( n216 , n211 , n215 );
and ( n217 , n210 , n215 );
or ( n218 , n212 , n216 , n217 );
and ( n219 , n85 , n129 );
and ( n220 , n90 , n172 );
and ( n221 , n219 , n220 );
buf ( n222 , n80 );
and ( n223 , n94 , n222 );
and ( n224 , n220 , n223 );
and ( n225 , n219 , n223 );
or ( n226 , n221 , n224 , n225 );
xor ( n227 , n169 , n170 );
xor ( n228 , n227 , n173 );
and ( n229 , n226 , n228 );
xor ( n230 , n178 , n179 );
and ( n231 , n228 , n230 );
and ( n232 , n226 , n230 );
or ( n233 , n229 , n231 , n232 );
xor ( n234 , n210 , n211 );
xor ( n235 , n234 , n215 );
and ( n236 , n233 , n235 );
xor ( n237 , n176 , n180 );
xor ( n238 , n237 , n183 );
and ( n239 , n235 , n238 );
and ( n240 , n233 , n238 );
or ( n241 , n236 , n239 , n240 );
and ( n242 , n218 , n241 );
xor ( n243 , n186 , n188 );
xor ( n244 , n243 , n191 );
and ( n245 , n241 , n244 );
and ( n246 , n218 , n244 );
or ( n247 , n242 , n245 , n246 );
and ( n248 , n207 , n247 );
xor ( n249 , n207 , n247 );
xor ( n250 , n218 , n241 );
xor ( n251 , n250 , n244 );
buf ( n252 , n72 );
and ( n253 , n252 , n91 );
and ( n254 , n177 , n95 );
and ( n255 , n253 , n254 );
and ( n256 , n123 , n137 );
and ( n257 , n254 , n256 );
and ( n258 , n253 , n256 );
or ( n259 , n255 , n257 , n258 );
not ( n260 , n252 );
and ( n261 , n87 , n252 );
nor ( n262 , n260 , n261 );
and ( n263 , n259 , n262 );
and ( n264 , n112 , n222 );
not ( n265 , n222 );
nor ( n266 , n264 , n265 );
and ( n267 , n262 , n266 );
and ( n268 , n259 , n266 );
or ( n269 , n263 , n267 , n268 );
and ( n270 , n85 , n172 );
and ( n271 , n90 , n222 );
and ( n272 , n270 , n271 );
buf ( n273 , n81 );
and ( n274 , n94 , n273 );
and ( n275 , n271 , n274 );
and ( n276 , n270 , n274 );
or ( n277 , n272 , n275 , n276 );
xor ( n278 , n253 , n254 );
xor ( n279 , n278 , n256 );
and ( n280 , n277 , n279 );
xor ( n281 , n219 , n220 );
xor ( n282 , n281 , n223 );
and ( n283 , n279 , n282 );
and ( n284 , n277 , n282 );
or ( n285 , n280 , n283 , n284 );
xor ( n286 , n259 , n262 );
xor ( n287 , n286 , n266 );
and ( n288 , n285 , n287 );
xor ( n289 , n226 , n228 );
xor ( n290 , n289 , n230 );
and ( n291 , n287 , n290 );
and ( n292 , n285 , n290 );
or ( n293 , n288 , n291 , n292 );
and ( n294 , n269 , n293 );
xor ( n295 , n233 , n235 );
xor ( n296 , n295 , n238 );
and ( n297 , n293 , n296 );
and ( n298 , n269 , n296 );
or ( n299 , n294 , n297 , n298 );
and ( n300 , n251 , n299 );
xor ( n301 , n251 , n299 );
xor ( n302 , n269 , n293 );
xor ( n303 , n302 , n296 );
buf ( n304 , n73 );
not ( n305 , n304 );
and ( n306 , n87 , n304 );
nor ( n307 , n305 , n306 );
and ( n308 , n112 , n273 );
not ( n309 , n273 );
nor ( n310 , n308 , n309 );
and ( n311 , n307 , n310 );
and ( n312 , n85 , n222 );
and ( n313 , n90 , n273 );
and ( n314 , n312 , n313 );
and ( n315 , n123 , n129 );
and ( n316 , n314 , n315 );
xor ( n317 , n270 , n271 );
xor ( n318 , n317 , n274 );
and ( n319 , n315 , n318 );
and ( n320 , n314 , n318 );
or ( n321 , n316 , n319 , n320 );
xor ( n322 , n277 , n279 );
xor ( n323 , n322 , n282 );
and ( n324 , n321 , n323 );
xor ( n325 , n307 , n310 );
and ( n326 , n323 , n325 );
and ( n327 , n321 , n325 );
or ( n328 , n324 , n326 , n327 );
and ( n329 , n311 , n328 );
xor ( n330 , n285 , n287 );
xor ( n331 , n330 , n290 );
and ( n332 , n328 , n331 );
and ( n333 , n311 , n331 );
or ( n334 , n329 , n332 , n333 );
and ( n335 , n303 , n334 );
xor ( n336 , n303 , n334 );
xor ( n337 , n311 , n328 );
xor ( n338 , n337 , n331 );
and ( n339 , n304 , n91 );
and ( n340 , n252 , n95 );
and ( n341 , n339 , n340 );
and ( n342 , n177 , n137 );
and ( n343 , n340 , n342 );
and ( n344 , n339 , n342 );
or ( n345 , n341 , n343 , n344 );
and ( n346 , n177 , n172 );
and ( n347 , n123 , n222 );
and ( n348 , n346 , n347 );
and ( n349 , n85 , n273 );
and ( n350 , n347 , n349 );
and ( n351 , n346 , n349 );
or ( n352 , n348 , n350 , n351 );
and ( n353 , n123 , n172 );
and ( n354 , n352 , n353 );
xor ( n355 , n312 , n313 );
and ( n356 , n353 , n355 );
and ( n357 , n352 , n355 );
or ( n358 , n354 , n356 , n357 );
xor ( n359 , n339 , n340 );
xor ( n360 , n359 , n342 );
and ( n361 , n358 , n360 );
xor ( n362 , n314 , n315 );
xor ( n363 , n362 , n318 );
and ( n364 , n360 , n363 );
and ( n365 , n358 , n363 );
or ( n366 , n361 , n364 , n365 );
and ( n367 , n345 , n366 );
xor ( n368 , n321 , n323 );
xor ( n369 , n368 , n325 );
and ( n370 , n366 , n369 );
and ( n371 , n345 , n369 );
or ( n372 , n367 , n370 , n371 );
and ( n373 , n338 , n372 );
xor ( n374 , n338 , n372 );
xor ( n375 , n345 , n366 );
xor ( n376 , n375 , n369 );
and ( n377 , n252 , n137 );
and ( n378 , n177 , n129 );
and ( n379 , n377 , n378 );
and ( n380 , n252 , n172 );
and ( n381 , n177 , n222 );
and ( n382 , n380 , n381 );
and ( n383 , n123 , n273 );
and ( n384 , n381 , n383 );
and ( n385 , n380 , n383 );
or ( n386 , n382 , n384 , n385 );
and ( n387 , n252 , n129 );
and ( n388 , n386 , n387 );
xor ( n389 , n346 , n347 );
xor ( n390 , n389 , n349 );
and ( n391 , n387 , n390 );
and ( n392 , n386 , n390 );
or ( n393 , n388 , n391 , n392 );
xor ( n394 , n377 , n378 );
and ( n395 , n393 , n394 );
xor ( n396 , n352 , n353 );
xor ( n397 , n396 , n355 );
and ( n398 , n394 , n397 );
and ( n399 , n393 , n397 );
or ( n400 , n395 , n398 , n399 );
and ( n401 , n379 , n400 );
xor ( n402 , n358 , n360 );
xor ( n403 , n402 , n363 );
and ( n404 , n400 , n403 );
and ( n405 , n379 , n403 );
or ( n406 , n401 , n404 , n405 );
and ( n407 , n376 , n406 );
xor ( n408 , n376 , n406 );
xor ( n409 , n379 , n400 );
xor ( n410 , n409 , n403 );
and ( n411 , n304 , n172 );
and ( n412 , n252 , n222 );
and ( n413 , n411 , n412 );
and ( n414 , n177 , n273 );
and ( n415 , n412 , n414 );
and ( n416 , n411 , n414 );
or ( n417 , n413 , n415 , n416 );
and ( n418 , n304 , n129 );
and ( n419 , n417 , n418 );
xor ( n420 , n380 , n381 );
xor ( n421 , n420 , n383 );
and ( n422 , n418 , n421 );
and ( n423 , n417 , n421 );
or ( n424 , n419 , n422 , n423 );
and ( n425 , n304 , n137 );
and ( n426 , n424 , n425 );
xor ( n427 , n386 , n387 );
xor ( n428 , n427 , n390 );
and ( n429 , n425 , n428 );
and ( n430 , n424 , n428 );
or ( n431 , n426 , n429 , n430 );
xor ( n432 , n393 , n394 );
xor ( n433 , n432 , n397 );
and ( n434 , n431 , n433 );
and ( n435 , n410 , n434 );
xor ( n436 , n410 , n434 );
and ( n437 , n304 , n95 );
xor ( n438 , n431 , n433 );
and ( n439 , n437 , n438 );
xor ( n440 , n437 , n438 );
xor ( n441 , n424 , n425 );
xor ( n442 , n441 , n428 );
xor ( n443 , n417 , n418 );
xor ( n444 , n443 , n421 );
xor ( n445 , n411 , n412 );
xor ( n446 , n445 , n414 );
and ( n447 , n304 , n222 );
and ( n448 , n252 , n273 );
and ( n449 , n447 , n448 );
and ( n450 , n446 , n449 );
and ( n451 , n444 , n450 );
and ( n452 , n442 , n451 );
and ( n453 , n440 , n452 );
or ( n454 , n439 , n453 );
and ( n455 , n436 , n454 );
or ( n456 , n435 , n455 );
and ( n457 , n408 , n456 );
or ( n458 , n407 , n457 );
and ( n459 , n374 , n458 );
or ( n460 , n373 , n459 );
and ( n461 , n336 , n460 );
or ( n462 , n335 , n461 );
and ( n463 , n301 , n462 );
or ( n464 , n300 , n463 );
and ( n465 , n249 , n464 );
or ( n466 , n248 , n465 );
and ( n467 , n205 , n466 );
or ( n468 , n204 , n467 );
and ( n469 , n166 , n468 );
or ( n470 , n165 , n469 );
and ( n471 , n120 , n470 );
or ( n472 , n119 , n471 );
buf ( n473 , n472 );
buf ( n474 , n473 );
xor ( n475 , n120 , n470 );
buf ( n476 , n475 );
buf ( n477 , n476 );
xor ( n478 , n166 , n468 );
buf ( n479 , n478 );
buf ( n480 , n479 );
xor ( n481 , n205 , n466 );
buf ( n482 , n481 );
buf ( n483 , n482 );
xor ( n484 , n249 , n464 );
buf ( n485 , n484 );
buf ( n486 , n485 );
xor ( n487 , n301 , n462 );
buf ( n488 , n487 );
buf ( n489 , n488 );
xor ( n490 , n336 , n460 );
buf ( n491 , n490 );
buf ( n492 , n491 );
xor ( n493 , n374 , n458 );
buf ( n494 , n493 );
buf ( n495 , n494 );
xor ( n496 , n408 , n456 );
buf ( n497 , n496 );
buf ( n498 , n497 );
xor ( n499 , n436 , n454 );
buf ( n500 , n499 );
buf ( n501 , n500 );
xor ( n502 , n440 , n452 );
buf ( n503 , n502 );
buf ( n504 , n503 );
xor ( n505 , n442 , n451 );
buf ( n506 , n505 );
buf ( n507 , n506 );
xor ( n508 , n444 , n450 );
buf ( n509 , n508 );
buf ( n510 , n509 );
xor ( n511 , n446 , n449 );
buf ( n512 , n511 );
buf ( n513 , n512 );
xor ( n514 , n447 , n448 );
buf ( n515 , n514 );
buf ( n516 , n515 );
and ( n517 , n304 , n273 );
buf ( n518 , n517 );
buf ( n519 , n518 );
endmodule

