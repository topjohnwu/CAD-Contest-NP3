//
// Conformal-LEC Version 16.10-d160 ( 04-Jul-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ;
output n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ;

wire n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , 
     n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , 
     n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , 
     n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , 
     n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , 
     n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , 
     n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , 
     n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
     n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
     n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , 
     n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , 
     n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , 
     n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , 
     n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , 
     n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , 
     n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , 
     n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , 
     n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , 
     n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , 
     n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , 
     n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , 
     n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
     n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
     n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
     n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
     n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , 
     n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 ;
buf ( n39 , n203 );
buf ( n42 , n220 );
buf ( n35 , n237 );
buf ( n43 , n254 );
buf ( n40 , n271 );
buf ( n38 , n288 );
buf ( n34 , n305 );
buf ( n36 , n315 );
buf ( n37 , n334 );
buf ( n41 , n348 );
buf ( n125 , n0 );
buf ( n126 , n29 );
buf ( n127 , n7 );
buf ( n128 , n14 );
buf ( n129 , n24 );
buf ( n130 , n4 );
buf ( n131 , n21 );
buf ( n132 , n28 );
buf ( n133 , n13 );
buf ( n134 , n30 );
buf ( n135 , n10 );
buf ( n136 , n31 );
buf ( n137 , n3 );
buf ( n138 , n27 );
buf ( n139 , n6 );
buf ( n140 , n9 );
buf ( n141 , n11 );
buf ( n142 , n25 );
buf ( n143 , n8 );
buf ( n144 , n33 );
buf ( n145 , n2 );
buf ( n146 , n32 );
buf ( n147 , n18 );
buf ( n148 , n19 );
buf ( n149 , n15 );
buf ( n150 , n20 );
buf ( n151 , n26 );
buf ( n152 , n22 );
buf ( n153 , n23 );
buf ( n154 , n16 );
buf ( n155 , n17 );
buf ( n156 , n12 );
buf ( n157 , n5 );
not ( n158 , n155 );
not ( n159 , n146 );
not ( n160 , n147 );
not ( n161 , n148 );
not ( n162 , n149 );
not ( n163 , n151 );
not ( n164 , n152 );
nor ( n165 , n159 , n160 , n161 , n162 , n150 , n163 , n164 , n153 , n154 );
not ( n166 , n165 );
and ( n167 , n166 , n125 );
not ( n168 , n135 );
and ( n169 , n168 , n125 );
buf ( n170 , n125 );
buf ( n171 , n126 );
buf ( n172 , n127 );
buf ( n173 , n128 );
buf ( n174 , n129 );
buf ( n175 , n130 );
buf ( n176 , n131 );
buf ( n177 , n132 );
buf ( n178 , n133 );
buf ( n179 , n134 );
and ( n180 , n178 , n179 );
and ( n181 , n177 , n180 );
and ( n182 , n176 , n181 );
and ( n183 , n175 , n182 );
and ( n184 , n174 , n183 );
and ( n185 , n173 , n184 );
and ( n186 , n172 , n185 );
and ( n187 , n171 , n186 );
xor ( n188 , n170 , n187 );
buf ( n189 , n188 );
and ( n190 , n189 , n135 );
or ( n191 , n169 , n190 );
not ( n192 , n138 );
not ( n193 , n139 );
not ( n194 , n145 );
or ( n195 , n136 , n137 , n192 , n193 , n140 , n141 , n142 , n143 , n144 , n194 );
and ( n196 , n191 , n195 );
or ( n197 , 1'b0 , n196 );
and ( n198 , n197 , n165 );
or ( n199 , n167 , n198 );
and ( n200 , n158 , n199 );
or ( n201 , n200 , 1'b0 );
buf ( n202 , n201 );
buf ( n203 , n202 );
not ( n204 , n155 );
not ( n205 , n165 );
and ( n206 , n205 , n126 );
not ( n207 , n135 );
and ( n208 , n207 , n126 );
xor ( n209 , n171 , n186 );
buf ( n210 , n209 );
and ( n211 , n210 , n135 );
or ( n212 , n208 , n211 );
and ( n213 , n212 , n195 );
or ( n214 , 1'b0 , n213 );
and ( n215 , n214 , n165 );
or ( n216 , n206 , n215 );
and ( n217 , n204 , n216 );
or ( n218 , n217 , 1'b0 );
buf ( n219 , n218 );
buf ( n220 , n219 );
not ( n221 , n155 );
not ( n222 , n165 );
and ( n223 , n222 , n127 );
not ( n224 , n135 );
and ( n225 , n224 , n127 );
xor ( n226 , n172 , n185 );
buf ( n227 , n226 );
and ( n228 , n227 , n135 );
or ( n229 , n225 , n228 );
and ( n230 , n229 , n195 );
or ( n231 , 1'b0 , n230 );
and ( n232 , n231 , n165 );
or ( n233 , n223 , n232 );
and ( n234 , n221 , n233 );
or ( n235 , n234 , 1'b0 );
buf ( n236 , n235 );
buf ( n237 , n236 );
not ( n238 , n155 );
not ( n239 , n165 );
and ( n240 , n239 , n128 );
not ( n241 , n135 );
and ( n242 , n241 , n128 );
xor ( n243 , n173 , n184 );
buf ( n244 , n243 );
and ( n245 , n244 , n135 );
or ( n246 , n242 , n245 );
and ( n247 , n246 , n195 );
or ( n248 , 1'b0 , n247 );
and ( n249 , n248 , n165 );
or ( n250 , n240 , n249 );
and ( n251 , n238 , n250 );
or ( n252 , n251 , 1'b0 );
buf ( n253 , n252 );
buf ( n254 , n253 );
not ( n255 , n155 );
not ( n256 , n165 );
and ( n257 , n256 , n129 );
not ( n258 , n135 );
and ( n259 , n258 , n129 );
xor ( n260 , n174 , n183 );
buf ( n261 , n260 );
and ( n262 , n261 , n135 );
or ( n263 , n259 , n262 );
and ( n264 , n263 , n195 );
or ( n265 , 1'b0 , n264 );
and ( n266 , n265 , n165 );
or ( n267 , n257 , n266 );
and ( n268 , n255 , n267 );
or ( n269 , n268 , 1'b0 );
buf ( n270 , n269 );
buf ( n271 , n270 );
not ( n272 , n155 );
not ( n273 , n165 );
and ( n274 , n273 , n130 );
not ( n275 , n135 );
and ( n276 , n275 , n130 );
xor ( n277 , n175 , n182 );
buf ( n278 , n277 );
and ( n279 , n278 , n135 );
or ( n280 , n276 , n279 );
and ( n281 , n280 , n195 );
or ( n282 , 1'b0 , n281 );
and ( n283 , n282 , n165 );
or ( n284 , n274 , n283 );
and ( n285 , n272 , n284 );
or ( n286 , n285 , 1'b0 );
buf ( n287 , n286 );
buf ( n288 , n287 );
not ( n289 , n155 );
not ( n290 , n165 );
and ( n291 , n290 , n131 );
not ( n292 , n135 );
and ( n293 , n292 , n131 );
xor ( n294 , n176 , n181 );
buf ( n295 , n294 );
and ( n296 , n295 , n135 );
or ( n297 , n293 , n296 );
and ( n298 , n297 , n195 );
or ( n299 , 1'b0 , n298 );
and ( n300 , n299 , n165 );
or ( n301 , n291 , n300 );
and ( n302 , n289 , n301 );
or ( n303 , n302 , 1'b0 );
buf ( n304 , n303 );
buf ( n305 , n304 );
or ( n306 , n155 , n165 );
not ( n307 , n306 );
nor ( n308 , n159 , n160 , n161 , n162 , n150 , n151 , n152 , n153 , n154 );
not ( n309 , n308 );
and ( n310 , n156 , n309 );
and ( n311 , n307 , n310 );
and ( n312 , 1'b1 , n306 );
or ( n313 , n311 , n312 );
buf ( n314 , n313 );
buf ( n315 , n314 );
not ( n316 , n155 );
not ( n317 , n165 );
and ( n318 , n317 , n157 );
nor ( n319 , n136 , n137 , n192 , n193 , n140 , n141 , n142 , n143 , n144 , n145 );
not ( n320 , n319 );
not ( n321 , n137 );
nor ( n322 , n136 , n321 , n138 , n193 , n140 , n141 , n142 , n143 , n144 , n145 );
not ( n323 , n322 );
and ( n324 , n157 , n323 );
and ( n325 , n320 , n324 );
and ( n326 , 1'b1 , n319 );
or ( n327 , n325 , n326 );
and ( n328 , n327 , n165 );
or ( n329 , n318 , n328 );
and ( n330 , n316 , n329 );
and ( n331 , 1'b1 , n155 );
or ( n332 , n330 , n331 );
buf ( n333 , n332 );
buf ( n334 , n333 );
not ( n335 , n155 );
not ( n336 , n165 );
and ( n337 , n336 , n136 );
buf ( n338 , n136 );
not ( n339 , n338 );
buf ( n340 , n339 );
and ( n341 , n340 , n195 );
or ( n342 , 1'b0 , n341 );
and ( n343 , n342 , n165 );
or ( n344 , n337 , n343 );
and ( n345 , n335 , n344 );
or ( n346 , n345 , 1'b0 );
buf ( n347 , n346 );
buf ( n348 , n347 );
not ( n349 , n195 );
not ( n350 , n195 );
not ( n351 , n195 );
not ( n352 , n195 );
not ( n353 , n195 );
not ( n354 , n195 );
not ( n355 , n195 );
not ( n356 , n195 );
endmodule

