//
// Conformal-LEC Version 16.10-d005 ( 21-Apr-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 ;
output n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 ;

wire n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
     n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
     n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
     n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
     n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
     n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
     n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
     n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
     n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
     n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
     n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
     n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
     n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
     n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
     n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
     n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
     n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
     n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
     n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
     n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
     n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
     n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
     n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
     n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
     n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , 
     n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , 
     n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
     n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , 
     n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
     n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , 
     n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
     n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
     n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
     n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , 
     n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
     n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
     n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
     n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
     n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
     n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
     n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
     n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
     n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
     n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
     n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
     n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
     n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , 
     n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , 
     n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , 
     n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , 
     n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , 
     n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , 
     n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , 
     n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
     n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , 
     n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , 
     n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , 
     n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , 
     n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , 
     n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , 
     n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , 
     n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , 
     n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , 
     n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , 
     n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , 
     n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , 
     n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , 
     n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , 
     n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
     n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
     n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
     n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
     n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
     n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
     n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
     n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
     n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
     n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
     n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
     n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
     n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
     n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
     n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , 
     n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , 
     n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
     n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , 
     n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , 
     n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , 
     n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , 
     n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , 
     n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , 
     n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , 
     n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , 
     n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
     n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , 
     n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , 
     n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , 
     n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
     n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , 
     n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , 
     n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
     n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , 
     n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , 
     n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , 
     n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , 
     n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , 
     n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , 
     n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , 
     n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , 
     n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , 
     n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , 
     n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , 
     n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , 
     n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , 
     n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , 
     n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , 
     n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , 
     n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , 
     n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , 
     n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
     n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , 
     n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , 
     n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , 
     n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , 
     n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , 
     n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , 
     n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , 
     n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , 
     n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , 
     n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , 
     n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , 
     n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , 
     n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , 
     n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , 
     n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , 
     n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , 
     n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , 
     n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , 
     n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , 
     n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , 
     n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , 
     n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , 
     n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , 
     n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , 
     n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , 
     n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , 
     n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , 
     n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , 
     n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , 
     n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , 
     n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , 
     n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , 
     n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , 
     n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , 
     n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , 
     n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , 
     n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , 
     n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , 
     n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , 
     n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , 
     n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , 
     n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , 
     n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , 
     n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , 
     n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , 
     n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , 
     n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , 
     n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , 
     n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , 
     n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , 
     n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , 
     n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , 
     n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , 
     n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , 
     n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , 
     n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , 
     n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , 
     n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , 
     n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , 
     n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , 
     n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , 
     n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , 
     n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , 
     n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , 
     n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , 
     n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , 
     n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , 
     n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , 
     n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , 
     n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , 
     n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , 
     n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , 
     n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , 
     n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , 
     n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , 
     n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , 
     n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , 
     n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , 
     n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , 
     n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , 
     n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , 
     n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , 
     n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , 
     n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , 
     n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , 
     n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , 
     n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , 
     n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , 
     n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , 
     n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , 
     n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , 
     n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , 
     n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , 
     n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , 
     n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , 
     n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , 
     n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , 
     n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , 
     n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , 
     n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , 
     n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , 
     n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , 
     n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , 
     n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , 
     n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , 
     n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , 
     n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , 
     n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , 
     n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , 
     n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , 
     n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , 
     n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , 
     n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , 
     n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , 
     n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , 
     n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , 
     n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , 
     n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , 
     n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , 
     n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , 
     n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , 
     n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , 
     n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , 
     n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , 
     n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , 
     n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , 
     n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , 
     n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , 
     n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , 
     n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , 
     n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , 
     n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , 
     n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , 
     n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , 
     n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , 
     n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , 
     n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , 
     n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , 
     n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , 
     n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , 
     n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , 
     n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , 
     n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , 
     n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , 
     n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , 
     n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , 
     n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , 
     n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , 
     n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , 
     n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , 
     n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , 
     n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , 
     n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , 
     n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , 
     n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , 
     n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , 
     n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , 
     n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , 
     n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , 
     n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , 
     n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , 
     n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , 
     n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , 
     n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , 
     n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , 
     n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , 
     n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , 
     n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , 
     n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , 
     n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , 
     n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , 
     n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , 
     n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , 
     n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , 
     n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , 
     n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , 
     n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , 
     n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , 
     n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , 
     n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , 
     n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , 
     n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , 
     n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , 
     n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , 
     n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , 
     n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , 
     n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , 
     n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , 
     n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , 
     n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , 
     n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , 
     n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , 
     n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , 
     n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , 
     n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , 
     n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , 
     n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , 
     n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , 
     n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , 
     n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , 
     n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , 
     n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , 
     n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , 
     n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , 
     n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , 
     n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , 
     n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , 
     n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , 
     n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , 
     n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , 
     n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , 
     n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , 
     n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , 
     n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , 
     n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , 
     n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , 
     n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , 
     n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , 
     n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , 
     n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , 
     n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , 
     n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , 
     n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , 
     n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , 
     n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , 
     n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , 
     n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , 
     n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , 
     n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , 
     n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , 
     n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , 
     n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , 
     n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , 
     n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , 
     n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , 
     n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , 
     n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , 
     n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , 
     n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , 
     n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , 
     n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , 
     n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , 
     n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , 
     n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , 
     n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , 
     n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , 
     n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , 
     n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , 
     n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , 
     n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , 
     n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , 
     n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , 
     n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , 
     n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , 
     n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , 
     n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , 
     n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , 
     n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , 
     n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , 
     n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , 
     n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , 
     n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , 
     n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , 
     n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , 
     n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , 
     n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , 
     n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , 
     n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , 
     n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , 
     n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , 
     n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , 
     n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , 
     n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , 
     n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , 
     n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , 
     n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , 
     n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , 
     n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , 
     n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , 
     n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , 
     n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , 
     n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , 
     n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , 
     n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , 
     n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , 
     n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , 
     n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , 
     n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , 
     n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , 
     n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , 
     n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , 
     n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , 
     n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , 
     n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , 
     n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , 
     n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , 
     n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , 
     n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , 
     n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , 
     n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , 
     n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , 
     n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , 
     n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , 
     n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , 
     n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , 
     n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , 
     n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , 
     n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , 
     n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , 
     n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , 
     n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , 
     n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , 
     n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , 
     n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , 
     n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , 
     n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , 
     n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , 
     n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , 
     n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , 
     n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , 
     n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , 
     n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , 
     n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , 
     n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , 
     n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , 
     n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , 
     n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , 
     n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , 
     n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , 
     n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , 
     n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , 
     n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , 
     n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , 
     n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , 
     n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , 
     n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , 
     n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , 
     n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , 
     n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , 
     n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , 
     n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , 
     n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , 
     n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , 
     n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , 
     n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , 
     n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , 
     n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , 
     n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , 
     n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , 
     n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , 
     n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , 
     n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , 
     n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , 
     n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , 
     n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , 
     n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , 
     n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , 
     n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , 
     n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , 
     n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , 
     n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , 
     n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , 
     n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , 
     n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , 
     n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , 
     n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , 
     n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , 
     n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , 
     n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , 
     n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , 
     n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , 
     n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , 
     n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , 
     n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , 
     n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , 
     n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , 
     n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , 
     n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , 
     n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , 
     n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , 
     n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , 
     n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , 
     n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , 
     n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , 
     n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , 
     n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , 
     n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , 
     n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , 
     n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , 
     n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , 
     n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , 
     n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , 
     n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , 
     n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , 
     n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , 
     n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , 
     n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , 
     n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , 
     n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , 
     n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , 
     n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , 
     n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , 
     n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , 
     n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , 
     n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , 
     n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , 
     n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , 
     n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , 
     n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , 
     n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , 
     n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , 
     n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , 
     n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , 
     n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , 
     n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , 
     n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , 
     n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , 
     n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , 
     n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , 
     n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , 
     n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , 
     n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , 
     n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , 
     n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , 
     n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , 
     n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , 
     n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , 
     n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , 
     n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , 
     n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , 
     n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , 
     n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , 
     n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , 
     n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , 
     n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , 
     n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , 
     n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , 
     n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , 
     n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , 
     n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , 
     n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , 
     n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , 
     n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , 
     n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , 
     n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , 
     n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , 
     n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , 
     n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , 
     n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , 
     n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , 
     n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , 
     n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , 
     n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , 
     n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , 
     n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , 
     n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , 
     n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , 
     n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , 
     n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , 
     n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , 
     n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , 
     n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , 
     n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , 
     n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , 
     n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , 
     n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , 
     n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , 
     n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , 
     n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , 
     n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , 
     n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , 
     n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , 
     n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , 
     n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , 
     n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , 
     n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , 
     n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , 
     n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , 
     n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , 
     n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , 
     n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , 
     n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , 
     n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , 
     n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , 
     n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , 
     n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , 
     n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , 
     n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , 
     n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , 
     n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , 
     n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , 
     n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , 
     n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , 
     n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , 
     n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , 
     n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , 
     n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , 
     n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , 
     n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , 
     n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , 
     n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , 
     n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , 
     n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , 
     n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , 
     n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , 
     n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , 
     n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , 
     n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , 
     n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , 
     n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , 
     n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , 
     n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , 
     n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , 
     n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , 
     n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , 
     n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , 
     n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , 
     n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , 
     n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , 
     n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , 
     n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , 
     n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , 
     n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , 
     n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , 
     n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , 
     n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , 
     n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , 
     n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , 
     n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , 
     n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , 
     n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , 
     n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , 
     n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , 
     n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , 
     n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , 
     n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , 
     n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , 
     n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , 
     n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , 
     n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , 
     n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , 
     n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , 
     n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , 
     n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , 
     n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , 
     n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , 
     n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , 
     n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , 
     n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , 
     n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , 
     n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , 
     n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , 
     n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , 
     n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , 
     n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , 
     n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , 
     n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , 
     n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , 
     n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , 
     n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , 
     n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , 
     n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , 
     n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , 
     n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , 
     n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , 
     n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , 
     n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , 
     n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , 
     n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , 
     n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , 
     n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , 
     n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , 
     n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , 
     n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , 
     n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , 
     n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , 
     n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , 
     n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , 
     n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , 
     n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , 
     n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , 
     n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , 
     n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , 
     n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , 
     n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , 
     n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , 
     n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , 
     n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , 
     n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , 
     n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , 
     n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , 
     n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , 
     n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , 
     n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , 
     n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , 
     n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , 
     n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , 
     n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , 
     n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , 
     n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , 
     n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , 
     n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , 
     n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , 
     n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , 
     n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , 
     n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , 
     n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , 
     n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , 
     n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , 
     n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , 
     n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , 
     n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , 
     n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , 
     n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , 
     n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , 
     n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , 
     n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , 
     n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , 
     n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , 
     n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , 
     n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , 
     n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , 
     n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , 
     n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , 
     n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , 
     n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , 
     n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , 
     n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , 
     n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , 
     n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , 
     n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , 
     n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , 
     n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , 
     n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , 
     n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , 
     n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , 
     n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , 
     n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , 
     n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , 
     n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , 
     n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , 
     n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , 
     n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , 
     n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , 
     n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , 
     n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , 
     n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , 
     n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , 
     n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , 
     n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , 
     n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , 
     n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , 
     n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , 
     n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , 
     n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , 
     n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , 
     n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , 
     n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , 
     n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , 
     n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , 
     n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , 
     n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , 
     n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , 
     n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , 
     n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , 
     n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , 
     n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , 
     n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , 
     n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , 
     n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , 
     n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , 
     n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , 
     n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , 
     n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , 
     n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , 
     n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , 
     n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , 
     n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , 
     n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , 
     n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , 
     n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , 
     n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , 
     n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , 
     n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , 
     n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , 
     n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , 
     n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , 
     n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , 
     n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , 
     n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , 
     n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , 
     n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , 
     n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , 
     n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , 
     n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , 
     n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , 
     n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , 
     n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , 
     n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , 
     n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , 
     n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , 
     n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , 
     n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , 
     n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , 
     n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , 
     n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , 
     n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , 
     n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , 
     n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , 
     n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , 
     n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , 
     n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , 
     n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , 
     n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , 
     n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , 
     n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , 
     n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , 
     n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , 
     n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , 
     n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , 
     n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , 
     n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , 
     n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , 
     n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , 
     n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , 
     n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , 
     n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , 
     n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , 
     n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , 
     n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , 
     n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , 
     n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , 
     n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , 
     n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , 
     n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , 
     n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , 
     n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , 
     n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , 
     n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , 
     n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , 
     n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , 
     n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , 
     n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , 
     n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , 
     n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , 
     n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , 
     n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , 
     n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , 
     n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , 
     n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , 
     n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , 
     n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , 
     n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , 
     n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , 
     n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , 
     n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , 
     n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , 
     n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , 
     n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , 
     n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , 
     n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , 
     n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , 
     n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , 
     n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , 
     n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , 
     n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , 
     n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , 
     n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , 
     n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , 
     n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , 
     n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , 
     n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , 
     n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , 
     n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , 
     n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , 
     n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , 
     n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , 
     n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , 
     n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , 
     n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , 
     n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , 
     n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , 
     n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , 
     n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , 
     n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , 
     n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , 
     n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , 
     n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , 
     n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , 
     n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , 
     n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , 
     n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , 
     n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , 
     n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , 
     n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , 
     n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , 
     n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , 
     n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , 
     n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , 
     n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , 
     n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , 
     n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , 
     n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , 
     n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , 
     n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , 
     n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , 
     n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , 
     n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , 
     n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , 
     n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , 
     n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , 
     n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , 
     n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , 
     n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , 
     n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , 
     n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , 
     n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , 
     n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , 
     n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , 
     n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , 
     n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , 
     n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , 
     n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , 
     n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , 
     n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , 
     n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , 
     n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , 
     n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , 
     n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , 
     n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , 
     n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , 
     n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , 
     n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , 
     n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , 
     n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , 
     n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , 
     n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , 
     n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , 
     n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , 
     n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , 
     n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , 
     n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , 
     n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , 
     n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , 
     n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , 
     n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , 
     n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , 
     n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , 
     n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , 
     n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , 
     n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , 
     n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , 
     n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , 
     n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , 
     n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , 
     n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , 
     n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , 
     n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , 
     n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , 
     n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , 
     n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , 
     n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , 
     n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , 
     n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , 
     n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , 
     n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , 
     n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , 
     n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , 
     n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , 
     n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , 
     n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , 
     n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , 
     n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , 
     n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , 
     n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , 
     n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , 
     n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , 
     n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , 
     n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , 
     n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , 
     n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , 
     n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , 
     n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , 
     n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , 
     n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , 
     n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , 
     n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , 
     n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , 
     n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , 
     n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , 
     n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , 
     n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , 
     n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , 
     n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , 
     n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , 
     n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , 
     n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , 
     n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , 
     n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , 
     n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , 
     n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , 
     n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , 
     n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , 
     n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , 
     n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , 
     n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , 
     n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , 
     n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , 
     n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , 
     n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , 
     n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , 
     n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , 
     n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , 
     n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , 
     n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , 
     n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , 
     n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , 
     n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , 
     n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , 
     n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , 
     n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , 
     n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , 
     n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , 
     n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , 
     n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , 
     n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , 
     n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , 
     n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , 
     n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , 
     n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , 
     n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , 
     n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , 
     n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , 
     n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , 
     n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , 
     n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , 
     n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , 
     n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , 
     n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , 
     n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , 
     n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , 
     n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , 
     n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , 
     n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , 
     n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , 
     n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , 
     n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , 
     n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , 
     n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , 
     n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , 
     n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , 
     n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , 
     n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , 
     n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , 
     n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , 
     n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , 
     n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , 
     n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , 
     n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , 
     n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , 
     n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , 
     n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , 
     n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , 
     n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , 
     n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , 
     n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , 
     n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , 
     n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , 
     n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , 
     n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , 
     n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , 
     n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , 
     n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , 
     n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , 
     n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , 
     n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , 
     n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , 
     n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , 
     n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , 
     n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , 
     n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , 
     n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , 
     n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , 
     n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , 
     n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , 
     n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , 
     n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , 
     n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , 
     n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , 
     n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , 
     n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , 
     n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , 
     n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , 
     n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , 
     n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , 
     n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , 
     n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , 
     n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , 
     n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , 
     n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , 
     n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , 
     n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , 
     n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , 
     n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , 
     n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , 
     n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , 
     n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , 
     n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , 
     n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , 
     n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , 
     n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , 
     n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , 
     n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , 
     n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , 
     n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , 
     n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , 
     n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , 
     n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , 
     n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , 
     n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , 
     n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , 
     n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , 
     n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , 
     n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , 
     n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , 
     n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , 
     n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , 
     n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , 
     n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , 
     n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , 
     n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , 
     n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , 
     n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , 
     n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , 
     n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , 
     n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , 
     n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , 
     n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , 
     n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , 
     n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , 
     n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , 
     n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , 
     n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , 
     n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , 
     n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , 
     n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , 
     n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , 
     n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , 
     n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , 
     n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , 
     n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , 
     n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , 
     n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , 
     n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , 
     n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , 
     n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , 
     n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , 
     n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , 
     n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , 
     n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , 
     n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , 
     n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , 
     n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , 
     n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , 
     n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , 
     n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , 
     n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , 
     n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , 
     n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , 
     n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , 
     n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , 
     n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , 
     n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , 
     n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , 
     n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , 
     n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , 
     n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , 
     n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , 
     n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , 
     n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , 
     n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , 
     n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , 
     n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , 
     n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , 
     n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , 
     n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , 
     n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , 
     n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , 
     n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , 
     n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , 
     n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , 
     n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , 
     n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , 
     n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , 
     n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , 
     n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , 
     n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , 
     n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , 
     n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , 
     n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , 
     n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , 
     n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , 
     n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , 
     n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , 
     n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , 
     n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , 
     n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , 
     n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , 
     n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , 
     n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , 
     n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , 
     n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , 
     n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , 
     n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , 
     n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , 
     n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , 
     n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , 
     n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , 
     n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , 
     n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , 
     n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , 
     n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , 
     n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , 
     n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , 
     n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , 
     n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , 
     n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , 
     n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , 
     n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , 
     n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , 
     n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , 
     n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , 
     n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , 
     n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , 
     n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , 
     n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , 
     n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , 
     n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , 
     n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , 
     n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , 
     n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , 
     n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , 
     n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , 
     n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , 
     n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , 
     n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , 
     n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , 
     n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , 
     n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , 
     n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , 
     n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , 
     n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , 
     n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , 
     n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , 
     n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , 
     n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , 
     n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , 
     n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , 
     n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , 
     n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , 
     n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , 
     n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , 
     n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , 
     n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , 
     n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , 
     n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , 
     n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , 
     n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , 
     n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , 
     n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , 
     n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , 
     n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , 
     n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , 
     n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , 
     n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , 
     n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , 
     n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , 
     n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , 
     n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , 
     n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , 
     n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , 
     n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , 
     n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , 
     n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , 
     n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , 
     n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , 
     n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , 
     n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , 
     n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , 
     n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , 
     n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , 
     n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , 
     n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , 
     n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , 
     n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , 
     n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , 
     n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , 
     n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , 
     n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , 
     n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , 
     n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , 
     n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , 
     n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , 
     n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , 
     n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , 
     n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , 
     n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , 
     n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , 
     n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , 
     n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , 
     n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , 
     n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , 
     n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , 
     n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , 
     n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , 
     n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , 
     n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , 
     n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , 
     n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , 
     n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , 
     n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , 
     n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , 
     n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , 
     n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , 
     n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , 
     n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , 
     n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , 
     n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , 
     n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , 
     n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , 
     n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , 
     n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , 
     n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , 
     n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , 
     n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , 
     n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , 
     n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , 
     n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , 
     n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , 
     n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , 
     n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , 
     n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , 
     n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , 
     n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , 
     n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , 
     n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , 
     n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , 
     n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , 
     n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , 
     n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , 
     n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , 
     n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , 
     n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , 
     n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , 
     n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , 
     n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , 
     n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , 
     n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , 
     n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , 
     n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , 
     n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , 
     n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , 
     n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , 
     n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , 
     n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , 
     n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , 
     n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , 
     n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , 
     n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , 
     n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , 
     n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , 
     n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , 
     n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , 
     n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , 
     n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , 
     n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , 
     n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , 
     n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , 
     n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , 
     n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , 
     n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , 
     n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , 
     n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , 
     n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , 
     n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , 
     n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , 
     n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , 
     n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , 
     n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , 
     n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , 
     n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , 
     n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , 
     n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , 
     n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , 
     n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , 
     n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , 
     n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , 
     n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , 
     n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , 
     n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , 
     n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , 
     n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , 
     n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , 
     n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , 
     n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , 
     n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , 
     n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , 
     n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , 
     n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , 
     n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , 
     n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , 
     n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , 
     n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , 
     n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , 
     n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , 
     n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , 
     n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , 
     n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , 
     n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , 
     n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , 
     n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , 
     n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , 
     n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , 
     n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , 
     n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , 
     n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , 
     n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , 
     n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , 
     n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , 
     n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , 
     n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , 
     n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , 
     n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , 
     n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , 
     n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , 
     n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , 
     n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , 
     n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , 
     n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , 
     n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , 
     n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , 
     n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , 
     n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , 
     n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , 
     n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , 
     n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , 
     n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , 
     n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , 
     n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , 
     n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , 
     n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , 
     n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , 
     n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , 
     n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , 
     n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , 
     n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , 
     n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , 
     n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , 
     n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , 
     n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , 
     n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , 
     n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , 
     n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , 
     n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , 
     n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , 
     n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , 
     n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , 
     n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , 
     n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , 
     n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , 
     n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , 
     n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , 
     n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , 
     n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , 
     n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , 
     n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , 
     n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , 
     n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , 
     n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , 
     n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , 
     n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , 
     n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , 
     n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , 
     n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , 
     n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , 
     n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , 
     n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , 
     n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , 
     n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , 
     n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , 
     n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , 
     n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , 
     n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , 
     n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , 
     n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , 
     n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , 
     n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , 
     n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , 
     n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , 
     n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , 
     n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , 
     n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , 
     n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , 
     n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , 
     n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , 
     n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , 
     n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , 
     n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , 
     n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , 
     n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , 
     n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , 
     n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , 
     n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , 
     n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , 
     n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , 
     n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , 
     n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , 
     n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , 
     n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , 
     n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , 
     n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , 
     n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , 
     n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , 
     n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , 
     n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , 
     n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , 
     n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , 
     n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , 
     n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , 
     n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , 
     n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , 
     n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , 
     n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , 
     n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , 
     n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , 
     n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , 
     n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , 
     n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , 
     n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , 
     n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , 
     n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , 
     n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , 
     n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , 
     n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , 
     n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , 
     n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , 
     n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , 
     n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , 
     n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , 
     n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , 
     n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , 
     n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , 
     n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , 
     n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , 
     n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , 
     n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , 
     n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , 
     n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , 
     n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , 
     n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , 
     n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , 
     n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , 
     n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , 
     n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , 
     n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , 
     n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , 
     n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , 
     n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , 
     n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , 
     n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , 
     n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , 
     n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , 
     n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , 
     n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , 
     n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , 
     n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , 
     n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , 
     n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , 
     n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , 
     n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , 
     n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , 
     n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , 
     n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , 
     n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , 
     n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , 
     n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , 
     n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , 
     n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , 
     n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , 
     n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , 
     n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , 
     n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , 
     n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , 
     n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , 
     n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , 
     n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , 
     n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , 
     n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , 
     n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , 
     n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , 
     n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , 
     n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , 
     n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , 
     n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , 
     n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , 
     n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , 
     n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , 
     n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , 
     n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , 
     n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , 
     n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , 
     n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , 
     n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , 
     n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , 
     n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , 
     n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , 
     n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , 
     n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , 
     n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , 
     n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , 
     n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , 
     n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , 
     n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , 
     n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , 
     n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , 
     n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , 
     n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , 
     n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , 
     n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , 
     n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , 
     n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , 
     n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , 
     n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , 
     n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , 
     n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , 
     n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , 
     n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , 
     n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , 
     n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , 
     n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , 
     n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , 
     n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , 
     n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , 
     n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , 
     n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , 
     n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , 
     n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , 
     n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , 
     n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , 
     n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , 
     n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , 
     n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , 
     n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , 
     n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , 
     n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , 
     n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , 
     n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , 
     n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , 
     n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , 
     n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , 
     n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , 
     n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , 
     n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , 
     n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , 
     n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , 
     n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , 
     n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , 
     n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , 
     n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , 
     n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , 
     n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , 
     n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , 
     n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , 
     n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , 
     n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , 
     n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , 
     n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , 
     n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , 
     n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , 
     n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , 
     n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , 
     n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , 
     n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , 
     n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , 
     n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , 
     n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , 
     n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , 
     n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , 
     n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , 
     n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , 
     n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , 
     n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , 
     n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , 
     n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , 
     n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , 
     n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , 
     n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , 
     n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , 
     n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , 
     n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , 
     n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , 
     n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , 
     n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , 
     n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , 
     n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , 
     n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , 
     n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , 
     n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , 
     n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , 
     n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , 
     n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , 
     n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , 
     n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , 
     n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , 
     n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , 
     n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , 
     n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , 
     n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , 
     n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , 
     n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , 
     n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , 
     n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , 
     n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , 
     n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , 
     n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , 
     n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , 
     n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , 
     n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , 
     n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , 
     n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , 
     n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , 
     n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , 
     n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , 
     n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , 
     n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , 
     n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , 
     n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , 
     n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , 
     n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , 
     n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , 
     n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , 
     n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , 
     n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , 
     n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , 
     n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , 
     n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , 
     n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , 
     n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , 
     n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , 
     n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , 
     n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , 
     n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , 
     n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , 
     n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , 
     n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , 
     n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , 
     n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , 
     n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , 
     n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , 
     n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , 
     n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , 
     n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , 
     n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , 
     n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , 
     n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , 
     n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , 
     n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , 
     n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , 
     n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , 
     n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , 
     n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , 
     n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , 
     n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , 
     n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , 
     n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , 
     n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , 
     n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , 
     n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , 
     n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , 
     n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , 
     n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , 
     n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , 
     n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , 
     n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , 
     n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , 
     n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , 
     n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , 
     n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , 
     n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , 
     n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , 
     n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , 
     n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , 
     n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , 
     n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , 
     n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , 
     n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , 
     n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , 
     n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , 
     n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , 
     n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , 
     n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , 
     n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , 
     n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , 
     n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , 
     n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , 
     n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , 
     n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , 
     n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , 
     n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , 
     n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , 
     n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , 
     n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , 
     n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , 
     n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , 
     n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , 
     n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , 
     n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , 
     n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , 
     n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , 
     n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , 
     n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , 
     n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , 
     n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , 
     n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , 
     n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , 
     n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , 
     n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , 
     n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , 
     n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , 
     n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , 
     n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , 
     n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , 
     n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , 
     n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , 
     n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , 
     n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , 
     n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , 
     n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , 
     n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , 
     n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , 
     n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , 
     n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , 
     n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , 
     n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , 
     n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , 
     n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , 
     n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , 
     n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , 
     n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , 
     n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , 
     n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , 
     n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , 
     n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , 
     n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , 
     n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , 
     n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , 
     n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , 
     n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , 
     n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , 
     n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , 
     n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , 
     n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , 
     n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , 
     n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , 
     n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , 
     n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , 
     n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , 
     n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , 
     n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , 
     n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , 
     n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , 
     n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , 
     n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , 
     n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , 
     n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , 
     n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , 
     n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , 
     n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , 
     n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , 
     n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , 
     n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , 
     n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , 
     n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , 
     n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , 
     n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , 
     n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , 
     n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , 
     n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , 
     n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , 
     n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , 
     n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , 
     n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , 
     n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , 
     n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , 
     n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , 
     n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , 
     n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , 
     n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , 
     n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , 
     n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , 
     n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , 
     n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , 
     n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , 
     n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , 
     n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , 
     n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , 
     n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , 
     n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , 
     n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , 
     n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , 
     n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , 
     n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , 
     n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , 
     n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , 
     n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , 
     n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , 
     n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , 
     n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , 
     n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , 
     n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , 
     n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , 
     n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , 
     n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , 
     n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , 
     n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , 
     n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , 
     n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , 
     n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , 
     n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , 
     n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , 
     n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , 
     n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , 
     n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , 
     n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , 
     n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , 
     n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , 
     n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , 
     n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , 
     n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , 
     n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , 
     n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , 
     n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , 
     n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , 
     n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , 
     n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , 
     n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , 
     n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , 
     n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , 
     n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , 
     n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , 
     n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , 
     n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , 
     n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , 
     n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , 
     n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , 
     n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , 
     n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , 
     n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , 
     n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , 
     n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , 
     n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , 
     n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , 
     n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , 
     n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , 
     n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , 
     n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , 
     n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , 
     n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , 
     n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , 
     n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , 
     n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , 
     n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , 
     n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , 
     n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , 
     n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , 
     n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , 
     n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , 
     n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , 
     n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , 
     n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , 
     n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , 
     n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , 
     n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , 
     n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , 
     n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , 
     n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , 
     n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , 
     n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , 
     n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , 
     n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , 
     n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , 
     n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , 
     n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , 
     n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , 
     n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , 
     n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , 
     n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , 
     n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , 
     n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , 
     n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , 
     n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , 
     n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , 
     n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , 
     n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , 
     n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , 
     n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , 
     n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , 
     n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , 
     n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , 
     n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , 
     n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , 
     n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , 
     n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , 
     n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , 
     n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , 
     n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , 
     n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , 
     n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , 
     n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , 
     n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , 
     n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , 
     n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , 
     n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , 
     n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , 
     n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , 
     n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , 
     n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , 
     n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , 
     n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , 
     n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , 
     n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , 
     n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , 
     n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , 
     n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , 
     n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , 
     n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , 
     n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , 
     n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , 
     n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , 
     n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , 
     n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , 
     n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , 
     n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , 
     n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , 
     n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , 
     n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , 
     n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , 
     n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , 
     n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , 
     n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , 
     n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , 
     n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , 
     n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , 
     n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , 
     n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , 
     n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , 
     n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , 
     n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , 
     n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , 
     n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , 
     n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , 
     n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , 
     n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , 
     n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , 
     n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , 
     n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , 
     n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , 
     n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , 
     n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , 
     n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , 
     n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , 
     n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , 
     n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , 
     n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , 
     n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , 
     n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , 
     n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , 
     n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , 
     n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , 
     n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , 
     n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , 
     n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , 
     n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , 
     n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , 
     n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , 
     n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , 
     n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , 
     n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , 
     n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , 
     n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , 
     n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , 
     n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , 
     n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , 
     n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , 
     n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , 
     n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , 
     n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , 
     n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , 
     n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , 
     n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , 
     n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , 
     n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , 
     n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , 
     n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , 
     n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , 
     n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , 
     n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , 
     n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , 
     n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , 
     n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , 
     n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , 
     n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , 
     n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , 
     n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , 
     n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , 
     n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , 
     n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , 
     n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , 
     n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , 
     n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , 
     n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , 
     n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , 
     n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , 
     n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , 
     n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , 
     n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , 
     n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , 
     n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , 
     n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , 
     n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , 
     n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , 
     n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , 
     n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , 
     n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , 
     n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , 
     n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , 
     n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , 
     n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , 
     n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , 
     n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , 
     n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , 
     n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , 
     n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , 
     n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , 
     n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , 
     n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , 
     n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , 
     n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , 
     n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , 
     n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , 
     n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , 
     n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , 
     n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , 
     n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , 
     n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , 
     n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , 
     n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , 
     n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , 
     n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , 
     n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , 
     n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , 
     n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , 
     n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , 
     n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , 
     n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , 
     n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , 
     n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , 
     n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , 
     n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , 
     n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , 
     n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , 
     n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , 
     n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , 
     n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , 
     n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , 
     n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , 
     n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , 
     n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , 
     n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , 
     n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , 
     n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , 
     n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , 
     n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , 
     n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , 
     n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , 
     n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , 
     n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , 
     n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , 
     n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , 
     n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , 
     n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , 
     n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , 
     n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , 
     n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , 
     n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , 
     n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , 
     n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , 
     n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , 
     n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , 
     n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , 
     n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , 
     n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , 
     n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , 
     n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , 
     n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , 
     n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , 
     n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , 
     n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , 
     n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , 
     n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , 
     n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , 
     n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , 
     n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , 
     n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , 
     n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , 
     n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , 
     n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , 
     n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , 
     n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , 
     n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , 
     n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , 
     n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , 
     n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , 
     n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , 
     n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , 
     n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , 
     n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , 
     n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , 
     n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , 
     n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , 
     n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , 
     n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , 
     n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , 
     n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , 
     n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , 
     n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , 
     n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , 
     n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , 
     n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , 
     n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , 
     n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , 
     n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , 
     n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , 
     n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , 
     n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , 
     n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , 
     n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , 
     n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , 
     n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , 
     n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , 
     n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , 
     n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , 
     n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , 
     n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , 
     n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , 
     n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , 
     n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , 
     n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , 
     n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , 
     n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , 
     n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , 
     n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , 
     n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , 
     n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , 
     n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , 
     n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , 
     n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , 
     n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , 
     n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , 
     n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , 
     n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , 
     n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , 
     n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , 
     n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , 
     n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , 
     n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , 
     n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , 
     n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , 
     n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , 
     n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , 
     n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , 
     n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , 
     n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , 
     n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , 
     n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , 
     n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , 
     n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , 
     n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , 
     n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , 
     n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , 
     n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , 
     n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , 
     n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , 
     n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , 
     n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , 
     n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , 
     n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , 
     n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , 
     n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , 
     n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , 
     n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , 
     n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , 
     n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , 
     n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , 
     n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , 
     n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , 
     n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , 
     n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , 
     n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , 
     n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , 
     n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , 
     n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , 
     n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , 
     n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , 
     n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , 
     n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , 
     n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , 
     n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , 
     n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , 
     n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , 
     n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , 
     n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , 
     n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , 
     n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , 
     n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , 
     n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , 
     n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , 
     n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , 
     n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , 
     n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , 
     n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , 
     n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , 
     n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , 
     n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , 
     n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , 
     n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , 
     n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , 
     n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , 
     n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , 
     n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , 
     n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , 
     n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , 
     n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , 
     n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , 
     n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , 
     n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , 
     n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , 
     n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , 
     n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , 
     n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , 
     n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , 
     n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , 
     n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , 
     n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , 
     n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , 
     n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , 
     n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , 
     n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , 
     n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , 
     n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , 
     n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , 
     n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , 
     n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , 
     n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , 
     n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , 
     n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , 
     n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , 
     n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , 
     n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , 
     n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , 
     n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , 
     n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , 
     n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , 
     n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , 
     n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , 
     n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , 
     n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , 
     n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , 
     n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , 
     n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , 
     n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , 
     n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , 
     n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , 
     n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , 
     n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , 
     n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , 
     n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , 
     n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , 
     n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , 
     n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , 
     n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , 
     n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , 
     n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , 
     n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , 
     n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , 
     n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , 
     n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , 
     n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , 
     n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , 
     n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , 
     n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , 
     n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , 
     n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , 
     n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , 
     n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , 
     n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , 
     n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , 
     n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , 
     n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , 
     n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , 
     n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , 
     n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , 
     n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , 
     n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , 
     n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , 
     n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , 
     n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , 
     n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , 
     n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , 
     n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , 
     n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , 
     n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , 
     n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , 
     n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , 
     n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , 
     n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , 
     n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , 
     n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , 
     n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , 
     n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , 
     n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , 
     n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , 
     n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , 
     n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , 
     n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , 
     n28941 , n28942 , n28943 , n28944 , n28945 , n28946 ;
buf ( n2192 , n13764 );
buf ( n2187 , n15439 );
buf ( n2190 , n19023 );
buf ( n2191 , n22066 );
buf ( n2193 , n23533 );
buf ( n2188 , n25011 );
buf ( n2189 , n26202 );
buf ( n2194 , n27139 );
buf ( n2195 , n28210 );
buf ( n2186 , n28946 );
buf ( n4394 , n2081 );
buf ( n4395 , n1581 );
buf ( n4396 , n1572 );
buf ( n4397 , n1274 );
buf ( n4398 , n811 );
buf ( n4399 , n1423 );
buf ( n4400 , n1546 );
buf ( n4401 , n664 );
buf ( n4402 , n918 );
buf ( n4403 , n413 );
buf ( n4404 , n2133 );
buf ( n4405 , n201 );
buf ( n4406 , n434 );
buf ( n4407 , n317 );
buf ( n4408 , n2023 );
buf ( n4409 , n882 );
buf ( n4410 , n1634 );
buf ( n4411 , n888 );
buf ( n4412 , n1142 );
buf ( n4413 , n349 );
buf ( n4414 , n729 );
buf ( n4415 , n1315 );
buf ( n4416 , n189 );
buf ( n4417 , n2176 );
buf ( n4418 , n168 );
buf ( n4419 , n164 );
buf ( n4420 , n831 );
buf ( n4421 , n979 );
buf ( n4422 , n1841 );
buf ( n4423 , n1855 );
buf ( n4424 , n1690 );
buf ( n4425 , n261 );
buf ( n4426 , n1901 );
buf ( n4427 , n1822 );
buf ( n4428 , n660 );
buf ( n4429 , n669 );
buf ( n4430 , n1715 );
buf ( n4431 , n684 );
buf ( n4432 , n2119 );
buf ( n4433 , n513 );
buf ( n4434 , n1828 );
buf ( n4435 , n4 );
buf ( n4436 , n716 );
buf ( n4437 , n1020 );
buf ( n4438 , n835 );
buf ( n4439 , n105 );
buf ( n4440 , n1615 );
buf ( n4441 , n397 );
buf ( n4442 , n1273 );
buf ( n4443 , n1550 );
buf ( n4444 , n1132 );
buf ( n4445 , n1804 );
buf ( n4446 , n1413 );
buf ( n4447 , n17 );
buf ( n4448 , n57 );
buf ( n4449 , n1023 );
buf ( n4450 , n1704 );
buf ( n4451 , n2039 );
buf ( n4452 , n120 );
buf ( n4453 , n1533 );
buf ( n4454 , n1650 );
buf ( n4455 , n1697 );
buf ( n4456 , n1563 );
buf ( n4457 , n984 );
buf ( n4458 , n2005 );
buf ( n4459 , n1552 );
buf ( n4460 , n1063 );
buf ( n4461 , n410 );
buf ( n4462 , n1995 );
buf ( n4463 , n1880 );
buf ( n4464 , n1117 );
buf ( n4465 , n1340 );
buf ( n4466 , n1971 );
buf ( n4467 , n1104 );
buf ( n4468 , n335 );
buf ( n4469 , n297 );
buf ( n4470 , n455 );
buf ( n4471 , n2018 );
buf ( n4472 , n804 );
buf ( n4473 , n374 );
buf ( n4474 , n0 );
buf ( n4475 , n1979 );
buf ( n4476 , n1625 );
buf ( n4477 , n296 );
buf ( n4478 , n304 );
buf ( n4479 , n1862 );
buf ( n4480 , n622 );
buf ( n4481 , n863 );
buf ( n4482 , n302 );
buf ( n4483 , n648 );
buf ( n4484 , n1433 );
buf ( n4485 , n850 );
buf ( n4486 , n80 );
buf ( n4487 , n1173 );
buf ( n4488 , n920 );
buf ( n4489 , n1022 );
buf ( n4490 , n584 );
buf ( n4491 , n173 );
buf ( n4492 , n219 );
buf ( n4493 , n1418 );
buf ( n4494 , n824 );
buf ( n4495 , n309 );
buf ( n4496 , n2076 );
buf ( n4497 , n659 );
buf ( n4498 , n2108 );
buf ( n4499 , n1842 );
buf ( n4500 , n1761 );
buf ( n4501 , n352 );
buf ( n4502 , n502 );
buf ( n4503 , n868 );
buf ( n4504 , n807 );
buf ( n4505 , n1976 );
buf ( n4506 , n631 );
buf ( n4507 , n332 );
buf ( n4508 , n1099 );
buf ( n4509 , n1577 );
buf ( n4510 , n2159 );
buf ( n4511 , n283 );
buf ( n4512 , n405 );
buf ( n4513 , n1989 );
buf ( n4514 , n1345 );
buf ( n4515 , n624 );
buf ( n4516 , n86 );
buf ( n4517 , n399 );
buf ( n4518 , n110 );
buf ( n4519 , n485 );
buf ( n4520 , n152 );
buf ( n4521 , n1566 );
buf ( n4522 , n1896 );
buf ( n4523 , n1900 );
buf ( n4524 , n954 );
buf ( n4525 , n518 );
buf ( n4526 , n1522 );
buf ( n4527 , n72 );
buf ( n4528 , n2153 );
buf ( n4529 , n114 );
buf ( n4530 , n1276 );
buf ( n4531 , n69 );
buf ( n4532 , n7 );
buf ( n4533 , n986 );
buf ( n4534 , n2096 );
buf ( n4535 , n890 );
buf ( n4536 , n1564 );
buf ( n4537 , n2052 );
buf ( n4538 , n74 );
buf ( n4539 , n1961 );
buf ( n4540 , n833 );
buf ( n4541 , n1261 );
buf ( n4542 , n2134 );
buf ( n4543 , n123 );
buf ( n4544 , n1654 );
buf ( n4545 , n849 );
buf ( n4546 , n1923 );
buf ( n4547 , n1348 );
buf ( n4548 , n151 );
buf ( n4549 , n1560 );
buf ( n4550 , n1685 );
buf ( n4551 , n577 );
buf ( n4552 , n969 );
buf ( n4553 , n1120 );
buf ( n4554 , n310 );
buf ( n4555 , n1435 );
buf ( n4556 , n77 );
buf ( n4557 , n533 );
buf ( n4558 , n761 );
buf ( n4559 , n1832 );
buf ( n4560 , n841 );
buf ( n4561 , n1228 );
buf ( n4562 , n504 );
buf ( n4563 , n756 );
buf ( n4564 , n2008 );
buf ( n4565 , n1622 );
buf ( n4566 , n205 );
buf ( n4567 , n864 );
buf ( n4568 , n1873 );
buf ( n4569 , n2012 );
buf ( n4570 , n1155 );
buf ( n4571 , n2014 );
buf ( n4572 , n323 );
buf ( n4573 , n337 );
buf ( n4574 , n842 );
buf ( n4575 , n598 );
buf ( n4576 , n1882 );
buf ( n4577 , n1585 );
buf ( n4578 , n486 );
buf ( n4579 , n388 );
buf ( n4580 , n1736 );
buf ( n4581 , n609 );
buf ( n4582 , n326 );
buf ( n4583 , n732 );
buf ( n4584 , n1477 );
buf ( n4585 , n12 );
buf ( n4586 , n357 );
buf ( n4587 , n1212 );
buf ( n4588 , n303 );
buf ( n4589 , n1876 );
buf ( n4590 , n776 );
buf ( n4591 , n1929 );
buf ( n4592 , n1919 );
buf ( n4593 , n401 );
buf ( n4594 , n953 );
buf ( n4595 , n1005 );
buf ( n4596 , n76 );
buf ( n4597 , n1946 );
buf ( n4598 , n412 );
buf ( n4599 , n55 );
buf ( n4600 , n1075 );
buf ( n4601 , n217 );
buf ( n4602 , n774 );
buf ( n4603 , n654 );
buf ( n4604 , n696 );
buf ( n4605 , n53 );
buf ( n4606 , n1883 );
buf ( n4607 , n1555 );
buf ( n4608 , n1621 );
buf ( n4609 , n1865 );
buf ( n4610 , n697 );
buf ( n4611 , n1283 );
buf ( n4612 , n1260 );
buf ( n4613 , n977 );
buf ( n4614 , n1993 );
buf ( n4615 , n725 );
buf ( n4616 , n163 );
buf ( n4617 , n741 );
buf ( n4618 , n1270 );
buf ( n4619 , n1877 );
buf ( n4620 , n1436 );
buf ( n4621 , n1514 );
buf ( n4622 , n1368 );
buf ( n4623 , n231 );
buf ( n4624 , n1707 );
buf ( n4625 , n524 );
buf ( n4626 , n1465 );
buf ( n4627 , n5 );
buf ( n4628 , n213 );
buf ( n4629 , n318 );
buf ( n4630 , n1352 );
buf ( n4631 , n2028 );
buf ( n4632 , n1308 );
buf ( n4633 , n921 );
buf ( n4634 , n508 );
buf ( n4635 , n320 );
buf ( n4636 , n243 );
buf ( n4637 , n22 );
buf ( n4638 , n793 );
buf ( n4639 , n1740 );
buf ( n4640 , n2055 );
buf ( n4641 , n1596 );
buf ( n4642 , n32 );
buf ( n4643 , n245 );
buf ( n4644 , n1028 );
buf ( n4645 , n992 );
buf ( n4646 , n1443 );
buf ( n4647 , n1358 );
buf ( n4648 , n149 );
buf ( n4649 , n1905 );
buf ( n4650 , n376 );
buf ( n4651 , n948 );
buf ( n4652 , n325 );
buf ( n4653 , n394 );
buf ( n4654 , n1893 );
buf ( n4655 , n468 );
buf ( n4656 , n1638 );
buf ( n4657 , n2074 );
buf ( n4658 , n1933 );
buf ( n4659 , n1516 );
buf ( n4660 , n364 );
buf ( n4661 , n1030 );
buf ( n4662 , n1609 );
buf ( n4663 , n340 );
buf ( n4664 , n246 );
buf ( n4665 , n2152 );
buf ( n4666 , n990 );
buf ( n4667 , n1363 );
buf ( n4668 , n663 );
buf ( n4669 , n652 );
buf ( n4670 , n2184 );
buf ( n4671 , n299 );
buf ( n4672 , n249 );
buf ( n4673 , n1612 );
buf ( n4674 , n1027 );
buf ( n4675 , n1366 );
buf ( n4676 , n235 );
buf ( n4677 , n2060 );
buf ( n4678 , n665 );
buf ( n4679 , n829 );
buf ( n4680 , n547 );
buf ( n4681 , n1911 );
buf ( n4682 , n955 );
buf ( n4683 , n1057 );
buf ( n4684 , n1805 );
buf ( n4685 , n1395 );
buf ( n4686 , n880 );
buf ( n4687 , n2021 );
buf ( n4688 , n579 );
buf ( n4689 , n1486 );
buf ( n4690 , n2162 );
buf ( n4691 , n1990 );
buf ( n4692 , n871 );
buf ( n4693 , n1932 );
buf ( n4694 , n505 );
buf ( n4695 , n2047 );
buf ( n4696 , n146 );
buf ( n4697 , n1216 );
buf ( n4698 , n1288 );
buf ( n4699 , n2066 );
buf ( n4700 , n1249 );
buf ( n4701 , n1518 );
buf ( n4702 , n2017 );
buf ( n4703 , n571 );
buf ( n4704 , n724 );
buf ( n4705 , n884 );
buf ( n4706 , n1215 );
buf ( n4707 , n1986 );
buf ( n4708 , n1046 );
buf ( n4709 , n1602 );
buf ( n4710 , n737 );
buf ( n4711 , n1498 );
buf ( n4712 , n98 );
buf ( n4713 , n1399 );
buf ( n4714 , n26 );
buf ( n4715 , n452 );
buf ( n4716 , n1408 );
buf ( n4717 , n1909 );
buf ( n4718 , n1233 );
buf ( n4719 , n1412 );
buf ( n4720 , n132 );
buf ( n4721 , n1000 );
buf ( n4722 , n530 );
buf ( n4723 , n1767 );
buf ( n4724 , n1515 );
buf ( n4725 , n1067 );
buf ( n4726 , n328 );
buf ( n4727 , n887 );
buf ( n4728 , n457 );
buf ( n4729 , n1992 );
buf ( n4730 , n1951 );
buf ( n4731 , n371 );
buf ( n4732 , n338 );
buf ( n4733 , n840 );
buf ( n4734 , n2138 );
buf ( n4735 , n933 );
buf ( n4736 , n1401 );
buf ( n4737 , n2129 );
buf ( n4738 , n1520 );
buf ( n4739 , n2168 );
buf ( n4740 , n260 );
buf ( n4741 , n18 );
buf ( n4742 , n1617 );
buf ( n4743 , n1907 );
buf ( n4744 , n1603 );
buf ( n4745 , n2090 );
buf ( n4746 , n1481 );
buf ( n4747 , n1508 );
buf ( n4748 , n594 );
buf ( n4749 , n2183 );
buf ( n4750 , n1610 );
buf ( n4751 , n1679 );
buf ( n4752 , n599 );
buf ( n4753 , n1079 );
buf ( n4754 , n589 );
buf ( n4755 , n830 );
buf ( n4756 , n95 );
buf ( n4757 , n140 );
buf ( n4758 , n568 );
buf ( n4759 , n1879 );
buf ( n4760 , n587 );
buf ( n4761 , n2013 );
buf ( n4762 , n674 );
buf ( n4763 , n788 );
buf ( n4764 , n1264 );
buf ( n4765 , n1683 );
buf ( n4766 , n723 );
buf ( n4767 , n2070 );
buf ( n4768 , n785 );
buf ( n4769 , n1831 );
buf ( n4770 , n2000 );
buf ( n4771 , n135 );
buf ( n4772 , n1637 );
buf ( n4773 , n33 );
buf ( n4774 , n1525 );
buf ( n4775 , n158 );
buf ( n4776 , n1013 );
buf ( n4777 , n2099 );
buf ( n4778 , n1776 );
buf ( n4779 , n2175 );
buf ( n4780 , n1833 );
buf ( n4781 , n828 );
buf ( n4782 , n744 );
buf ( n4783 , n1298 );
buf ( n4784 , n2125 );
buf ( n4785 , n653 );
buf ( n4786 , n1968 );
buf ( n4787 , n503 );
buf ( n4788 , n1984 );
buf ( n4789 , n1047 );
buf ( n4790 , n1431 );
buf ( n4791 , n2082 );
buf ( n4792 , n772 );
buf ( n4793 , n813 );
buf ( n4794 , n1152 );
buf ( n4795 , n982 );
buf ( n4796 , n1997 );
buf ( n4797 , n1278 );
buf ( n4798 , n1179 );
buf ( n4799 , n1280 );
buf ( n4800 , n211 );
buf ( n4801 , n386 );
buf ( n4802 , n1269 );
buf ( n4803 , n254 );
buf ( n4804 , n1620 );
buf ( n4805 , n2149 );
buf ( n4806 , n826 );
buf ( n4807 , n854 );
buf ( n4808 , n759 );
buf ( n4809 , n1664 );
buf ( n4810 , n980 );
buf ( n4811 , n543 );
buf ( n4812 , n119 );
buf ( n4813 , n2095 );
buf ( n4814 , n934 );
buf ( n4815 , n188 );
buf ( n4816 , n927 );
buf ( n4817 , n495 );
buf ( n4818 , n435 );
buf ( n4819 , n630 );
buf ( n4820 , n1076 );
buf ( n4821 , n75 );
buf ( n4822 , n1207 );
buf ( n4823 , n658 );
buf ( n4824 , n1912 );
buf ( n4825 , n1749 );
buf ( n4826 , n1648 );
buf ( n4827 , n1497 );
buf ( n4828 , n974 );
buf ( n4829 , n1474 );
buf ( n4830 , n1641 );
buf ( n4831 , n1836 );
buf ( n4832 , n102 );
buf ( n4833 , n1802 );
buf ( n4834 , n731 );
buf ( n4835 , n606 );
buf ( n4836 , n150 );
buf ( n4837 , n1999 );
buf ( n4838 , n1245 );
buf ( n4839 , n509 );
buf ( n4840 , n1405 );
buf ( n4841 , n2139 );
buf ( n4842 , n1972 );
buf ( n4843 , n1604 );
buf ( n4844 , n2062 );
buf ( n4845 , n1529 );
buf ( n4846 , n1854 );
buf ( n4847 , n1209 );
buf ( n4848 , n1386 );
buf ( n4849 , n629 );
buf ( n4850 , n1981 );
buf ( n4851 , n1895 );
buf ( n4852 , n592 );
buf ( n4853 , n672 );
buf ( n4854 , n1045 );
buf ( n4855 , n1591 );
buf ( n4856 , n1955 );
buf ( n4857 , n363 );
buf ( n4858 , n1821 );
buf ( n4859 , n1387 );
buf ( n4860 , n298 );
buf ( n4861 , n1226 );
buf ( n4862 , n968 );
buf ( n4863 , n1452 );
buf ( n4864 , n91 );
buf ( n4865 , n492 );
buf ( n4866 , n1456 );
buf ( n4867 , n2004 );
buf ( n4868 , n699 );
buf ( n4869 , n626 );
buf ( n4870 , n789 );
buf ( n4871 , n1475 );
buf ( n4872 , n1642 );
buf ( n4873 , n1784 );
buf ( n4874 , n329 );
buf ( n4875 , n705 );
buf ( n4876 , n681 );
buf ( n4877 , n962 );
buf ( n4878 , n1191 );
buf ( n4879 , n268 );
buf ( n4880 , n9 );
buf ( n4881 , n2078 );
buf ( n4882 , n604 );
buf ( n4883 , n1427 );
buf ( n4884 , n1250 );
buf ( n4885 , n65 );
buf ( n4886 , n2177 );
buf ( n4887 , n1942 );
buf ( n4888 , n1379 );
buf ( n4889 , n666 );
buf ( n4890 , n2140 );
buf ( n4891 , n964 );
buf ( n4892 , n290 );
buf ( n4893 , n700 );
buf ( n4894 , n1314 );
buf ( n4895 , n1128 );
buf ( n4896 , n676 );
buf ( n4897 , n1820 );
buf ( n4898 , n633 );
buf ( n4899 , n575 );
buf ( n4900 , n1187 );
buf ( n4901 , n1248 );
buf ( n4902 , n1917 );
buf ( n4903 , n469 );
buf ( n4904 , n1328 );
buf ( n4905 , n541 );
buf ( n4906 , n1597 );
buf ( n4907 , n1960 );
buf ( n4908 , n645 );
buf ( n4909 , n407 );
buf ( n4910 , n430 );
buf ( n4911 , n966 );
buf ( n4912 , n2169 );
buf ( n4913 , n1246 );
buf ( n4914 , n701 );
buf ( n4915 , n1757 );
buf ( n4916 , n855 );
buf ( n4917 , n1201 );
buf ( n4918 , n1019 );
buf ( n4919 , n1496 );
buf ( n4920 , n1175 );
buf ( n4921 , n1014 );
buf ( n4922 , n1561 );
buf ( n4923 , n601 );
buf ( n4924 , n448 );
buf ( n4925 , n368 );
buf ( n4926 , n1015 );
buf ( n4927 , n1744 );
buf ( n4928 , n898 );
buf ( n4929 , n2093 );
buf ( n4930 , n514 );
buf ( n4931 , n360 );
buf ( n4932 , n1220 );
buf ( n4933 , n1869 );
buf ( n4934 , n190 );
buf ( n4935 , n1872 );
buf ( n4936 , n1827 );
buf ( n4937 , n1674 );
buf ( n4938 , n221 );
buf ( n4939 , n770 );
buf ( n4940 , n1826 );
buf ( n4941 , n2043 );
buf ( n4942 , n1780 );
buf ( n4943 , n753 );
buf ( n4944 , n1904 );
buf ( n4945 , n1655 );
buf ( n4946 , n1502 );
buf ( n4947 , n1823 );
buf ( n4948 , n1819 );
buf ( n4949 , n816 );
buf ( n4950 , n616 );
buf ( n4951 , n902 );
buf ( n4952 , n825 );
buf ( n4953 , n1086 );
buf ( n4954 , n2006 );
buf ( n4955 , n1171 );
buf ( n4956 , n441 );
buf ( n4957 , n1967 );
buf ( n4958 , n29 );
buf ( n4959 , n195 );
buf ( n4960 , n1480 );
buf ( n4961 , n212 );
buf ( n4962 , n236 );
buf ( n4963 , n1705 );
buf ( n4964 , n1186 );
buf ( n4965 , n1102 );
buf ( n4966 , n1962 );
buf ( n4967 , n550 );
buf ( n4968 , n248 );
buf ( n4969 , n286 );
buf ( n4970 , n1856 );
buf ( n4971 , n1599 );
buf ( n4972 , n2077 );
buf ( n4973 , n628 );
buf ( n4974 , n935 );
buf ( n4975 , n963 );
buf ( n4976 , n160 );
buf ( n4977 , n1899 );
buf ( n4978 , n2020 );
buf ( n4979 , n768 );
buf ( n4980 , n1991 );
buf ( n4981 , n1208 );
buf ( n4982 , n2071 );
buf ( n4983 , n499 );
buf ( n4984 , n15 );
buf ( n4985 , n1772 );
buf ( n4986 , n1943 );
buf ( n4987 , n852 );
buf ( n4988 , n1875 );
buf ( n4989 , n817 );
buf ( n4990 , n71 );
buf ( n4991 , n557 );
buf ( n4992 , n1732 );
buf ( n4993 , n2024 );
buf ( n4994 , n50 );
buf ( n4995 , n1948 );
buf ( n4996 , n1853 );
buf ( n4997 , n1285 );
buf ( n4998 , n688 );
buf ( n4999 , n1157 );
buf ( n5000 , n1567 );
buf ( n5001 , n634 );
buf ( n5002 , n1162 );
buf ( n5003 , n178 );
buf ( n5004 , n536 );
buf ( n5005 , n906 );
buf ( n5006 , n1039 );
buf ( n5007 , n951 );
buf ( n5008 , n1380 );
buf ( n5009 , n1501 );
buf ( n5010 , n1381 );
buf ( n5011 , n108 );
buf ( n5012 , n746 );
buf ( n5013 , n2118 );
buf ( n5014 , n1537 );
buf ( n5015 , n432 );
buf ( n5016 , n2059 );
buf ( n5017 , n937 );
buf ( n5018 , n347 );
buf ( n5019 , n1606 );
buf ( n5020 , n501 );
buf ( n5021 , n1672 );
buf ( n5022 , n1031 );
buf ( n5023 , n88 );
buf ( n5024 , n1859 );
buf ( n5025 , n965 );
buf ( n5026 , n1286 );
buf ( n5027 , n300 );
buf ( n5028 , n1090 );
buf ( n5029 , n949 );
buf ( n5030 , n1794 );
buf ( n5031 , n1439 );
buf ( n5032 , n2073 );
buf ( n5033 , n563 );
buf ( n5034 , n2115 );
buf ( n5035 , n1354 );
buf ( n5036 , n1791 );
buf ( n5037 , n1367 );
buf ( n5038 , n30 );
buf ( n5039 , n784 );
buf ( n5040 , n815 );
buf ( n5041 , n943 );
buf ( n5042 , n1448 );
buf ( n5043 , n461 );
buf ( n5044 , n794 );
buf ( n5045 , n1032 );
buf ( n5046 , n554 );
buf ( n5047 , n2064 );
buf ( n5048 , n1463 );
buf ( n5049 , n20 );
buf ( n5050 , n1341 );
buf ( n5051 , n348 );
buf ( n5052 , n1969 );
buf ( n5053 , n295 );
buf ( n5054 , n1965 );
buf ( n5055 , n1107 );
buf ( n5056 , n433 );
buf ( n5057 , n316 );
buf ( n5058 , n1316 );
buf ( n5059 , n561 );
buf ( n5060 , n1973 );
buf ( n5061 , n1292 );
buf ( n5062 , n498 );
buf ( n5063 , n301 );
buf ( n5064 , n460 );
buf ( n5065 , n500 );
buf ( n5066 , n444 );
buf ( n5067 , n58 );
buf ( n5068 , n143 );
buf ( n5069 , n428 );
buf ( n5070 , n893 );
buf ( n5071 , n82 );
buf ( n5072 , n449 );
buf ( n5073 , n1103 );
buf ( n5074 , n714 );
buf ( n5075 , n641 );
buf ( n5076 , n379 );
buf ( n5077 , n1491 );
buf ( n5078 , n1489 );
buf ( n5079 , n1825 );
buf ( n5080 , n1816 );
buf ( n5081 , n709 );
buf ( n5082 , n42 );
buf ( n5083 , n754 );
buf ( n5084 , n782 );
buf ( n5085 , n981 );
buf ( n5086 , n1198 );
buf ( n5087 , n226 );
buf ( n5088 , n595 );
buf ( n5089 , n284 );
buf ( n5090 , n1695 );
buf ( n5091 , n2051 );
buf ( n5092 , n944 );
buf ( n5093 , n1614 );
buf ( n5094 , n1160 );
buf ( n5095 , n1845 );
buf ( n5096 , n230 );
buf ( n5097 , n764 );
buf ( n5098 , n156 );
buf ( n5099 , n800 );
buf ( n5100 , n956 );
buf ( n5101 , n2075 );
buf ( n5102 , n472 );
buf ( n5103 , n2136 );
buf ( n5104 , n1631 );
buf ( n5105 , n1575 );
buf ( n5106 , n978 );
buf ( n5107 , n1579 );
buf ( n5108 , n1582 );
buf ( n5109 , n1410 );
buf ( n5110 , n484 );
buf ( n5111 , n278 );
buf ( n5112 , n1526 );
buf ( n5113 , n1636 );
buf ( n5114 , n1289 );
buf ( n5115 , n1926 );
buf ( n5116 , n1726 );
buf ( n5117 , n172 );
buf ( n5118 , n1665 );
buf ( n5119 , n266 );
buf ( n5120 , n1196 );
buf ( n5121 , n895 );
buf ( n5122 , n605 );
buf ( n5123 , n1663 );
buf ( n5124 , n610 );
buf ( n5125 , n398 );
buf ( n5126 , n220 );
buf ( n5127 , n958 );
buf ( n5128 , n137 );
buf ( n5129 , n881 );
buf ( n5130 , n889 );
buf ( n5131 , n1257 );
buf ( n5132 , n113 );
buf ( n5133 , n851 );
buf ( n5134 , n1524 );
buf ( n5135 , n999 );
buf ( n5136 , n61 );
buf ( n5137 , n1008 );
buf ( n5138 , n1759 );
buf ( n5139 , n1910 );
buf ( n5140 , n569 );
buf ( n5141 , n67 );
buf ( n5142 , n345 );
buf ( n5143 , n834 );
buf ( n5144 , n856 );
buf ( n5145 , n1817 );
buf ( n5146 , n1043 );
buf ( n5147 , n1370 );
buf ( n5148 , n240 );
buf ( n5149 , n930 );
buf ( n5150 , n1513 );
buf ( n5151 , n1885 );
buf ( n5152 , n1239 );
buf ( n5153 , n19 );
buf ( n5154 , n2067 );
buf ( n5155 , n1768 );
buf ( n5156 , n2042 );
buf ( n5157 , n1710 );
buf ( n5158 , n564 );
buf ( n5159 , n623 );
buf ( n5160 , n1469 );
buf ( n5161 , n1098 );
buf ( n5162 , n845 );
buf ( n5163 , n1130 );
buf ( n5164 , n1199 );
buf ( n5165 , n1584 );
buf ( n5166 , n293 );
buf ( n5167 , n253 );
buf ( n5168 , n1483 );
buf ( n5169 , n265 );
buf ( n5170 , n1908 );
buf ( n5171 , n1139 );
buf ( n5172 , n973 );
buf ( n5173 , n1077 );
buf ( n5174 , n1108 );
buf ( n5175 , n1009 );
buf ( n5176 , n1897 );
buf ( n5177 , n130 );
buf ( n5178 , n1750 );
buf ( n5179 , n1952 );
buf ( n5180 , n755 );
buf ( n5181 , n1059 );
buf ( n5182 , n1033 );
buf ( n5183 , n972 );
buf ( n5184 , n2174 );
buf ( n5185 , n1072 );
buf ( n5186 , n506 );
buf ( n5187 , n988 );
buf ( n5188 , n1070 );
buf ( n5189 , n751 );
buf ( n5190 , n528 );
buf ( n5191 , n1742 );
buf ( n5192 , n493 );
buf ( n5193 , n1134 );
buf ( n5194 , n608 );
buf ( n5195 , n2097 );
buf ( n5196 , n531 );
buf ( n5197 , n1123 );
buf ( n5198 , n2178 );
buf ( n5199 , n689 );
buf ( n5200 , n1864 );
buf ( n5201 , n1332 );
buf ( n5202 , n2056 );
buf ( n5203 , n1263 );
buf ( n5204 , n2083 );
buf ( n5205 , n1738 );
buf ( n5206 , n1416 );
buf ( n5207 , n87 );
buf ( n5208 , n1361 );
buf ( n5209 , n415 );
buf ( n5210 , n101 );
buf ( n5211 , n1321 );
buf ( n5212 , n1646 );
buf ( n5213 , n928 );
buf ( n5214 , n1921 );
buf ( n5215 , n2101 );
buf ( n5216 , n1578 );
buf ( n5217 , n704 );
buf ( n5218 , n778 );
buf ( n5219 , n184 );
buf ( n5220 , n1766 );
buf ( n5221 , n1994 );
buf ( n5222 , n1562 );
buf ( n5223 , n1906 );
buf ( n5224 , n1195 );
buf ( n5225 , n1217 );
buf ( n5226 , n1868 );
buf ( n5227 , n1049 );
buf ( n5228 , n878 );
buf ( n5229 , n1781 );
buf ( n5230 , n1116 );
buf ( n5231 , n305 );
buf ( n5232 , n343 );
buf ( n5233 , n1225 );
buf ( n5234 , n2041 );
buf ( n5235 , n2167 );
buf ( n5236 , n996 );
buf ( n5237 , n703 );
buf ( n5238 , n1213 );
buf ( n5239 , n277 );
buf ( n5240 , n1396 );
buf ( n5241 , n2179 );
buf ( n5242 , n1093 );
buf ( n5243 , n1197 );
buf ( n5244 , n192 );
buf ( n5245 , n270 );
buf ( n5246 , n1016 );
buf ( n5247 , n1607 );
buf ( n5248 , n590 );
buf ( n5249 , n389 );
buf ( n5250 , n1141 );
buf ( n5251 , n210 );
buf ( n5252 , n1623 );
buf ( n5253 , n1957 );
buf ( n5254 , n511 );
buf ( n5255 , n2130 );
buf ( n5256 , n1126 );
buf ( n5257 , n1645 );
buf ( n5258 , n1056 );
buf ( n5259 , n186 );
buf ( n5260 , n1748 );
buf ( n5261 , n812 );
buf ( n5262 , n1037 );
buf ( n5263 , n593 );
buf ( n5264 , n239 );
buf ( n5265 , n447 );
buf ( n5266 , n607 );
buf ( n5267 , n177 );
buf ( n5268 , n549 );
buf ( n5269 , n1717 );
buf ( n5270 , n313 );
buf ( n5271 , n1505 );
buf ( n5272 , n2146 );
buf ( n5273 , n1454 );
buf ( n5274 , n1884 );
buf ( n5275 , n667 );
buf ( n5276 , n534 );
buf ( n5277 , n142 );
buf ( n5278 , n382 );
buf ( n5279 , n1041 );
buf ( n5280 , n1632 );
buf ( n5281 , n1982 );
buf ( n5282 , n581 );
buf ( n5283 , n707 );
buf ( n5284 , n1656 );
buf ( n5285 , n2166 );
buf ( n5286 , n1343 );
buf ( n5287 , n1756 );
buf ( n5288 , n848 );
buf ( n5289 , n946 );
buf ( n5290 , n1538 );
buf ( n5291 , n1357 );
buf ( n5292 , n762 );
buf ( n5293 , n344 );
buf ( n5294 , n2058 );
buf ( n5295 , n1402 );
buf ( n5296 , n367 );
buf ( n5297 , n1588 );
buf ( n5298 , n1806 );
buf ( n5299 , n68 );
buf ( n5300 , n1810 );
buf ( n5301 , n532 );
buf ( n5302 , n721 );
buf ( n5303 , n642 );
buf ( n5304 , n411 );
buf ( n5305 , n1970 );
buf ( n5306 , n1193 );
buf ( n5307 , n93 );
buf ( n5308 , n1587 );
buf ( n5309 , n92 );
buf ( n5310 , n60 );
buf ( n5311 , n1445 );
buf ( n5312 , n289 );
buf ( n5313 , n155 );
buf ( n5314 , n803 );
buf ( n5315 , n1846 );
buf ( n5316 , n2105 );
buf ( n5317 , n429 );
buf ( n5318 , n478 );
buf ( n5319 , n526 );
buf ( n5320 , n263 );
buf ( n5321 , n1799 );
buf ( n5322 , n2025 );
buf ( n5323 , n952 );
buf ( n5324 , n1662 );
buf ( n5325 , n154 );
buf ( n5326 , n994 );
buf ( n5327 , n1432 );
buf ( n5328 , n1192 );
buf ( n5329 , n169 );
buf ( n5330 , n420 );
buf ( n5331 , n1026 );
buf ( n5332 , n1773 );
buf ( n5333 , n2015 );
buf ( n5334 , n765 );
buf ( n5335 , n757 );
buf ( n5336 , n214 );
buf ( n5337 , n341 );
buf ( n5338 , n1383 );
buf ( n5339 , n822 );
buf ( n5340 , n1040 );
buf ( n5341 , n1692 );
buf ( n5342 , n1793 );
buf ( n5343 , n1282 );
buf ( n5344 , n378 );
buf ( n5345 , n1807 );
buf ( n5346 , n2009 );
buf ( n5347 , n913 );
buf ( n5348 , n40 );
buf ( n5349 , n1210 );
buf ( n5350 , n1788 );
buf ( n5351 , n1953 );
buf ( n5352 , n442 );
buf ( n5353 , n914 );
buf ( n5354 , n1360 );
buf ( n5355 , n1898 );
buf ( n5356 , n1291 );
buf ( n5357 , n867 );
buf ( n5358 , n1699 );
buf ( n5359 , n436 );
buf ( n5360 , n1012 );
buf ( n5361 , n1034 );
buf ( n5362 , n691 );
buf ( n5363 , n733 );
buf ( n5364 , n423 );
buf ( n5365 , n234 );
buf ( n5366 , n1156 );
buf ( n5367 , n1188 );
buf ( n5368 , n1741 );
buf ( n5369 , n1874 );
buf ( n5370 , n1221 );
buf ( n5371 , n462 );
buf ( n5372 , n170 );
buf ( n5373 , n148 );
buf ( n5374 , n1442 );
buf ( n5375 , n670 );
buf ( n5376 , n1222 );
buf ( n5377 , n677 );
buf ( n5378 , n1421 );
buf ( n5379 , n1643 );
buf ( n5380 , n1149 );
buf ( n5381 , n1301 );
buf ( n5382 , n819 );
buf ( n5383 , n1440 );
buf ( n5384 , n1441 );
buf ( n5385 , n2007 );
buf ( n5386 , n1004 );
buf ( n5387 , n1558 );
buf ( n5388 , n1327 );
buf ( n5389 , n256 );
buf ( n5390 , n1887 );
buf ( n5391 , n479 );
buf ( n5392 , n1534 );
buf ( n5393 , n175 );
buf ( n5394 , n1818 );
buf ( n5395 , n2092 );
buf ( n5396 , n51 );
buf ( n5397 , n161 );
buf ( n5398 , n1119 );
buf ( n5399 , n1472 );
buf ( n5400 , n1922 );
buf ( n5401 , n339 );
buf ( n5402 , n229 );
buf ( n5403 , n414 );
buf ( n5404 , n1111 );
buf ( n5405 , n1809 );
buf ( n5406 , n287 );
buf ( n5407 , n1290 );
buf ( n5408 , n1085 );
buf ( n5409 , n2151 );
buf ( n5410 , n385 );
buf ( n5411 , n720 );
buf ( n5412 , n1499 );
buf ( n5413 , n1996 );
buf ( n5414 , n2116 );
buf ( n5415 , n1131 );
buf ( n5416 , n116 );
buf ( n5417 , n615 );
buf ( n5418 , n621 );
buf ( n5419 , n191 );
buf ( n5420 , n1745 );
buf ( n5421 , n85 );
buf ( n5422 , n1493 );
buf ( n5423 , n1153 );
buf ( n5424 , n873 );
buf ( n5425 , n1109 );
buf ( n5426 , n827 );
buf ( n5427 , n1415 );
buf ( n5428 , n939 );
buf ( n5429 , n1696 );
buf ( n5430 , n2180 );
buf ( n5431 , n1203 );
buf ( n5432 , n1688 );
buf ( n5433 , n876 );
buf ( n5434 , n8 );
buf ( n5435 , n1590 );
buf ( n5436 , n1305 );
buf ( n5437 , n747 );
buf ( n5438 , n1815 );
buf ( n5439 , n1318 );
buf ( n5440 , n750 );
buf ( n5441 , n380 );
buf ( n5442 , n1758 );
buf ( n5443 , n1871 );
buf ( n5444 , n771 );
buf ( n5445 , n742 );
buf ( n5446 , n967 );
buf ( n5447 , n603 );
buf ( n5448 , n1754 );
buf ( n5449 , n719 );
buf ( n5450 , n1194 );
buf ( n5451 , n133 );
buf ( n5452 , n1653 );
buf ( n5453 , n1492 );
buf ( n5454 , n353 );
buf ( n5455 , n1605 );
buf ( n5456 , n1852 );
buf ( n5457 , n49 );
buf ( n5458 , n656 );
buf ( n5459 , n2157 );
buf ( n5460 , n425 );
buf ( n5461 , n1739 );
buf ( n5462 , n839 );
buf ( n5463 , n1002 );
buf ( n5464 , n1927 );
buf ( n5465 , n144 );
buf ( n5466 , n960 );
buf ( n5467 , n1528 );
buf ( n5468 , n1091 );
buf ( n5469 , n1523 );
buf ( n5470 , n45 );
buf ( n5471 , n1135 );
buf ( n5472 , n1267 );
buf ( n5473 , n975 );
buf ( n5474 , n997 );
buf ( n5475 , n1189 );
buf ( n5476 , n1729 );
buf ( n5477 , n1959 );
buf ( n5478 , n242 );
buf ( n5479 , n1071 );
buf ( n5480 , n1613 );
buf ( n5481 , n321 );
buf ( n5482 , n1789 );
buf ( n5483 , n662 );
buf ( n5484 , n2063 );
buf ( n5485 , n1935 );
buf ( n5486 , n1129 );
buf ( n5487 , n1170 );
buf ( n5488 , n1694 );
buf ( n5489 , n1671 );
buf ( n5490 , n34 );
buf ( n5491 , n546 );
buf ( n5492 , n1236 );
buf ( n5493 , n799 );
buf ( n5494 , n553 );
buf ( n5495 , n127 );
buf ( n5496 , n1451 );
buf ( n5497 , n2161 );
buf ( n5498 , n207 );
buf ( n5499 , n2122 );
buf ( n5500 , n111 );
buf ( n5501 , n1698 );
buf ( n5502 , n875 );
buf ( n5503 , n23 );
buf ( n5504 , n182 );
buf ( n5505 , n866 );
buf ( n5506 , n474 );
buf ( n5507 , n877 );
buf ( n5508 , n307 );
buf ( n5509 , n1568 );
buf ( n5510 , n1064 );
buf ( n5511 , n1765 );
buf ( n5512 , n279 );
buf ( n5513 , n271 );
buf ( n5514 , n1110 );
buf ( n5515 , n1223 );
buf ( n5516 , n1018 );
buf ( n5517 , n139 );
buf ( n5518 , n1813 );
buf ( n5519 , n1545 );
buf ( n5520 , n1097 );
buf ( n5521 , n2121 );
buf ( n5522 , n134 );
buf ( n5523 , n695 );
buf ( n5524 , n2141 );
buf ( n5525 , n272 );
buf ( n5526 , n471 );
buf ( n5527 , n527 );
buf ( n5528 , n145 );
buf ( n5529 , n24 );
buf ( n5530 , n1087 );
buf ( n5531 , n1271 );
buf ( n5532 , n905 );
buf ( n5533 , n907 );
buf ( n5534 , n1182 );
buf ( n5535 , n2085 );
buf ( n5536 , n1362 );
buf ( n5537 , n273 );
buf ( n5538 , n1089 );
buf ( n5539 , n333 );
buf ( n5540 , n2032 );
buf ( n5541 , n281 );
buf ( n5542 , n1916 );
buf ( n5543 , n1122 );
buf ( n5544 , n558 );
buf ( n5545 , n1272 );
buf ( n5546 , n1243 );
buf ( n5547 , n1556 );
buf ( n5548 , n923 );
buf ( n5549 , n308 );
buf ( n5550 , n1764 );
buf ( n5551 , n56 );
buf ( n5552 , n1322 );
buf ( n5553 , n206 );
buf ( n5554 , n1785 );
buf ( n5555 , n560 );
buf ( n5556 , n255 );
buf ( n5557 , n1677 );
buf ( n5558 , n1931 );
buf ( n5559 , n453 );
buf ( n5560 , n1800 );
buf ( n5561 , n247 );
buf ( n5562 , n976 );
buf ( n5563 , n1743 );
buf ( n5564 , n1394 );
buf ( n5565 , n2027 );
buf ( n5566 , n2040 );
buf ( n5567 , n1172 );
buf ( n5568 , n1468 );
buf ( n5569 , n985 );
buf ( n5570 , n1547 );
buf ( n5571 , n421 );
buf ( n5572 , n950 );
buf ( n5573 , n365 );
buf ( n5574 , n802 );
buf ( n5575 , n1455 );
buf ( n5576 , n1500 );
buf ( n5577 , n1920 );
buf ( n5578 , n1176 );
buf ( n5579 , n1275 );
buf ( n5580 , n1302 );
buf ( n5581 , n758 );
buf ( n5582 , n59 );
buf ( n5583 , n1062 );
buf ( n5584 , n331 );
buf ( n5585 , n2114 );
buf ( n5586 , n312 );
buf ( n5587 , n1392 );
buf ( n5588 , n1336 );
buf ( n5589 , n1391 );
buf ( n5590 , n1035 );
buf ( n5591 , n1342 );
buf ( n5592 , n525 );
buf ( n5593 , n1324 );
buf ( n5594 , n1466 );
buf ( n5595 , n1204 );
buf ( n5596 , n1375 );
buf ( n5597 , n556 );
buf ( n5598 , n451 );
buf ( n5599 , n971 );
buf ( n5600 , n1262 );
buf ( n5601 , n427 );
buf ( n5602 , n847 );
buf ( n5603 , n961 );
buf ( n5604 , n1038 );
buf ( n5605 , n1762 );
buf ( n5606 , n1151 );
buf ( n5607 , n1300 );
buf ( n5608 , n1792 );
buf ( n5609 , n64 );
buf ( n5610 , n668 );
buf ( n5611 , n2137 );
buf ( n5612 , n3 );
buf ( n5613 , n2182 );
buf ( n5614 , n1174 );
buf ( n5615 , n1752 );
buf ( n5616 , n1319 );
buf ( n5617 , n1691 );
buf ( n5618 , n2154 );
buf ( n5619 , n391 );
buf ( n5620 , n1945 );
buf ( n5621 , n1600 );
buf ( n5622 , n1036 );
buf ( n5623 , n282 );
buf ( n5624 , n529 );
buf ( n5625 , n780 );
buf ( n5626 , n552 );
buf ( n5627 , n1242 );
buf ( n5628 , n1232 );
buf ( n5629 , n1573 );
buf ( n5630 , n369 );
buf ( n5631 , n682 );
buf ( n5632 , n1219 );
buf ( n5633 , n439 );
buf ( n5634 , n661 );
buf ( n5635 , n995 );
buf ( n5636 , n406 );
buf ( n5637 , n698 );
buf ( n5638 , n1678 );
buf ( n5639 , n90 );
buf ( n5640 , n1886 );
buf ( n5641 , n947 );
buf ( n5642 , n708 );
buf ( n5643 , n1797 );
buf ( n5644 , n267 );
buf ( n5645 , n570 );
buf ( n5646 , n1494 );
buf ( n5647 , n783 );
buf ( n5648 , n1530 );
buf ( n5649 , n1303 );
buf ( n5650 , n1479 );
buf ( n5651 , n131 );
buf ( n5652 , n440 );
buf ( n5653 , n1593 );
buf ( n5654 , n779 );
buf ( n5655 , n124 );
buf ( n5656 , n36 );
buf ( n5657 , n174 );
buf ( n5658 , n1725 );
buf ( n5659 , n1938 );
buf ( n5660 , n710 );
buf ( n5661 , n537 );
buf ( n5662 , n1716 );
buf ( n5663 , n346 );
buf ( n5664 , n926 );
buf ( n5665 , n1867 );
buf ( n5666 , n294 );
buf ( n5667 , n1985 );
buf ( n5668 , n931 );
buf ( n5669 , n580 );
buf ( n5670 , n1121 );
buf ( n5671 , n1385 );
buf ( n5672 , n351 );
buf ( n5673 , n1870 );
buf ( n5674 , n922 );
buf ( n5675 , n745 );
buf ( n5676 , n1424 );
buf ( n5677 , n957 );
buf ( n5678 , n1055 );
buf ( n5679 , n901 );
buf ( n5680 , n859 );
buf ( n5681 , n2102 );
buf ( n5682 , n919 );
buf ( n5683 , n1052 );
buf ( n5684 , n280 );
buf ( n5685 , n602 );
buf ( n5686 , n740 );
buf ( n5687 , n1180 );
buf ( n5688 , n1658 );
buf ( n5689 , n2135 );
buf ( n5690 , n915 );
buf ( n5691 , n1251 );
buf ( n5692 , n749 );
buf ( n5693 , n857 );
buf ( n5694 , n1651 );
buf ( n5695 , n1746 );
buf ( n5696 , n916 );
buf ( n5697 , n2080 );
buf ( n5698 , n356 );
buf ( n5699 , n257 );
buf ( n5700 , n208 );
buf ( n5701 , n496 );
buf ( n5702 , n79 );
buf ( n5703 , n2128 );
buf ( n5704 , n1420 );
buf ( n5705 , n1594 );
buf ( n5706 , n259 );
buf ( n5707 , n1202 );
buf ( n5708 , n483 );
buf ( n5709 , n1406 );
buf ( n5710 , n41 );
buf ( n5711 , n1782 );
buf ( n5712 , n1824 );
buf ( n5713 , n488 );
buf ( n5714 , n1148 );
buf ( n5715 , n1544 );
buf ( n5716 , n115 );
buf ( n5717 , n760 );
buf ( n5718 , n2022 );
buf ( n5719 , n1335 );
buf ( n5720 , n1371 );
buf ( n5721 , n38 );
buf ( n5722 , n687 );
buf ( n5723 , n1700 );
buf ( n5724 , n702 );
buf ( n5725 , n179 );
buf ( n5726 , n1733 );
buf ( n5727 , n646 );
buf ( n5728 , n1894 );
buf ( n5729 , n1281 );
buf ( n5730 , n1574 );
buf ( n5731 , n1720 );
buf ( n5732 , n1987 );
buf ( n5733 , n620 );
buf ( n5734 , n712 );
buf ( n5735 , n879 );
buf ( n5736 , n1178 );
buf ( n5737 , n1258 );
buf ( n5738 , n1080 );
buf ( n5739 , n1238 );
buf ( n5740 , n1181 );
buf ( n5741 , n1007 );
buf ( n5742 , n767 );
buf ( n5743 , n651 );
buf ( n5744 , n1706 );
buf ( n5745 , n404 );
buf ( n5746 , n1892 );
buf ( n5747 , n129 );
buf ( n5748 , n1428 );
buf ( n5749 , n1751 );
buf ( n5750 , n1137 );
buf ( n5751 , n47 );
buf ( n5752 , n1346 );
buf ( n5753 , n1266 );
buf ( n5754 , n786 );
buf ( n5755 , n1101 );
buf ( n5756 , n1539 );
buf ( n5757 , n1670 );
buf ( n5758 , n1095 );
buf ( n5759 , n78 );
buf ( n5760 , n193 );
buf ( n5761 , n862 );
buf ( n5762 , n727 );
buf ( n5763 , n909 );
buf ( n5764 , n1438 );
buf ( n5765 , n2001 );
buf ( n5766 , n1722 );
buf ( n5767 , n1586 );
buf ( n5768 , n1675 );
buf ( n5769 , n2110 );
buf ( n5770 , n925 );
buf ( n5771 , n180 );
buf ( n5772 , n692 );
buf ( n5773 , n136 );
buf ( n5774 , n1980 );
buf ( n5775 , n640 );
buf ( n5776 , n1100 );
buf ( n5777 , n1163 );
buf ( n5778 , n1796 );
buf ( n5779 , n39 );
buf ( n5780 , n1551 );
buf ( n5781 , n1521 );
buf ( n5782 , n1747 );
buf ( n5783 , n327 );
buf ( n5784 , n128 );
buf ( n5785 , n1488 );
buf ( n5786 , n2132 );
buf ( n5787 , n21 );
buf ( n5788 , n467 );
buf ( n5789 , n791 );
buf ( n5790 , n1786 );
buf ( n5791 , n1553 );
buf ( n5792 , n233 );
buf ( n5793 , n1310 );
buf ( n5794 , n1639 );
buf ( n5795 , n387 );
buf ( n5796 , n250 );
buf ( n5797 , n276 );
buf ( n5798 , n520 );
buf ( n5799 , n1069 );
buf ( n5800 , n1312 );
buf ( n5801 , n1025 );
buf ( n5802 , n734 );
buf ( n5803 , n2010 );
buf ( n5804 , n322 );
buf ( n5805 , n2172 );
buf ( n5806 , n2165 );
buf ( n5807 , n384 );
buf ( n5808 , n836 );
buf ( n5809 , n1029 );
buf ( n5810 , n106 );
buf ( n5811 , n1378 );
buf ( n5812 , n726 );
buf ( n5813 , n1471 );
buf ( n5814 , n1461 );
buf ( n5815 , n2016 );
buf ( n5816 , n1652 );
buf ( n5817 , n11 );
buf ( n5818 , n25 );
buf ( n5819 , n426 );
buf ( n5820 , n2037 );
buf ( n5821 , n1304 );
buf ( n5822 , n1914 );
buf ( n5823 , n1934 );
buf ( n5824 , n832 );
buf ( n5825 , n1624 );
buf ( n5826 , n355 );
buf ( n5827 , n1835 );
buf ( n5828 , n970 );
buf ( n5829 , n285 );
buf ( n5830 , n1229 );
buf ( n5831 , n315 );
buf ( n5832 , n319 );
buf ( n5833 , n1627 );
buf ( n5834 , n336 );
buf ( n5835 , n62 );
buf ( n5836 , n1003 );
buf ( n5837 , n1074 );
buf ( n5838 , n1183 );
buf ( n5839 , n1058 );
buf ( n5840 , n1808 );
buf ( n5841 , n1549 );
buf ( n5842 , n924 );
buf ( n5843 , n512 );
buf ( n5844 , n521 );
buf ( n5845 , n1891 );
buf ( n5846 , n354 );
buf ( n5847 , n861 );
buf ( n5848 , n171 );
buf ( n5849 , n2100 );
buf ( n5850 , n517 );
buf ( n5851 , n565 );
buf ( n5852 , n936 );
buf ( n5853 , n1255 );
buf ( n5854 , n358 );
buf ( n5855 , n393 );
buf ( n5856 , n264 );
buf ( n5857 , n126 );
buf ( n5858 , n1339 );
buf ( n5859 , n1535 );
buf ( n5860 , n618 );
buf ( n5861 , n2061 );
buf ( n5862 , n1644 );
buf ( n5863 , n1459 );
buf ( n5864 , n324 );
buf ( n5865 , n1589 );
buf ( n5866 , n1559 );
buf ( n5867 , n1068 );
buf ( n5868 , n1913 );
buf ( n5869 , n2123 );
buf ( n5870 , n1517 );
buf ( n5871 , n1447 );
buf ( n5872 , n480 );
buf ( n5873 , n1218 );
buf ( n5874 , n1949 );
buf ( n5875 , n1487 );
buf ( n5876 , n843 );
buf ( n5877 , n475 );
buf ( n5878 , n2142 );
buf ( n5879 , n477 );
buf ( n5880 , n1977 );
buf ( n5881 , n650 );
buf ( n5882 , n1667 );
buf ( n5883 , n1769 );
buf ( n5884 , n1640 );
buf ( n5885 , n1450 );
buf ( n5886 , n1734 );
buf ( n5887 , n619 );
buf ( n5888 , n350 );
buf ( n5889 , n1760 );
buf ( n5890 , n1510 );
buf ( n5891 , n1364 );
buf ( n5892 , n361 );
buf ( n5893 , n892 );
buf ( n5894 , n617 );
buf ( n5895 , n2104 );
buf ( n5896 , n1256 );
buf ( n5897 , n1006 );
buf ( n5898 , n655 );
buf ( n5899 , n1947 );
buf ( n5900 , n1241 );
buf ( n5901 , n1338 );
buf ( n5902 , n1365 );
buf ( n5903 , n614 );
buf ( n5904 , n2046 );
buf ( n5905 , n373 );
buf ( n5906 , n766 );
buf ( n5907 , n542 );
buf ( n5908 , n1214 );
buf ( n5909 , n431 );
buf ( n5910 , n1444 );
buf ( n5911 , n1790 );
buf ( n5912 , n1347 );
buf ( n5913 , n1113 );
buf ( n5914 , n2003 );
buf ( n5915 , n1878 );
buf ( n5916 , n2113 );
buf ( n5917 , n157 );
buf ( n5918 , n2026 );
buf ( n5919 , n578 );
buf ( n5920 , n14 );
buf ( n5921 , n1048 );
buf ( n5922 , n1133 );
buf ( n5923 , n16 );
buf ( n5924 , n1840 );
buf ( n5925 , n1414 );
buf ( n5926 , n416 );
buf ( n5927 , n1777 );
buf ( n5928 , n2036 );
buf ( n5929 , n1311 );
buf ( n5930 , n1088 );
buf ( n5931 , n989 );
buf ( n5932 , n403 );
buf ( n5933 , n680 );
buf ( n5934 , n362 );
buf ( n5935 , n1390 );
buf ( n5936 , n1453 );
buf ( n5937 , n1941 );
buf ( n5938 , n419 );
buf ( n5939 , n1084 );
buf ( n5940 , n1592 );
buf ( n5941 , n2 );
buf ( n5942 , n1096 );
buf ( n5943 , n539 );
buf ( n5944 , n2150 );
buf ( n5945 , n1778 );
buf ( n5946 , n643 );
buf ( n5947 , n1400 );
buf ( n5948 , n1713 );
buf ( n5949 , n1419 );
buf ( n5950 , n1915 );
buf ( n5951 , n10 );
buf ( n5952 , n292 );
buf ( n5953 , n1881 );
buf ( n5954 , n456 );
buf ( n5955 , n1426 );
buf ( n5956 , n2173 );
buf ( n5957 , n1106 );
buf ( n5958 , n657 );
buf ( n5959 , n463 );
buf ( n5960 , n258 );
buf ( n5961 , n773 );
buf ( n5962 , n377 );
buf ( n5963 , n932 );
buf ( n5964 , n2087 );
buf ( n5965 , n1446 );
buf ( n5966 , n572 );
buf ( n5967 , n196 );
buf ( n5968 , n1154 );
buf ( n5969 , n408 );
buf ( n5970 , n52 );
buf ( n5971 , n1429 );
buf ( n5972 , n73 );
buf ( n5973 , n1731 );
buf ( n5974 , n743 );
buf ( n5975 , n591 );
buf ( n5976 , n885 );
buf ( n5977 , n1168 );
buf ( n5978 , n94 );
buf ( n5979 , n1983 );
buf ( n5980 , n722 );
buf ( n5981 , n1629 );
buf ( n5982 , n1950 );
buf ( n5983 , n1138 );
buf ( n5984 , n798 );
buf ( n5985 , n2107 );
buf ( n5986 , n775 );
buf ( n5987 , n215 );
buf ( n5988 , n2033 );
buf ( n5989 , n805 );
buf ( n5990 , n1657 );
buf ( n5991 , n1681 );
buf ( n5992 , n400 );
buf ( n5993 , n1659 );
buf ( n5994 , n1661 );
buf ( n5995 , n1268 );
buf ( n5996 , n1323 );
buf ( n5997 , n1889 );
buf ( n5998 , n2155 );
buf ( n5999 , n647 );
buf ( n6000 , n1190 );
buf ( n6001 , n2171 );
buf ( n6002 , n216 );
buf ( n6003 , n1723 );
buf ( n6004 , n1703 );
buf ( n6005 , n198 );
buf ( n6006 , n2181 );
buf ( n6007 , n81 );
buf ( n6008 , n1277 );
buf ( n6009 , n1711 );
buf ( n6010 , n1861 );
buf ( n6011 , n238 );
buf ( n6012 , n538 );
buf ( n6013 , n1177 );
buf ( n6014 , n899 );
buf ( n6015 , n510 );
buf ( n6016 , n2098 );
buf ( n6017 , n31 );
buf ( n6018 , n1571 );
buf ( n6019 , n1583 );
buf ( n6020 , n375 );
buf ( n6021 , n683 );
buf ( n6022 , n685 );
buf ( n6023 , n1684 );
buf ( n6024 , n222 );
buf ( n6025 , n2086 );
buf ( n6026 , n551 );
buf ( n6027 , n1206 );
buf ( n6028 , n1701 );
buf ( n6029 , n1333 );
buf ( n6030 , n612 );
buf ( n6031 , n2145 );
buf ( n6032 , n181 );
buf ( n6033 , n1235 );
buf ( n6034 , n2079 );
buf ( n6035 , n929 );
buf ( n6036 , n808 );
buf ( n6037 , n910 );
buf ( n6038 , n1144 );
buf ( n6039 , n555 );
buf ( n6040 , n176 );
buf ( n6041 , n1811 );
buf ( n6042 , n713 );
buf ( n6043 , n2044 );
buf ( n6044 , n1755 );
buf ( n6045 , n736 );
buf ( n6046 , n1422 );
buf ( n6047 , n904 );
buf ( n6048 , n1458 );
buf ( n6049 , n1737 );
buf ( n6050 , n482 );
buf ( n6051 , n1668 );
buf ( n6052 , n366 );
buf ( n6053 , n1847 );
buf ( n6054 , n1532 );
buf ( n6055 , n2127 );
buf ( n6056 , n422 );
buf ( n6057 , n883 );
buf ( n6058 , n2030 );
buf ( n6059 , n1355 );
buf ( n6060 , n1078 );
buf ( n6061 , n1061 );
buf ( n6062 , n1580 );
buf ( n6063 , n1476 );
buf ( n6064 , n109 );
buf ( n6065 , n1398 );
buf ( n6066 , n491 );
buf ( n6067 , n806 );
buf ( n6068 , n795 );
buf ( n6069 , n838 );
buf ( n6070 , n1925 );
buf ( n6071 , n1377 );
buf ( n6072 , n2094 );
buf ( n6073 , n2160 );
buf ( n6074 , n1164 );
buf ( n6075 , n2126 );
buf ( n6076 , n1265 );
buf ( n6077 , n818 );
buf ( n6078 , n639 );
buf ( n6079 , n1462 );
buf ( n6080 , n625 );
buf ( n6081 , n2109 );
buf ( n6082 , n613 );
buf ( n6083 , n1843 );
buf ( n6084 , n2117 );
buf ( n6085 , n1936 );
buf ( n6086 , n1403 );
buf ( n6087 , n1 );
buf ( n6088 , n237 );
buf ( n6089 , n84 );
buf ( n6090 , n1351 );
buf ( n6091 , n717 );
buf ( n6092 , n1687 );
buf ( n6093 , n675 );
buf ( n6094 , n1702 );
buf ( n6095 , n121 );
buf ( n6096 , n1073 );
buf ( n6097 , n1850 );
buf ( n6098 , n627 );
buf ( n6099 , n637 );
buf ( n6100 , n1844 );
buf ( n6101 , n1230 );
buf ( n6102 , n1094 );
buf ( n6103 , n1158 );
buf ( n6104 , n244 );
buf ( n6105 , n70 );
buf ( n6106 , n187 );
buf ( n6107 , n1185 );
buf ( n6108 , n251 );
buf ( n6109 , n1680 );
buf ( n6110 , n585 );
buf ( n6111 , n1143 );
buf ( n6112 , n1112 );
buf ( n6113 , n706 );
buf ( n6114 , n1457 );
buf ( n6115 , n1166 );
buf ( n6116 , n1812 );
buf ( n6117 , n1115 );
buf ( n6118 , n1712 );
buf ( n6119 , n1252 );
buf ( n6120 , n1858 );
buf ( n6121 , n894 );
buf ( n6122 , n1127 );
buf ( n6123 , n1417 );
buf ( n6124 , n1066 );
buf ( n6125 , n1147 );
buf ( n6126 , n801 );
buf ( n6127 , n540 );
buf ( n6128 , n911 );
buf ( n6129 , n1601 );
buf ( n6130 , n1709 );
buf ( n6131 , n1295 );
buf ( n6132 , n1374 );
buf ( n6133 , n489 );
buf ( n6134 , n814 );
buf ( n6135 , n241 );
buf ( n6136 , n1830 );
buf ( n6137 , n1159 );
buf ( n6138 , n66 );
buf ( n6139 , n1849 );
buf ( n6140 , n2124 );
buf ( n6141 , n1888 );
buf ( n6142 , n1307 );
buf ( n6143 , n476 );
buf ( n6144 , n1081 );
buf ( n6145 , n418 );
buf ( n6146 , n1783 );
buf ( n6147 , n228 );
buf ( n6148 , n600 );
buf ( n6149 , n544 );
buf ( n6150 , n1284 );
buf ( n6151 , n562 );
buf ( n6152 , n1140 );
buf ( n6153 , n1669 );
buf ( n6154 , n2011 );
buf ( n6155 , n497 );
buf ( n6156 , n1146 );
buf ( n6157 , n940 );
buf ( n6158 , n2069 );
buf ( n6159 , n673 );
buf ( n6160 , n1724 );
buf ( n6161 , n872 );
buf ( n6162 , n1224 );
buf ( n6163 , n738 );
buf ( n6164 , n1814 );
buf ( n6165 , n735 );
buf ( n6166 , n2111 );
buf ( n6167 , n2034 );
buf ( n6168 , n224 );
buf ( n6169 , n43 );
buf ( n6170 , n125 );
buf ( n6171 , n1434 );
buf ( n6172 , n671 );
buf ( n6173 , n162 );
buf ( n6174 , n1050 );
buf ( n6175 , n1964 );
buf ( n6176 , n1608 );
buf ( n6177 , n1647 );
buf ( n6178 , n796 );
buf ( n6179 , n1930 );
buf ( n6180 , n1630 );
buf ( n6181 , n1334 );
buf ( n6182 , n821 );
buf ( n6183 , n197 );
buf ( n6184 , n993 );
buf ( n6185 , n2163 );
buf ( n6186 , n288 );
buf ( n6187 , n2156 );
buf ( n6188 , n991 );
buf ( n6189 , n218 );
buf ( n6190 , n507 );
buf ( n6191 , n1349 );
buf ( n6192 , n1237 );
buf ( n6193 , n2120 );
buf ( n6194 , n1259 );
buf ( n6195 , n797 );
buf ( n6196 , n443 );
buf ( n6197 , n2144 );
buf ( n6198 , n153 );
buf ( n6199 , n1042 );
buf ( n6200 , n381 );
buf ( n6201 , n104 );
buf ( n6202 , n1404 );
buf ( n6203 , n1205 );
buf ( n6204 , n1393 );
buf ( n6205 , n858 );
buf ( n6206 , n1834 );
buf ( n6207 , n1689 );
buf ( n6208 , n1954 );
buf ( n6209 , n1124 );
buf ( n6210 , n548 );
buf ( n6211 , n1719 );
buf ( n6212 , n938 );
buf ( n6213 , n522 );
buf ( n6214 , n470 );
buf ( n6215 , n1331 );
buf ( n6216 , n678 );
buf ( n6217 , n103 );
buf ( n6218 , n1279 );
buf ( n6219 , n1082 );
buf ( n6220 , n1554 );
buf ( n6221 , n199 );
buf ( n6222 , n1411 );
buf ( n6223 , n54 );
buf ( n6224 , n194 );
buf ( n6225 , n1317 );
buf ( n6226 , n1350 );
buf ( n6227 , n516 );
buf ( n6228 , n185 );
buf ( n6229 , n1369 );
buf ( n6230 , n1863 );
buf ( n6231 , n1839 );
buf ( n6232 , n897 );
buf ( n6233 , n1244 );
buf ( n6234 , n1519 );
buf ( n6235 , n1598 );
buf ( n6236 , n596 );
buf ( n6237 , n252 );
buf ( n6238 , n959 );
buf ( n6239 , n167 );
buf ( n6240 , n1373 );
buf ( n6241 , n820 );
buf ( n6242 , n1253 );
buf ( n6243 , n559 );
buf ( n6244 , n165 );
buf ( n6245 , n396 );
buf ( n6246 , n409 );
buf ( n6247 , n1313 );
buf ( n6248 , n2112 );
buf ( n6249 , n1676 );
buf ( n6250 , n1167 );
buf ( n6251 , n1998 );
buf ( n6252 , n1051 );
buf ( n6253 , n466 );
buf ( n6254 , n1978 );
buf ( n6255 , n1918 );
buf ( n6256 , n1626 );
buf ( n6257 , n446 );
buf ( n6258 , n1125 );
buf ( n6259 , n588 );
buf ( n6260 , n1485 );
buf ( n6261 , n112 );
buf ( n6262 , n1092 );
buf ( n6263 , n395 );
buf ( n6264 , n183 );
buf ( n6265 , n2147 );
buf ( n6266 , n748 );
buf ( n6267 , n117 );
buf ( n6268 , n390 );
buf ( n6269 , n823 );
buf ( n6270 , n896 );
buf ( n6271 , n2038 );
buf ( n6272 , n853 );
buf ( n6273 , n694 );
buf ( n6274 , n1902 );
buf ( n6275 , n1054 );
buf ( n6276 , n1803 );
buf ( n6277 , n769 );
buf ( n6278 , n330 );
buf ( n6279 , n1635 );
buf ( n6280 , n1866 );
buf ( n6281 , n1114 );
buf ( n6282 , n1460 );
buf ( n6283 , n1306 );
buf ( n6284 , n1512 );
buf ( n6285 , n1618 );
buf ( n6286 , n402 );
buf ( n6287 , n1329 );
buf ( n6288 , n1287 );
buf ( n6289 , n100 );
buf ( n6290 , n1718 );
buf ( n6291 , n1024 );
buf ( n6292 , n777 );
buf ( n6293 , n2072 );
buf ( n6294 , n1963 );
buf ( n6295 , n1211 );
buf ( n6296 , n1543 );
buf ( n6297 , n465 );
buf ( n6298 , n1727 );
buf ( n6299 , n611 );
buf ( n6300 , n1326 );
buf ( n6301 , n1372 );
buf ( n6302 , n1247 );
buf ( n6303 , n473 );
buf ( n6304 , n1682 );
buf ( n6305 , n1507 );
buf ( n6306 , n1320 );
buf ( n6307 , n752 );
buf ( n6308 , n1344 );
buf ( n6309 , n1473 );
buf ( n6310 , n1975 );
buf ( n6311 , n97 );
buf ( n6312 , n718 );
buf ( n6313 , n342 );
buf ( n6314 , n1388 );
buf ( n6315 , n83 );
buf ( n6316 , n37 );
buf ( n6317 , n912 );
buf ( n6318 , n644 );
buf ( n6319 , n1944 );
buf ( n6320 , n147 );
buf ( n6321 , n1437 );
buf ( n6322 , n535 );
buf ( n6323 , n2049 );
buf ( n6324 , n35 );
buf ( n6325 , n1105 );
buf ( n6326 , n1771 );
buf ( n6327 , n1017 );
buf ( n6328 , n424 );
buf ( n6329 , n1169 );
buf ( n6330 , n1382 );
buf ( n6331 , n1735 );
buf ( n6332 , n1557 );
buf ( n6333 , n1254 );
buf ( n6334 , n1633 );
buf ( n6335 , n1795 );
buf ( n6336 , n1857 );
buf ( n6337 , n1509 );
buf ( n6338 , n809 );
buf ( n6339 , n458 );
buf ( n6340 , n523 );
buf ( n6341 , n1234 );
buf ( n6342 , n1937 );
buf ( n6343 , n573 );
buf ( n6344 , n2091 );
buf ( n6345 , n1359 );
buf ( n6346 , n359 );
buf ( n6347 , n1470 );
buf ( n6348 , n1053 );
buf ( n6349 , n122 );
buf ( n6350 , n649 );
buf ( n6351 , n1449 );
buf ( n6352 , n1083 );
buf ( n6353 , n2019 );
buf ( n6354 , n586 );
buf ( n6355 , n574 );
buf ( n6356 , n44 );
buf ( n6357 , n1787 );
buf ( n6358 , n632 );
buf ( n6359 , n711 );
buf ( n6360 , n1798 );
buf ( n6361 , n28 );
buf ( n6362 , n417 );
buf ( n6363 , n1548 );
buf ( n6364 , n274 );
buf ( n6365 , n63 );
buf ( n6366 , n1988 );
buf ( n6367 , n2035 );
buf ( n6368 , n2002 );
buf ( n6369 , n1309 );
buf ( n6370 , n787 );
buf ( n6371 , n763 );
buf ( n6372 , n370 );
buf ( n6373 , n1570 );
buf ( n6374 , n790 );
buf ( n6375 , n1478 );
buf ( n6376 , n2084 );
buf ( n6377 , n515 );
buf ( n6378 , n2031 );
buf ( n6379 , n1484 );
buf ( n6380 , n1693 );
buf ( n6381 , n232 );
buf ( n6382 , n1890 );
buf ( n6383 , n1595 );
buf ( n6384 , n1240 );
buf ( n6385 , n1136 );
buf ( n6386 , n225 );
buf ( n6387 , n1021 );
buf ( n6388 , n1353 );
buf ( n6389 , n202 );
buf ( n6390 , n1200 );
buf ( n6391 , n1467 );
buf ( n6392 , n2089 );
buf ( n6393 , n941 );
buf ( n6394 , n481 );
buf ( n6395 , n1464 );
buf ( n6396 , n2143 );
buf ( n6397 , n1531 );
buf ( n6398 , n874 );
buf ( n6399 , n2131 );
buf ( n6400 , n545 );
buf ( n6401 , n1673 );
buf ( n6402 , n1325 );
buf ( n6403 , n1297 );
buf ( n6404 , n1389 );
buf ( n6405 , n869 );
buf ( n6406 , n227 );
buf ( n6407 , n166 );
buf ( n6408 , n2106 );
buf ( n6409 , n141 );
buf ( n6410 , n846 );
buf ( n6411 , n1619 );
buf ( n6412 , n1541 );
buf ( n6413 , n844 );
buf ( n6414 , n1060 );
buf ( n6415 , n567 );
buf ( n6416 , n1425 );
buf ( n6417 , n494 );
buf ( n6418 , n1775 );
buf ( n6419 , n223 );
buf ( n6420 , n454 );
buf ( n6421 , n1721 );
buf ( n6422 , n1150 );
buf ( n6423 , n1001 );
buf ( n6424 , n1940 );
buf ( n6425 , n908 );
buf ( n6426 , n1956 );
buf ( n6427 , n576 );
buf ( n6428 , n1848 );
buf ( n6429 , n1829 );
buf ( n6430 , n1482 );
buf ( n6431 , n1730 );
buf ( n6432 , n1011 );
buf ( n6433 , n2050 );
buf ( n6434 , n837 );
buf ( n6435 , n138 );
buf ( n6436 , n1903 );
buf ( n6437 , n1161 );
buf ( n6438 , n891 );
buf ( n6439 , n638 );
buf ( n6440 , n269 );
buf ( n6441 , n1536 );
buf ( n6442 , n203 );
buf ( n6443 , n582 );
buf ( n6444 , n1616 );
buf ( n6445 , n1958 );
buf ( n6446 , n1542 );
buf ( n6447 , n445 );
buf ( n6448 , n1714 );
buf ( n6449 , n1708 );
buf ( n6450 , n2068 );
buf ( n6451 , n487 );
buf ( n6452 , n200 );
buf ( n6453 , n275 );
buf ( n6454 , n1231 );
buf ( n6455 , n1939 );
buf ( n6456 , n1330 );
buf ( n6457 , n1506 );
buf ( n6458 , n118 );
buf ( n6459 , n945 );
buf ( n6460 , n1838 );
buf ( n6461 , n13 );
buf ( n6462 , n1924 );
buf ( n6463 , n2088 );
buf ( n6464 , n1294 );
buf ( n6465 , n1686 );
buf ( n6466 , n209 );
buf ( n6467 , n636 );
buf ( n6468 , n2053 );
buf ( n6469 , n942 );
buf ( n6470 , n792 );
buf ( n6471 , n1763 );
buf ( n6472 , n1376 );
buf ( n6473 , n1044 );
buf ( n6474 , n1576 );
buf ( n6475 , n490 );
buf ( n6476 , n96 );
buf ( n6477 , n1299 );
buf ( n6478 , n730 );
buf ( n6479 , n1753 );
buf ( n6480 , n2054 );
buf ( n6481 , n2045 );
buf ( n6482 , n566 );
buf ( n6483 , n107 );
buf ( n6484 , n334 );
buf ( n6485 , n204 );
buf ( n6486 , n2048 );
buf ( n6487 , n383 );
buf ( n6488 , n2103 );
buf ( n6489 , n900 );
buf ( n6490 , n1628 );
buf ( n6491 , n1504 );
buf ( n6492 , n1065 );
buf ( n6493 , n1384 );
buf ( n6494 , n987 );
buf ( n6495 , n1407 );
buf ( n6496 , n886 );
buf ( n6497 , n1337 );
buf ( n6498 , n1184 );
buf ( n6499 , n392 );
buf ( n6500 , n1511 );
buf ( n6501 , n1527 );
buf ( n6502 , n1837 );
buf ( n6503 , n1145 );
buf ( n6504 , n1356 );
buf ( n6505 , n1165 );
buf ( n6506 , n583 );
buf ( n6507 , n27 );
buf ( n6508 , n2185 );
buf ( n6509 , n306 );
buf ( n6510 , n2158 );
buf ( n6511 , n159 );
buf ( n6512 , n89 );
buf ( n6513 , n870 );
buf ( n6514 , n1966 );
buf ( n6515 , n690 );
buf ( n6516 , n597 );
buf ( n6517 , n635 );
buf ( n6518 , n1296 );
buf ( n6519 , n314 );
buf ( n6520 , n1409 );
buf ( n6521 , n438 );
buf ( n6522 , n983 );
buf ( n6523 , n1569 );
buf ( n6524 , n437 );
buf ( n6525 , n1565 );
buf ( n6526 , n739 );
buf ( n6527 , n1397 );
buf ( n6528 , n810 );
buf ( n6529 , n1490 );
buf ( n6530 , n728 );
buf ( n6531 , n686 );
buf ( n6532 , n1801 );
buf ( n6533 , n1227 );
buf ( n6534 , n450 );
buf ( n6535 , n1293 );
buf ( n6536 , n715 );
buf ( n6537 , n519 );
buf ( n6538 , n1779 );
buf ( n6539 , n1649 );
buf ( n6540 , n865 );
buf ( n6541 , n262 );
buf ( n6542 , n860 );
buf ( n6543 , n1495 );
buf ( n6544 , n998 );
buf ( n6545 , n1010 );
buf ( n6546 , n1860 );
buf ( n6547 , n1974 );
buf ( n6548 , n464 );
buf ( n6549 , n1770 );
buf ( n6550 , n1666 );
buf ( n6551 , n311 );
buf ( n6552 , n1611 );
buf ( n6553 , n6 );
buf ( n6554 , n291 );
buf ( n6555 , n2170 );
buf ( n6556 , n2065 );
buf ( n6557 , n2148 );
buf ( n6558 , n1660 );
buf ( n6559 , n781 );
buf ( n6560 , n459 );
buf ( n6561 , n1503 );
buf ( n6562 , n46 );
buf ( n6563 , n917 );
buf ( n6564 , n1928 );
buf ( n6565 , n1540 );
buf ( n6566 , n99 );
buf ( n6567 , n1728 );
buf ( n6568 , n48 );
buf ( n6569 , n679 );
buf ( n6570 , n372 );
buf ( n6571 , n2057 );
buf ( n6572 , n1118 );
buf ( n6573 , n2029 );
buf ( n6574 , n1774 );
buf ( n6575 , n1851 );
buf ( n6576 , n903 );
buf ( n6577 , n2164 );
buf ( n6578 , n1430 );
buf ( n6579 , n693 );
buf ( n6580 , n4394 );
buf ( n6581 , n6580 );
not ( n6582 , n6581 );
buf ( n6583 , n4395 );
buf ( n6584 , n6583 );
not ( n6585 , n6584 );
buf ( n6586 , n4396 );
not ( n6587 , n6586 );
not ( n6588 , n6587 );
or ( n6589 , n6585 , n6588 );
not ( n6590 , n6583 );
buf ( n6591 , n6586 );
nand ( n6592 , n6590 , n6591 );
nand ( n6593 , n6589 , n6592 );
buf ( n6594 , n4397 );
buf ( n6595 , n6594 );
and ( n6596 , n6593 , n6595 );
not ( n6597 , n6593 );
not ( n6598 , n6594 );
and ( n6599 , n6597 , n6598 );
nor ( n6600 , n6596 , n6599 );
buf ( n6601 , n4398 );
not ( n6602 , n6601 );
buf ( n6603 , n4399 );
nand ( n6604 , n6602 , n6603 );
not ( n6605 , n6604 );
buf ( n6606 , n6605 );
buf ( n6607 , n6606 );
buf ( n6608 , n6607 );
buf ( n6609 , n4400 );
nand ( n6610 , n6608 , n6609 );
buf ( n6611 , n4401 );
not ( n6612 , n6611 );
and ( n6613 , n6610 , n6612 );
not ( n6614 , n6610 );
buf ( n6615 , n6611 );
and ( n6616 , n6614 , n6615 );
nor ( n6617 , n6613 , n6616 );
not ( n6618 , n6617 );
xor ( n6619 , n6600 , n6618 );
buf ( n6620 , n6605 );
buf ( n6621 , n6620 );
buf ( n6622 , n6621 );
buf ( n6623 , n4402 );
nand ( n6624 , n6622 , n6623 );
buf ( n6625 , n4403 );
buf ( n6626 , n6625 );
and ( n6627 , n6624 , n6626 );
not ( n6628 , n6624 );
not ( n6629 , n6625 );
and ( n6630 , n6628 , n6629 );
nor ( n6631 , n6627 , n6630 );
buf ( n6632 , n6631 );
xor ( n6633 , n6619 , n6632 );
not ( n6634 , n6633 );
not ( n6635 , n6634 );
or ( n6636 , n6582 , n6635 );
xor ( n6637 , n6600 , n6631 );
xnor ( n6638 , n6637 , n6617 );
not ( n6639 , n6638 );
or ( n6640 , n6639 , n6581 );
nand ( n6641 , n6636 , n6640 );
not ( n6642 , n6641 );
buf ( n6643 , n4404 );
buf ( n6644 , n6643 );
not ( n6645 , n6644 );
buf ( n6646 , n4405 );
not ( n6647 , n6646 );
not ( n6648 , n6647 );
or ( n6649 , n6645 , n6648 );
not ( n6650 , n6643 );
buf ( n6651 , n6646 );
nand ( n6652 , n6650 , n6651 );
nand ( n6653 , n6649 , n6652 );
not ( n6654 , n6653 );
buf ( n6655 , n4406 );
buf ( n6656 , n4407 );
xor ( n6657 , n6655 , n6656 );
buf ( n6658 , n6605 );
buf ( n6659 , n6658 );
buf ( n6660 , n6659 );
buf ( n6661 , n4408 );
nand ( n6662 , n6660 , n6661 );
buf ( n6663 , n4409 );
not ( n6664 , n6663 );
and ( n6665 , n6662 , n6664 );
not ( n6666 , n6662 );
buf ( n6667 , n6663 );
and ( n6668 , n6666 , n6667 );
nor ( n6669 , n6665 , n6668 );
xnor ( n6670 , n6657 , n6669 );
not ( n6671 , n6670 );
or ( n6672 , n6654 , n6671 );
not ( n6673 , n6670 );
not ( n6674 , n6653 );
nand ( n6675 , n6673 , n6674 );
nand ( n6676 , n6672 , n6675 );
not ( n6677 , n6676 );
buf ( n6678 , n6677 );
not ( n6679 , n6678 );
or ( n6680 , n6642 , n6679 );
not ( n6681 , n6641 );
not ( n6682 , n6677 );
nand ( n6683 , n6681 , n6682 );
nand ( n6684 , n6680 , n6683 );
not ( n6685 , n6684 );
buf ( n6686 , n4410 );
not ( n6687 , n6686 );
buf ( n6688 , n4411 );
buf ( n6689 , n6688 );
not ( n6690 , n6689 );
buf ( n6691 , n4412 );
not ( n6692 , n6691 );
not ( n6693 , n6692 );
or ( n6694 , n6690 , n6693 );
not ( n6695 , n6688 );
buf ( n6696 , n6691 );
nand ( n6697 , n6695 , n6696 );
nand ( n6698 , n6694 , n6697 );
buf ( n6699 , n4413 );
not ( n6700 , n6699 );
and ( n6701 , n6698 , n6700 );
not ( n6702 , n6698 );
buf ( n6703 , n6699 );
and ( n6704 , n6702 , n6703 );
nor ( n6705 , n6701 , n6704 );
buf ( n6706 , n6621 );
buf ( n6707 , n4414 );
nand ( n6708 , n6706 , n6707 );
buf ( n6709 , n4415 );
buf ( n6710 , n6709 );
and ( n6711 , n6708 , n6710 );
not ( n6712 , n6708 );
not ( n6713 , n6709 );
and ( n6714 , n6712 , n6713 );
nor ( n6715 , n6711 , n6714 );
xor ( n6716 , n6705 , n6715 );
buf ( n6717 , n4416 );
nand ( n6718 , n6706 , n6717 );
buf ( n6719 , n4417 );
buf ( n6720 , n6719 );
and ( n6721 , n6718 , n6720 );
not ( n6722 , n6718 );
not ( n6723 , n6719 );
and ( n6724 , n6722 , n6723 );
nor ( n6725 , n6721 , n6724 );
not ( n6726 , n6725 );
xnor ( n6727 , n6716 , n6726 );
not ( n6728 , n6727 );
or ( n6729 , n6687 , n6728 );
or ( n6730 , n6727 , n6686 );
nand ( n6731 , n6729 , n6730 );
buf ( n6732 , n4418 );
buf ( n6733 , n6732 );
not ( n6734 , n6733 );
buf ( n6735 , n4419 );
not ( n6736 , n6735 );
not ( n6737 , n6736 );
or ( n6738 , n6734 , n6737 );
not ( n6739 , n6732 );
buf ( n6740 , n6735 );
nand ( n6741 , n6739 , n6740 );
nand ( n6742 , n6738 , n6741 );
buf ( n6743 , n4420 );
not ( n6744 , n6743 );
and ( n6745 , n6742 , n6744 );
not ( n6746 , n6742 );
buf ( n6747 , n6743 );
and ( n6748 , n6746 , n6747 );
nor ( n6749 , n6745 , n6748 );
buf ( n6750 , n4421 );
nand ( n6751 , n6706 , n6750 );
buf ( n6752 , n4422 );
buf ( n6753 , n6752 );
and ( n6754 , n6751 , n6753 );
not ( n6755 , n6751 );
not ( n6756 , n6752 );
and ( n6757 , n6755 , n6756 );
nor ( n6758 , n6754 , n6757 );
xor ( n6759 , n6749 , n6758 );
buf ( n6760 , n6606 );
buf ( n6761 , n6760 );
buf ( n6762 , n4423 );
nand ( n6763 , n6761 , n6762 );
buf ( n6764 , n4424 );
not ( n6765 , n6764 );
and ( n6766 , n6763 , n6765 );
not ( n6767 , n6763 );
buf ( n6768 , n6764 );
and ( n6769 , n6767 , n6768 );
nor ( n6770 , n6766 , n6769 );
xnor ( n6771 , n6759 , n6770 );
buf ( n6772 , n6771 );
buf ( n6773 , n6772 );
and ( n6774 , n6731 , n6773 );
not ( n6775 , n6731 );
not ( n6776 , n6772 );
and ( n6777 , n6775 , n6776 );
nor ( n6778 , n6774 , n6777 );
not ( n6779 , n6778 );
nand ( n6780 , n6685 , n6779 );
not ( n6781 , n6780 );
buf ( n6782 , n4425 );
buf ( n6783 , n6782 );
not ( n6784 , n6783 );
buf ( n6785 , n4426 );
buf ( n6786 , n6785 );
not ( n6787 , n6786 );
buf ( n6788 , n4427 );
not ( n6789 , n6788 );
not ( n6790 , n6789 );
or ( n6791 , n6787 , n6790 );
not ( n6792 , n6785 );
buf ( n6793 , n6788 );
nand ( n6794 , n6792 , n6793 );
nand ( n6795 , n6791 , n6794 );
buf ( n6796 , n4428 );
buf ( n6797 , n6796 );
and ( n6798 , n6795 , n6797 );
not ( n6799 , n6795 );
not ( n6800 , n6796 );
and ( n6801 , n6799 , n6800 );
nor ( n6802 , n6798 , n6801 );
buf ( n6803 , n6620 );
buf ( n6804 , n6803 );
buf ( n6805 , n4429 );
nand ( n6806 , n6804 , n6805 );
buf ( n6807 , n4430 );
buf ( n6808 , n6807 );
and ( n6809 , n6806 , n6808 );
not ( n6810 , n6806 );
not ( n6811 , n6807 );
and ( n6812 , n6810 , n6811 );
nor ( n6813 , n6809 , n6812 );
xor ( n6814 , n6802 , n6813 );
buf ( n6815 , n6658 );
buf ( n6816 , n6815 );
buf ( n6817 , n6816 );
buf ( n6818 , n4431 );
nand ( n6819 , n6817 , n6818 );
buf ( n6820 , n4432 );
buf ( n6821 , n6820 );
and ( n6822 , n6819 , n6821 );
not ( n6823 , n6819 );
not ( n6824 , n6820 );
and ( n6825 , n6823 , n6824 );
nor ( n6826 , n6822 , n6825 );
xnor ( n6827 , n6814 , n6826 );
buf ( n6828 , n6827 );
not ( n6829 , n6828 );
or ( n6830 , n6784 , n6829 );
or ( n6831 , n6828 , n6783 );
nand ( n6832 , n6830 , n6831 );
buf ( n6833 , n4433 );
buf ( n6834 , n6833 );
not ( n6835 , n6834 );
buf ( n6836 , n4434 );
not ( n6837 , n6836 );
not ( n6838 , n6837 );
or ( n6839 , n6835 , n6838 );
not ( n6840 , n6833 );
buf ( n6841 , n6836 );
nand ( n6842 , n6840 , n6841 );
nand ( n6843 , n6839 , n6842 );
buf ( n6844 , n4435 );
buf ( n6845 , n6844 );
and ( n6846 , n6843 , n6845 );
not ( n6847 , n6843 );
not ( n6848 , n6844 );
and ( n6849 , n6847 , n6848 );
nor ( n6850 , n6846 , n6849 );
buf ( n6851 , n6815 );
buf ( n6852 , n4436 );
nand ( n6853 , n6851 , n6852 );
buf ( n6854 , n4437 );
buf ( n6855 , n6854 );
and ( n6856 , n6853 , n6855 );
not ( n6857 , n6853 );
not ( n6858 , n6854 );
and ( n6859 , n6857 , n6858 );
nor ( n6860 , n6856 , n6859 );
xor ( n6861 , n6850 , n6860 );
buf ( n6862 , n6605 );
buf ( n6863 , n6862 );
buf ( n6864 , n4438 );
nand ( n6865 , n6863 , n6864 );
buf ( n6866 , n4439 );
buf ( n6867 , n6866 );
and ( n6868 , n6865 , n6867 );
not ( n6869 , n6865 );
not ( n6870 , n6866 );
and ( n6871 , n6869 , n6870 );
nor ( n6872 , n6868 , n6871 );
xor ( n6873 , n6861 , n6872 );
not ( n6874 , n6873 );
and ( n6875 , n6832 , n6874 );
not ( n6876 , n6832 );
not ( n6877 , n6874 );
and ( n6878 , n6876 , n6877 );
nor ( n6879 , n6875 , n6878 );
not ( n6880 , n6879 );
not ( n6881 , n6880 );
and ( n6882 , n6781 , n6881 );
and ( n6883 , n6780 , n6880 );
nor ( n6884 , n6882 , n6883 );
not ( n6885 , n6884 );
not ( n6886 , n6885 );
buf ( n6887 , n4440 );
buf ( n6888 , n6887 );
not ( n6889 , n6888 );
buf ( n6890 , n4441 );
buf ( n6891 , n6890 );
buf ( n6892 , n4442 );
not ( n6893 , n6892 );
buf ( n6894 , n4443 );
buf ( n6895 , n6894 );
and ( n6896 , n6893 , n6895 );
not ( n6897 , n6893 );
not ( n6898 , n6894 );
and ( n6899 , n6897 , n6898 );
nor ( n6900 , n6896 , n6899 );
xor ( n6901 , n6891 , n6900 );
buf ( n6902 , n4444 );
buf ( n6903 , n4445 );
xor ( n6904 , n6902 , n6903 );
buf ( n6905 , n6815 );
buf ( n6906 , n6905 );
buf ( n6907 , n4446 );
nand ( n6908 , n6906 , n6907 );
xnor ( n6909 , n6904 , n6908 );
xor ( n6910 , n6901 , n6909 );
not ( n6911 , n6910 );
or ( n6912 , n6889 , n6911 );
or ( n6913 , n6910 , n6888 );
nand ( n6914 , n6912 , n6913 );
buf ( n6915 , n4447 );
buf ( n6916 , n6915 );
not ( n6917 , n6916 );
buf ( n6918 , n4448 );
not ( n6919 , n6918 );
not ( n6920 , n6919 );
or ( n6921 , n6917 , n6920 );
not ( n6922 , n6915 );
buf ( n6923 , n6918 );
nand ( n6924 , n6922 , n6923 );
nand ( n6925 , n6921 , n6924 );
buf ( n6926 , n4449 );
not ( n6927 , n6926 );
and ( n6928 , n6925 , n6927 );
not ( n6929 , n6925 );
buf ( n6930 , n6926 );
and ( n6931 , n6929 , n6930 );
nor ( n6932 , n6928 , n6931 );
buf ( n6933 , n6620 );
buf ( n6934 , n6933 );
buf ( n6935 , n4450 );
nand ( n6936 , n6934 , n6935 );
buf ( n6937 , n4451 );
buf ( n6938 , n6937 );
and ( n6939 , n6936 , n6938 );
not ( n6940 , n6936 );
not ( n6941 , n6937 );
and ( n6942 , n6940 , n6941 );
nor ( n6943 , n6939 , n6942 );
xor ( n6944 , n6932 , n6943 );
buf ( n6945 , n6851 );
buf ( n6946 , n4452 );
nand ( n6947 , n6945 , n6946 );
buf ( n6948 , n4453 );
buf ( n6949 , n6948 );
and ( n6950 , n6947 , n6949 );
not ( n6951 , n6947 );
not ( n6952 , n6948 );
and ( n6953 , n6951 , n6952 );
nor ( n6954 , n6950 , n6953 );
xnor ( n6955 , n6944 , n6954 );
buf ( n6956 , n6955 );
not ( n6957 , n6956 );
and ( n6958 , n6914 , n6957 );
not ( n6959 , n6914 );
not ( n6960 , n6956 );
not ( n6961 , n6960 );
and ( n6962 , n6959 , n6961 );
nor ( n6963 , n6958 , n6962 );
buf ( n6964 , n4454 );
buf ( n6965 , n6964 );
not ( n6966 , n6965 );
buf ( n6967 , n4455 );
buf ( n6968 , n6967 );
not ( n6969 , n6968 );
buf ( n6970 , n4456 );
not ( n6971 , n6970 );
not ( n6972 , n6971 );
or ( n6973 , n6969 , n6972 );
not ( n6974 , n6967 );
buf ( n6975 , n6970 );
nand ( n6976 , n6974 , n6975 );
nand ( n6977 , n6973 , n6976 );
buf ( n6978 , n4457 );
not ( n6979 , n6978 );
and ( n6980 , n6977 , n6979 );
not ( n6981 , n6977 );
buf ( n6982 , n6978 );
and ( n6983 , n6981 , n6982 );
nor ( n6984 , n6980 , n6983 );
buf ( n6985 , n6621 );
buf ( n6986 , n4458 );
nand ( n6987 , n6985 , n6986 );
buf ( n6988 , n4459 );
buf ( n6989 , n6988 );
and ( n6990 , n6987 , n6989 );
not ( n6991 , n6987 );
not ( n6992 , n6988 );
and ( n6993 , n6991 , n6992 );
nor ( n6994 , n6990 , n6993 );
xor ( n6995 , n6984 , n6994 );
buf ( n6996 , n6622 );
buf ( n6997 , n4460 );
nand ( n6998 , n6996 , n6997 );
buf ( n6999 , n4461 );
not ( n7000 , n6999 );
and ( n7001 , n6998 , n7000 );
not ( n7002 , n6998 );
buf ( n7003 , n6999 );
and ( n7004 , n7002 , n7003 );
nor ( n7005 , n7001 , n7004 );
xnor ( n7006 , n6995 , n7005 );
not ( n7007 , n7006 );
or ( n7008 , n6966 , n7007 );
not ( n7009 , n6965 );
not ( n7010 , n6994 );
xor ( n7011 , n6984 , n7010 );
xnor ( n7012 , n7011 , n7005 );
nand ( n7013 , n7009 , n7012 );
nand ( n7014 , n7008 , n7013 );
buf ( n7015 , n4462 );
buf ( n7016 , n7015 );
not ( n7017 , n7016 );
buf ( n7018 , n4463 );
not ( n7019 , n7018 );
not ( n7020 , n7019 );
or ( n7021 , n7017 , n7020 );
not ( n7022 , n7015 );
buf ( n7023 , n7018 );
nand ( n7024 , n7022 , n7023 );
nand ( n7025 , n7021 , n7024 );
buf ( n7026 , n4464 );
buf ( n7027 , n7026 );
and ( n7028 , n7025 , n7027 );
not ( n7029 , n7025 );
not ( n7030 , n7026 );
and ( n7031 , n7029 , n7030 );
nor ( n7032 , n7028 , n7031 );
buf ( n7033 , n4465 );
nand ( n7034 , n6607 , n7033 );
buf ( n7035 , n4466 );
buf ( n7036 , n7035 );
and ( n7037 , n7034 , n7036 );
not ( n7038 , n7034 );
not ( n7039 , n7035 );
and ( n7040 , n7038 , n7039 );
nor ( n7041 , n7037 , n7040 );
xor ( n7042 , n7032 , n7041 );
buf ( n7043 , n6621 );
buf ( n7044 , n4467 );
nand ( n7045 , n7043 , n7044 );
buf ( n7046 , n4468 );
not ( n7047 , n7046 );
and ( n7048 , n7045 , n7047 );
not ( n7049 , n7045 );
buf ( n7050 , n7046 );
and ( n7051 , n7049 , n7050 );
nor ( n7052 , n7048 , n7051 );
xor ( n7053 , n7042 , n7052 );
not ( n7054 , n7053 );
not ( n7055 , n7054 );
and ( n7056 , n7014 , n7055 );
not ( n7057 , n7014 );
and ( n7058 , n7057 , n7054 );
nor ( n7059 , n7056 , n7058 );
not ( n7060 , n7059 );
nand ( n7061 , n6963 , n7060 );
not ( n7062 , n7061 );
buf ( n7063 , n4469 );
buf ( n7064 , n4470 );
buf ( n7065 , n7064 );
not ( n7066 , n7065 );
buf ( n7067 , n4471 );
not ( n7068 , n7067 );
not ( n7069 , n7068 );
or ( n7070 , n7066 , n7069 );
not ( n7071 , n7064 );
buf ( n7072 , n7067 );
nand ( n7073 , n7071 , n7072 );
nand ( n7074 , n7070 , n7073 );
buf ( n7075 , n4472 );
buf ( n7076 , n7075 );
and ( n7077 , n7074 , n7076 );
not ( n7078 , n7074 );
not ( n7079 , n7075 );
and ( n7080 , n7078 , n7079 );
nor ( n7081 , n7077 , n7080 );
buf ( n7082 , n6933 );
buf ( n7083 , n4473 );
nand ( n7084 , n7082 , n7083 );
buf ( n7085 , n4474 );
buf ( n7086 , n7085 );
and ( n7087 , n7084 , n7086 );
not ( n7088 , n7084 );
not ( n7089 , n7085 );
and ( n7090 , n7088 , n7089 );
nor ( n7091 , n7087 , n7090 );
xor ( n7092 , n7081 , n7091 );
buf ( n7093 , n6620 );
buf ( n7094 , n7093 );
buf ( n7095 , n4475 );
nand ( n7096 , n7094 , n7095 );
buf ( n7097 , n4476 );
buf ( n7098 , n7097 );
and ( n7099 , n7096 , n7098 );
not ( n7100 , n7096 );
not ( n7101 , n7097 );
and ( n7102 , n7100 , n7101 );
nor ( n7103 , n7099 , n7102 );
not ( n7104 , n7103 );
xnor ( n7105 , n7092 , n7104 );
xor ( n7106 , n7063 , n7105 );
buf ( n7107 , n4477 );
buf ( n7108 , n7107 );
not ( n7109 , n7108 );
buf ( n7110 , n4478 );
not ( n7111 , n7110 );
not ( n7112 , n7111 );
or ( n7113 , n7109 , n7112 );
not ( n7114 , n7107 );
buf ( n7115 , n7110 );
nand ( n7116 , n7114 , n7115 );
nand ( n7117 , n7113 , n7116 );
buf ( n7118 , n4479 );
buf ( n7119 , n7118 );
and ( n7120 , n7117 , n7119 );
not ( n7121 , n7117 );
not ( n7122 , n7118 );
and ( n7123 , n7121 , n7122 );
nor ( n7124 , n7120 , n7123 );
buf ( n7125 , n6658 );
buf ( n7126 , n7125 );
buf ( n7127 , n4480 );
nand ( n7128 , n7126 , n7127 );
buf ( n7129 , n4481 );
xor ( n7130 , n7128 , n7129 );
xor ( n7131 , n7124 , n7130 );
buf ( n7132 , n6605 );
buf ( n7133 , n7132 );
buf ( n7134 , n7133 );
buf ( n7135 , n4482 );
nand ( n7136 , n7134 , n7135 );
buf ( n7137 , n4483 );
buf ( n7138 , n7137 );
and ( n7139 , n7136 , n7138 );
not ( n7140 , n7136 );
not ( n7141 , n7137 );
and ( n7142 , n7140 , n7141 );
nor ( n7143 , n7139 , n7142 );
xnor ( n7144 , n7131 , n7143 );
xnor ( n7145 , n7106 , n7144 );
not ( n7146 , n7145 );
and ( n7147 , n7062 , n7146 );
not ( n7148 , n7059 );
nand ( n7149 , n7148 , n6963 );
and ( n7150 , n7149 , n7145 );
nor ( n7151 , n7147 , n7150 );
nand ( n7152 , n6684 , n6879 );
buf ( n7153 , n4484 );
nand ( n7154 , n6706 , n7153 );
buf ( n7155 , n4485 );
buf ( n7156 , n7155 );
and ( n7157 , n7154 , n7156 );
not ( n7158 , n7154 );
not ( n7159 , n7155 );
and ( n7160 , n7158 , n7159 );
nor ( n7161 , n7157 , n7160 );
buf ( n7162 , n7161 );
not ( n7163 , n7162 );
buf ( n7164 , n4486 );
buf ( n7165 , n7164 );
not ( n7166 , n7165 );
buf ( n7167 , n4487 );
not ( n7168 , n7167 );
not ( n7169 , n7168 );
or ( n7170 , n7166 , n7169 );
not ( n7171 , n7164 );
buf ( n7172 , n7167 );
nand ( n7173 , n7171 , n7172 );
nand ( n7174 , n7170 , n7173 );
buf ( n7175 , n4488 );
buf ( n7176 , n7175 );
and ( n7177 , n7174 , n7176 );
not ( n7178 , n7174 );
not ( n7179 , n7175 );
and ( n7180 , n7178 , n7179 );
nor ( n7181 , n7177 , n7180 );
not ( n7182 , n7181 );
buf ( n7183 , n7125 );
buf ( n7184 , n7183 );
buf ( n7185 , n4489 );
nand ( n7186 , n7184 , n7185 );
buf ( n7187 , n4490 );
not ( n7188 , n7187 );
and ( n7189 , n7186 , n7188 );
not ( n7190 , n7186 );
buf ( n7191 , n7187 );
and ( n7192 , n7190 , n7191 );
nor ( n7193 , n7189 , n7192 );
xor ( n7194 , n7182 , n7193 );
buf ( n7195 , n6620 );
buf ( n7196 , n7195 );
buf ( n7197 , n4491 );
nand ( n7198 , n7196 , n7197 );
buf ( n7199 , n4492 );
buf ( n7200 , n7199 );
and ( n7201 , n7198 , n7200 );
not ( n7202 , n7198 );
not ( n7203 , n7199 );
and ( n7204 , n7202 , n7203 );
nor ( n7205 , n7201 , n7204 );
not ( n7206 , n7205 );
xnor ( n7207 , n7194 , n7206 );
not ( n7208 , n7207 );
or ( n7209 , n7163 , n7208 );
or ( n7210 , n7207 , n7162 );
nand ( n7211 , n7209 , n7210 );
buf ( n7212 , n4493 );
buf ( n7213 , n7212 );
not ( n7214 , n7213 );
buf ( n7215 , n4494 );
not ( n7216 , n7215 );
not ( n7217 , n7216 );
or ( n7218 , n7214 , n7217 );
not ( n7219 , n7212 );
buf ( n7220 , n7215 );
nand ( n7221 , n7219 , n7220 );
nand ( n7222 , n7218 , n7221 );
buf ( n7223 , n4495 );
not ( n7224 , n7223 );
and ( n7225 , n7222 , n7224 );
not ( n7226 , n7222 );
buf ( n7227 , n7223 );
and ( n7228 , n7226 , n7227 );
nor ( n7229 , n7225 , n7228 );
buf ( n7230 , n6659 );
buf ( n7231 , n4496 );
nand ( n7232 , n7230 , n7231 );
buf ( n7233 , n4497 );
buf ( n7234 , n7233 );
and ( n7235 , n7232 , n7234 );
not ( n7236 , n7232 );
not ( n7237 , n7233 );
and ( n7238 , n7236 , n7237 );
nor ( n7239 , n7235 , n7238 );
xor ( n7240 , n7229 , n7239 );
buf ( n7241 , n4498 );
nand ( n7242 , n7184 , n7241 );
buf ( n7243 , n4499 );
not ( n7244 , n7243 );
and ( n7245 , n7242 , n7244 );
not ( n7246 , n7242 );
buf ( n7247 , n7243 );
and ( n7248 , n7246 , n7247 );
nor ( n7249 , n7245 , n7248 );
xnor ( n7250 , n7240 , n7249 );
not ( n7251 , n7250 );
buf ( n7252 , n7251 );
and ( n7253 , n7211 , n7252 );
not ( n7254 , n7211 );
not ( n7255 , n7250 );
not ( n7256 , n7255 );
and ( n7257 , n7254 , n7256 );
nor ( n7258 , n7253 , n7257 );
buf ( n7259 , n7258 );
not ( n7260 , n7259 );
and ( n7261 , n7152 , n7260 );
not ( n7262 , n7152 );
and ( n7263 , n7262 , n7259 );
nor ( n7264 , n7261 , n7263 );
or ( n7265 , n7151 , n7264 );
nand ( n7266 , n7264 , n7151 );
nand ( n7267 , n7265 , n7266 );
buf ( n7268 , n4500 );
buf ( n7269 , n7268 );
buf ( n7270 , n4501 );
buf ( n7271 , n7270 );
not ( n7272 , n7271 );
buf ( n7273 , n4502 );
not ( n7274 , n7273 );
not ( n7275 , n7274 );
or ( n7276 , n7272 , n7275 );
not ( n7277 , n7270 );
buf ( n7278 , n7273 );
nand ( n7279 , n7277 , n7278 );
nand ( n7280 , n7276 , n7279 );
buf ( n7281 , n4503 );
buf ( n7282 , n7281 );
and ( n7283 , n7280 , n7282 );
not ( n7284 , n7280 );
not ( n7285 , n7281 );
and ( n7286 , n7284 , n7285 );
nor ( n7287 , n7283 , n7286 );
buf ( n7288 , n6815 );
buf ( n7289 , n4504 );
nand ( n7290 , n7288 , n7289 );
buf ( n7291 , n4505 );
buf ( n7292 , n7291 );
and ( n7293 , n7290 , n7292 );
not ( n7294 , n7290 );
not ( n7295 , n7291 );
and ( n7296 , n7294 , n7295 );
nor ( n7297 , n7293 , n7296 );
xor ( n7298 , n7287 , n7297 );
buf ( n7299 , n6659 );
buf ( n7300 , n4506 );
nand ( n7301 , n7299 , n7300 );
buf ( n7302 , n4507 );
buf ( n7303 , n7302 );
and ( n7304 , n7301 , n7303 );
not ( n7305 , n7301 );
not ( n7306 , n7302 );
and ( n7307 , n7305 , n7306 );
nor ( n7308 , n7304 , n7307 );
not ( n7309 , n7308 );
xnor ( n7310 , n7298 , n7309 );
not ( n7311 , n7310 );
not ( n7312 , n7311 );
xor ( n7313 , n7269 , n7312 );
buf ( n7314 , n4508 );
buf ( n7315 , n7314 );
buf ( n7316 , n4509 );
buf ( n7317 , n7316 );
not ( n7318 , n7317 );
buf ( n7319 , n4510 );
not ( n7320 , n7319 );
not ( n7321 , n7320 );
or ( n7322 , n7318 , n7321 );
not ( n7323 , n7316 );
buf ( n7324 , n7319 );
nand ( n7325 , n7323 , n7324 );
nand ( n7326 , n7322 , n7325 );
xor ( n7327 , n7315 , n7326 );
buf ( n7328 , n4511 );
buf ( n7329 , n4512 );
xor ( n7330 , n7328 , n7329 );
buf ( n7331 , n4513 );
nand ( n7332 , n7134 , n7331 );
xnor ( n7333 , n7330 , n7332 );
xnor ( n7334 , n7327 , n7333 );
not ( n7335 , n7334 );
not ( n7336 , n7335 );
xnor ( n7337 , n7313 , n7336 );
buf ( n7338 , n4514 );
buf ( n7339 , n7338 );
not ( n7340 , n7339 );
buf ( n7341 , n4515 );
not ( n7342 , n7341 );
not ( n7343 , n7342 );
or ( n7344 , n7340 , n7343 );
not ( n7345 , n7338 );
buf ( n7346 , n7341 );
nand ( n7347 , n7345 , n7346 );
nand ( n7348 , n7344 , n7347 );
buf ( n7349 , n4516 );
buf ( n7350 , n7349 );
and ( n7351 , n7348 , n7350 );
not ( n7352 , n7348 );
not ( n7353 , n7349 );
and ( n7354 , n7352 , n7353 );
nor ( n7355 , n7351 , n7354 );
buf ( n7356 , n7195 );
buf ( n7357 , n4517 );
nand ( n7358 , n7356 , n7357 );
buf ( n7359 , n4518 );
buf ( n7360 , n7359 );
and ( n7361 , n7358 , n7360 );
not ( n7362 , n7358 );
not ( n7363 , n7359 );
and ( n7364 , n7362 , n7363 );
nor ( n7365 , n7361 , n7364 );
xor ( n7366 , n7355 , n7365 );
buf ( n7367 , n4519 );
nand ( n7368 , n6706 , n7367 );
buf ( n7369 , n4520 );
buf ( n7370 , n7369 );
and ( n7371 , n7368 , n7370 );
not ( n7372 , n7368 );
not ( n7373 , n7369 );
and ( n7374 , n7372 , n7373 );
nor ( n7375 , n7371 , n7374 );
xor ( n7376 , n7366 , n7375 );
not ( n7377 , n7376 );
buf ( n7378 , n7377 );
not ( n7379 , n7378 );
buf ( n7380 , n4521 );
buf ( n7381 , n7380 );
not ( n7382 , n7381 );
buf ( n7383 , n4522 );
buf ( n7384 , n7383 );
not ( n7385 , n7384 );
buf ( n7386 , n4523 );
not ( n7387 , n7386 );
not ( n7388 , n7387 );
or ( n7389 , n7385 , n7388 );
not ( n7390 , n7383 );
buf ( n7391 , n7386 );
nand ( n7392 , n7390 , n7391 );
nand ( n7393 , n7389 , n7392 );
buf ( n7394 , n4524 );
not ( n7395 , n7394 );
and ( n7396 , n7393 , n7395 );
not ( n7397 , n7393 );
buf ( n7398 , n7394 );
and ( n7399 , n7397 , n7398 );
nor ( n7400 , n7396 , n7399 );
buf ( n7401 , n6659 );
buf ( n7402 , n4525 );
nand ( n7403 , n7401 , n7402 );
buf ( n7404 , n4526 );
not ( n7405 , n7404 );
and ( n7406 , n7403 , n7405 );
not ( n7407 , n7403 );
buf ( n7408 , n7404 );
and ( n7409 , n7407 , n7408 );
nor ( n7410 , n7406 , n7409 );
xor ( n7411 , n7400 , n7410 );
buf ( n7412 , n6620 );
buf ( n7413 , n7412 );
buf ( n7414 , n4527 );
nand ( n7415 , n7413 , n7414 );
buf ( n7416 , n4528 );
buf ( n7417 , n7416 );
and ( n7418 , n7415 , n7417 );
not ( n7419 , n7415 );
not ( n7420 , n7416 );
and ( n7421 , n7419 , n7420 );
nor ( n7422 , n7418 , n7421 );
xor ( n7423 , n7411 , n7422 );
buf ( n7424 , n7423 );
not ( n7425 , n7424 );
not ( n7426 , n7425 );
or ( n7427 , n7382 , n7426 );
not ( n7428 , n7423 );
not ( n7429 , n7428 );
not ( n7430 , n7380 );
nand ( n7431 , n7429 , n7430 );
nand ( n7432 , n7427 , n7431 );
not ( n7433 , n7432 );
or ( n7434 , n7379 , n7433 );
buf ( n7435 , n7376 );
not ( n7436 , n7435 );
or ( n7437 , n7432 , n7436 );
nand ( n7438 , n7434 , n7437 );
not ( n7439 , n7438 );
nand ( n7440 , n7337 , n7439 );
not ( n7441 , n7440 );
buf ( n7442 , n6760 );
buf ( n7443 , n4529 );
nand ( n7444 , n7442 , n7443 );
buf ( n7445 , n4530 );
not ( n7446 , n7445 );
and ( n7447 , n7444 , n7446 );
not ( n7448 , n7444 );
buf ( n7449 , n7445 );
and ( n7450 , n7448 , n7449 );
nor ( n7451 , n7447 , n7450 );
not ( n7452 , n7451 );
buf ( n7453 , n4531 );
buf ( n7454 , n7453 );
not ( n7455 , n7454 );
buf ( n7456 , n4532 );
not ( n7457 , n7456 );
not ( n7458 , n7457 );
or ( n7459 , n7455 , n7458 );
not ( n7460 , n7453 );
buf ( n7461 , n7456 );
nand ( n7462 , n7460 , n7461 );
nand ( n7463 , n7459 , n7462 );
buf ( n7464 , n4533 );
buf ( n7465 , n7464 );
and ( n7466 , n7463 , n7465 );
not ( n7467 , n7463 );
not ( n7468 , n7464 );
and ( n7469 , n7467 , n7468 );
nor ( n7470 , n7466 , n7469 );
buf ( n7471 , n6606 );
buf ( n7472 , n4534 );
nand ( n7473 , n7471 , n7472 );
buf ( n7474 , n4535 );
xor ( n7475 , n7473 , n7474 );
xor ( n7476 , n7470 , n7475 );
buf ( n7477 , n7132 );
buf ( n7478 , n7477 );
buf ( n7479 , n4536 );
nand ( n7480 , n7478 , n7479 );
buf ( n7481 , n4537 );
buf ( n7482 , n7481 );
and ( n7483 , n7480 , n7482 );
not ( n7484 , n7480 );
not ( n7485 , n7481 );
and ( n7486 , n7484 , n7485 );
nor ( n7487 , n7483 , n7486 );
xnor ( n7488 , n7476 , n7487 );
buf ( n7489 , n7488 );
not ( n7490 , n7489 );
or ( n7491 , n7452 , n7490 );
not ( n7492 , n7451 );
xor ( n7493 , n7470 , n7475 );
not ( n7494 , n7487 );
xnor ( n7495 , n7493 , n7494 );
nand ( n7496 , n7492 , n7495 );
nand ( n7497 , n7491 , n7496 );
not ( n7498 , n7497 );
buf ( n7499 , n4538 );
not ( n7500 , n7499 );
buf ( n7501 , n4539 );
not ( n7502 , n7501 );
buf ( n7503 , n4540 );
buf ( n7504 , n7503 );
nand ( n7505 , n7502 , n7504 );
not ( n7506 , n7503 );
buf ( n7507 , n7501 );
nand ( n7508 , n7506 , n7507 );
and ( n7509 , n7505 , n7508 );
xor ( n7510 , n7500 , n7509 );
buf ( n7511 , n4541 );
buf ( n7512 , n4542 );
buf ( n7513 , n7512 );
xor ( n7514 , n7511 , n7513 );
buf ( n7515 , n6933 );
buf ( n7516 , n7515 );
buf ( n7517 , n4543 );
nand ( n7518 , n7516 , n7517 );
xnor ( n7519 , n7514 , n7518 );
xnor ( n7520 , n7510 , n7519 );
buf ( n7521 , n7520 );
not ( n7522 , n7521 );
and ( n7523 , n7498 , n7522 );
and ( n7524 , n7497 , n7521 );
nor ( n7525 , n7523 , n7524 );
not ( n7526 , n7525 );
not ( n7527 , n7526 );
and ( n7528 , n7441 , n7527 );
and ( n7529 , n7440 , n7526 );
nor ( n7530 , n7528 , n7529 );
buf ( n7531 , n7530 );
not ( n7532 , n7531 );
and ( n7533 , n7267 , n7532 );
not ( n7534 , n7267 );
and ( n7535 , n7534 , n7531 );
nor ( n7536 , n7533 , n7535 );
buf ( n7537 , n4544 );
buf ( n7538 , n7537 );
not ( n7539 , n7538 );
buf ( n7540 , n4545 );
buf ( n7541 , n7540 );
not ( n7542 , n7541 );
buf ( n7543 , n4546 );
not ( n7544 , n7543 );
not ( n7545 , n7544 );
or ( n7546 , n7542 , n7545 );
not ( n7547 , n7540 );
buf ( n7548 , n7543 );
nand ( n7549 , n7547 , n7548 );
nand ( n7550 , n7546 , n7549 );
buf ( n7551 , n4547 );
not ( n7552 , n7551 );
and ( n7553 , n7550 , n7552 );
not ( n7554 , n7550 );
buf ( n7555 , n7551 );
and ( n7556 , n7554 , n7555 );
nor ( n7557 , n7553 , n7556 );
buf ( n7558 , n4548 );
nand ( n7559 , n6851 , n7558 );
buf ( n7560 , n4549 );
buf ( n7561 , n7560 );
and ( n7562 , n7559 , n7561 );
not ( n7563 , n7559 );
not ( n7564 , n7560 );
and ( n7565 , n7563 , n7564 );
nor ( n7566 , n7562 , n7565 );
xor ( n7567 , n7557 , n7566 );
buf ( n7568 , n4550 );
nand ( n7569 , n7413 , n7568 );
buf ( n7570 , n4551 );
not ( n7571 , n7570 );
and ( n7572 , n7569 , n7571 );
not ( n7573 , n7569 );
buf ( n7574 , n7570 );
and ( n7575 , n7573 , n7574 );
nor ( n7576 , n7572 , n7575 );
xnor ( n7577 , n7567 , n7576 );
not ( n7578 , n7577 );
buf ( n7579 , n7578 );
not ( n7580 , n7579 );
not ( n7581 , n7580 );
or ( n7582 , n7539 , n7581 );
buf ( n7583 , n7577 );
not ( n7584 , n7583 );
not ( n7585 , n7537 );
nand ( n7586 , n7584 , n7585 );
nand ( n7587 , n7582 , n7586 );
buf ( n7588 , n4552 );
buf ( n7589 , n7588 );
not ( n7590 , n7589 );
buf ( n7591 , n4553 );
not ( n7592 , n7591 );
not ( n7593 , n7592 );
or ( n7594 , n7590 , n7593 );
not ( n7595 , n7588 );
buf ( n7596 , n7591 );
nand ( n7597 , n7595 , n7596 );
nand ( n7598 , n7594 , n7597 );
buf ( n7599 , n4554 );
not ( n7600 , n7599 );
and ( n7601 , n7598 , n7600 );
not ( n7602 , n7598 );
buf ( n7603 , n7599 );
and ( n7604 , n7602 , n7603 );
nor ( n7605 , n7601 , n7604 );
buf ( n7606 , n4555 );
nand ( n7607 , n7288 , n7606 );
buf ( n7608 , n4556 );
buf ( n7609 , n7608 );
and ( n7610 , n7607 , n7609 );
not ( n7611 , n7607 );
not ( n7612 , n7608 );
and ( n7613 , n7611 , n7612 );
nor ( n7614 , n7610 , n7613 );
xor ( n7615 , n7605 , n7614 );
buf ( n7616 , n6815 );
buf ( n7617 , n7616 );
buf ( n7618 , n4557 );
nand ( n7619 , n7617 , n7618 );
buf ( n7620 , n4558 );
not ( n7621 , n7620 );
and ( n7622 , n7619 , n7621 );
not ( n7623 , n7619 );
buf ( n7624 , n7620 );
and ( n7625 , n7623 , n7624 );
nor ( n7626 , n7622 , n7625 );
xnor ( n7627 , n7615 , n7626 );
buf ( n7628 , n7627 );
buf ( n7629 , n7628 );
xnor ( n7630 , n7587 , n7629 );
buf ( n7631 , n4559 );
buf ( n7632 , n7631 );
not ( n7633 , n7632 );
buf ( n7634 , n4560 );
buf ( n7635 , n7634 );
not ( n7636 , n7635 );
buf ( n7637 , n4561 );
not ( n7638 , n7637 );
not ( n7639 , n7638 );
or ( n7640 , n7636 , n7639 );
not ( n7641 , n7634 );
buf ( n7642 , n7637 );
nand ( n7643 , n7641 , n7642 );
nand ( n7644 , n7640 , n7643 );
buf ( n7645 , n4562 );
not ( n7646 , n7645 );
and ( n7647 , n7644 , n7646 );
not ( n7648 , n7644 );
buf ( n7649 , n7645 );
and ( n7650 , n7648 , n7649 );
nor ( n7651 , n7647 , n7650 );
buf ( n7652 , n4563 );
nand ( n7653 , n7515 , n7652 );
buf ( n7654 , n4564 );
buf ( n7655 , n7654 );
and ( n7656 , n7653 , n7655 );
not ( n7657 , n7653 );
not ( n7658 , n7654 );
and ( n7659 , n7657 , n7658 );
nor ( n7660 , n7656 , n7659 );
xor ( n7661 , n7651 , n7660 );
buf ( n7662 , n4565 );
nand ( n7663 , n6996 , n7662 );
buf ( n7664 , n4566 );
not ( n7665 , n7664 );
and ( n7666 , n7663 , n7665 );
not ( n7667 , n7663 );
buf ( n7668 , n7664 );
and ( n7669 , n7667 , n7668 );
nor ( n7670 , n7666 , n7669 );
xnor ( n7671 , n7661 , n7670 );
buf ( n7672 , n7671 );
not ( n7673 , n7672 );
or ( n7674 , n7633 , n7673 );
or ( n7675 , n7672 , n7632 );
nand ( n7676 , n7674 , n7675 );
not ( n7677 , n7676 );
buf ( n7678 , n4567 );
buf ( n7679 , n7678 );
not ( n7680 , n7679 );
buf ( n7681 , n4568 );
not ( n7682 , n7681 );
not ( n7683 , n7682 );
or ( n7684 , n7680 , n7683 );
not ( n7685 , n7678 );
buf ( n7686 , n7681 );
nand ( n7687 , n7685 , n7686 );
nand ( n7688 , n7684 , n7687 );
buf ( n7689 , n4569 );
not ( n7690 , n7689 );
and ( n7691 , n7688 , n7690 );
not ( n7692 , n7688 );
buf ( n7693 , n7689 );
and ( n7694 , n7692 , n7693 );
nor ( n7695 , n7691 , n7694 );
buf ( n7696 , n4570 );
nand ( n7697 , n7195 , n7696 );
buf ( n7698 , n4571 );
buf ( n7699 , n7698 );
and ( n7700 , n7697 , n7699 );
not ( n7701 , n7697 );
not ( n7702 , n7698 );
and ( n7703 , n7701 , n7702 );
nor ( n7704 , n7700 , n7703 );
xor ( n7705 , n7695 , n7704 );
buf ( n7706 , n4572 );
nand ( n7707 , n7196 , n7706 );
buf ( n7708 , n4573 );
buf ( n7709 , n7708 );
and ( n7710 , n7707 , n7709 );
not ( n7711 , n7707 );
not ( n7712 , n7708 );
and ( n7713 , n7711 , n7712 );
nor ( n7714 , n7710 , n7713 );
xnor ( n7715 , n7705 , n7714 );
not ( n7716 , n7715 );
not ( n7717 , n7716 );
and ( n7718 , n7677 , n7717 );
and ( n7719 , n7676 , n7716 );
nor ( n7720 , n7718 , n7719 );
nand ( n7721 , n7630 , n7720 );
not ( n7722 , n7721 );
buf ( n7723 , n4574 );
nand ( n7724 , n7356 , n7723 );
buf ( n7725 , n4575 );
not ( n7726 , n7725 );
and ( n7727 , n7724 , n7726 );
not ( n7728 , n7724 );
buf ( n7729 , n7725 );
and ( n7730 , n7728 , n7729 );
nor ( n7731 , n7727 , n7730 );
not ( n7732 , n7731 );
buf ( n7733 , n4576 );
buf ( n7734 , n4577 );
buf ( n7735 , n7734 );
not ( n7736 , n7735 );
buf ( n7737 , n4578 );
not ( n7738 , n7737 );
not ( n7739 , n7738 );
or ( n7740 , n7736 , n7739 );
not ( n7741 , n7734 );
buf ( n7742 , n7737 );
nand ( n7743 , n7741 , n7742 );
nand ( n7744 , n7740 , n7743 );
xor ( n7745 , n7733 , n7744 );
buf ( n7746 , n4579 );
buf ( n7747 , n4580 );
not ( n7748 , n7747 );
xor ( n7749 , n7746 , n7748 );
buf ( n7750 , n6606 );
buf ( n7751 , n4581 );
nand ( n7752 , n7750 , n7751 );
xnor ( n7753 , n7749 , n7752 );
xnor ( n7754 , n7745 , n7753 );
buf ( n7755 , n7754 );
not ( n7756 , n7755 );
not ( n7757 , n7756 );
or ( n7758 , n7732 , n7757 );
not ( n7759 , n7731 );
nand ( n7760 , n7759 , n7755 );
nand ( n7761 , n7758 , n7760 );
buf ( n7762 , n4582 );
buf ( n7763 , n7762 );
not ( n7764 , n7763 );
buf ( n7765 , n4583 );
not ( n7766 , n7765 );
not ( n7767 , n7766 );
or ( n7768 , n7764 , n7767 );
not ( n7769 , n7762 );
buf ( n7770 , n7765 );
nand ( n7771 , n7769 , n7770 );
nand ( n7772 , n7768 , n7771 );
buf ( n7773 , n4584 );
not ( n7774 , n7773 );
and ( n7775 , n7772 , n7774 );
not ( n7776 , n7772 );
buf ( n7777 , n7773 );
and ( n7778 , n7776 , n7777 );
nor ( n7779 , n7775 , n7778 );
buf ( n7780 , n4585 );
nand ( n7781 , n7412 , n7780 );
buf ( n7782 , n4586 );
xor ( n7783 , n7781 , n7782 );
xor ( n7784 , n7779 , n7783 );
buf ( n7785 , n7471 );
buf ( n7786 , n4587 );
nand ( n7787 , n7785 , n7786 );
buf ( n7788 , n4588 );
not ( n7789 , n7788 );
and ( n7790 , n7787 , n7789 );
not ( n7791 , n7787 );
buf ( n7792 , n7788 );
and ( n7793 , n7791 , n7792 );
nor ( n7794 , n7790 , n7793 );
xnor ( n7795 , n7784 , n7794 );
buf ( n7796 , n7795 );
xor ( n7797 , n7761 , n7796 );
not ( n7798 , n7797 );
not ( n7799 , n7798 );
and ( n7800 , n7722 , n7799 );
and ( n7801 , n7721 , n7798 );
nor ( n7802 , n7800 , n7801 );
not ( n7803 , n7802 );
buf ( n7804 , n4589 );
buf ( n7805 , n7804 );
buf ( n7806 , n4590 );
buf ( n7807 , n7806 );
not ( n7808 , n7807 );
buf ( n7809 , n4591 );
not ( n7810 , n7809 );
not ( n7811 , n7810 );
or ( n7812 , n7808 , n7811 );
not ( n7813 , n7806 );
buf ( n7814 , n7809 );
nand ( n7815 , n7813 , n7814 );
nand ( n7816 , n7812 , n7815 );
buf ( n7817 , n4592 );
buf ( n7818 , n7817 );
and ( n7819 , n7816 , n7818 );
not ( n7820 , n7816 );
not ( n7821 , n7817 );
and ( n7822 , n7820 , n7821 );
nor ( n7823 , n7819 , n7822 );
buf ( n7824 , n4593 );
nand ( n7825 , n7195 , n7824 );
buf ( n7826 , n4594 );
buf ( n7827 , n7826 );
and ( n7828 , n7825 , n7827 );
not ( n7829 , n7825 );
not ( n7830 , n7826 );
and ( n7831 , n7829 , n7830 );
nor ( n7832 , n7828 , n7831 );
xor ( n7833 , n7823 , n7832 );
buf ( n7834 , n4595 );
nand ( n7835 , n7126 , n7834 );
buf ( n7836 , n4596 );
buf ( n7837 , n7836 );
and ( n7838 , n7835 , n7837 );
not ( n7839 , n7835 );
not ( n7840 , n7836 );
and ( n7841 , n7839 , n7840 );
nor ( n7842 , n7838 , n7841 );
not ( n7843 , n7842 );
xnor ( n7844 , n7833 , n7843 );
xor ( n7845 , n7805 , n7844 );
buf ( n7846 , n4597 );
buf ( n7847 , n4598 );
buf ( n7848 , n7847 );
not ( n7849 , n7848 );
buf ( n7850 , n4599 );
not ( n7851 , n7850 );
not ( n7852 , n7851 );
or ( n7853 , n7849 , n7852 );
not ( n7854 , n7847 );
buf ( n7855 , n7850 );
nand ( n7856 , n7854 , n7855 );
nand ( n7857 , n7853 , n7856 );
xor ( n7858 , n7846 , n7857 );
buf ( n7859 , n4600 );
nand ( n7860 , n7195 , n7859 );
not ( n7861 , n7860 );
buf ( n7862 , n4601 );
not ( n7863 , n7862 );
and ( n7864 , n7861 , n7863 );
buf ( n7865 , n7125 );
nand ( n7866 , n7865 , n7859 );
and ( n7867 , n7866 , n7862 );
nor ( n7868 , n7864 , n7867 );
not ( n7869 , n7868 );
buf ( n7870 , n4602 );
nand ( n7871 , n6660 , n7870 );
buf ( n7872 , n4603 );
not ( n7873 , n7872 );
and ( n7874 , n7871 , n7873 );
not ( n7875 , n7871 );
buf ( n7876 , n7872 );
and ( n7877 , n7875 , n7876 );
nor ( n7878 , n7874 , n7877 );
not ( n7879 , n7878 );
or ( n7880 , n7869 , n7879 );
not ( n7881 , n7878 );
not ( n7882 , n7868 );
nand ( n7883 , n7881 , n7882 );
nand ( n7884 , n7880 , n7883 );
xnor ( n7885 , n7858 , n7884 );
buf ( n7886 , n7885 );
xnor ( n7887 , n7845 , n7886 );
buf ( n7888 , n4604 );
buf ( n7889 , n7888 );
not ( n7890 , n7889 );
buf ( n7891 , n4605 );
buf ( n7892 , n7891 );
not ( n7893 , n7892 );
buf ( n7894 , n4606 );
not ( n7895 , n7894 );
not ( n7896 , n7895 );
or ( n7897 , n7893 , n7896 );
not ( n7898 , n7891 );
buf ( n7899 , n7894 );
nand ( n7900 , n7898 , n7899 );
nand ( n7901 , n7897 , n7900 );
buf ( n7902 , n4607 );
buf ( n7903 , n7902 );
and ( n7904 , n7901 , n7903 );
not ( n7905 , n7901 );
not ( n7906 , n7902 );
and ( n7907 , n7905 , n7906 );
nor ( n7908 , n7904 , n7907 );
buf ( n7909 , n6606 );
buf ( n7910 , n4608 );
nand ( n7911 , n7909 , n7910 );
buf ( n7912 , n4609 );
buf ( n7913 , n7912 );
and ( n7914 , n7911 , n7913 );
not ( n7915 , n7911 );
not ( n7916 , n7912 );
and ( n7917 , n7915 , n7916 );
nor ( n7918 , n7914 , n7917 );
xor ( n7919 , n7908 , n7918 );
buf ( n7920 , n6862 );
buf ( n7921 , n7920 );
buf ( n7922 , n4610 );
nand ( n7923 , n7921 , n7922 );
buf ( n7924 , n4611 );
not ( n7925 , n7924 );
and ( n7926 , n7923 , n7925 );
not ( n7927 , n7923 );
buf ( n7928 , n7924 );
and ( n7929 , n7927 , n7928 );
nor ( n7930 , n7926 , n7929 );
xnor ( n7931 , n7919 , n7930 );
buf ( n7932 , n7931 );
not ( n7933 , n7932 );
not ( n7934 , n7933 );
or ( n7935 , n7890 , n7934 );
or ( n7936 , n7933 , n7889 );
nand ( n7937 , n7935 , n7936 );
buf ( n7938 , n4612 );
not ( n7939 , n7938 );
buf ( n7940 , n4613 );
buf ( n7941 , n7940 );
not ( n7942 , n7941 );
buf ( n7943 , n4614 );
not ( n7944 , n7943 );
not ( n7945 , n7944 );
or ( n7946 , n7942 , n7945 );
not ( n7947 , n7940 );
buf ( n7948 , n7943 );
nand ( n7949 , n7947 , n7948 );
nand ( n7950 , n7946 , n7949 );
not ( n7951 , n7950 );
xor ( n7952 , n7939 , n7951 );
buf ( n7953 , n4615 );
not ( n7954 , n7953 );
buf ( n7955 , n6815 );
buf ( n7956 , n4616 );
nand ( n7957 , n7955 , n7956 );
buf ( n7958 , n4617 );
buf ( n7959 , n7958 );
and ( n7960 , n7957 , n7959 );
not ( n7961 , n7957 );
not ( n7962 , n7958 );
and ( n7963 , n7961 , n7962 );
nor ( n7964 , n7960 , n7963 );
not ( n7965 , n7964 );
or ( n7966 , n7954 , n7965 );
or ( n7967 , n7964 , n7953 );
nand ( n7968 , n7966 , n7967 );
xnor ( n7969 , n7952 , n7968 );
buf ( n7970 , n7969 );
and ( n7971 , n7937 , n7970 );
not ( n7972 , n7937 );
buf ( n7973 , n7938 );
xor ( n7974 , n7973 , n7950 );
not ( n7975 , n7968 );
xnor ( n7976 , n7974 , n7975 );
buf ( n7977 , n7976 );
and ( n7978 , n7972 , n7977 );
nor ( n7979 , n7971 , n7978 );
nand ( n7980 , n7887 , n7979 );
buf ( n7981 , n7125 );
buf ( n7982 , n4618 );
nand ( n7983 , n7981 , n7982 );
buf ( n7984 , n4619 );
buf ( n7985 , n7984 );
and ( n7986 , n7983 , n7985 );
not ( n7987 , n7983 );
not ( n7988 , n7984 );
and ( n7989 , n7987 , n7988 );
nor ( n7990 , n7986 , n7989 );
buf ( n7991 , n7990 );
not ( n7992 , n7991 );
buf ( n7993 , n4620 );
buf ( n7994 , n7993 );
not ( n7995 , n7994 );
buf ( n7996 , n4621 );
not ( n7997 , n7996 );
not ( n7998 , n7997 );
or ( n7999 , n7995 , n7998 );
not ( n8000 , n7993 );
buf ( n8001 , n7996 );
nand ( n8002 , n8000 , n8001 );
nand ( n8003 , n7999 , n8002 );
buf ( n8004 , n4622 );
not ( n8005 , n8004 );
and ( n8006 , n8003 , n8005 );
not ( n8007 , n8003 );
buf ( n8008 , n8004 );
and ( n8009 , n8007 , n8008 );
nor ( n8010 , n8006 , n8009 );
buf ( n8011 , n4623 );
nand ( n8012 , n7043 , n8011 );
buf ( n8013 , n4624 );
xor ( n8014 , n8012 , n8013 );
xor ( n8015 , n8010 , n8014 );
buf ( n8016 , n4625 );
nand ( n8017 , n6996 , n8016 );
buf ( n8018 , n4626 );
not ( n8019 , n8018 );
and ( n8020 , n8017 , n8019 );
not ( n8021 , n8017 );
buf ( n8022 , n8018 );
and ( n8023 , n8021 , n8022 );
nor ( n8024 , n8020 , n8023 );
xnor ( n8025 , n8015 , n8024 );
buf ( n8026 , n8025 );
not ( n8027 , n8026 );
not ( n8028 , n8027 );
or ( n8029 , n7992 , n8028 );
or ( n8030 , n8027 , n7991 );
nand ( n8031 , n8029 , n8030 );
not ( n8032 , n8031 );
buf ( n8033 , n4627 );
buf ( n8034 , n8033 );
not ( n8035 , n8034 );
buf ( n8036 , n4628 );
not ( n8037 , n8036 );
not ( n8038 , n8037 );
or ( n8039 , n8035 , n8038 );
not ( n8040 , n8033 );
buf ( n8041 , n8036 );
nand ( n8042 , n8040 , n8041 );
nand ( n8043 , n8039 , n8042 );
not ( n8044 , n8043 );
not ( n8045 , n8044 );
buf ( n8046 , n4629 );
buf ( n8047 , n4630 );
buf ( n8048 , n8047 );
not ( n8049 , n8048 );
buf ( n8050 , n4631 );
nand ( n8051 , n7750 , n8050 );
not ( n8052 , n8051 );
or ( n8053 , n8049 , n8052 );
not ( n8054 , n8047 );
nand ( n8055 , n7471 , n8054 , n8050 );
nand ( n8056 , n8053 , n8055 );
xor ( n8057 , n8046 , n8056 );
buf ( n8058 , n4632 );
nand ( n8059 , n6706 , n8058 );
buf ( n8060 , n4633 );
not ( n8061 , n8060 );
and ( n8062 , n8059 , n8061 );
not ( n8063 , n8059 );
buf ( n8064 , n8060 );
and ( n8065 , n8063 , n8064 );
nor ( n8066 , n8062 , n8065 );
xnor ( n8067 , n8057 , n8066 );
not ( n8068 , n8067 );
not ( n8069 , n8068 );
or ( n8070 , n8045 , n8069 );
nand ( n8071 , n8067 , n8043 );
nand ( n8072 , n8070 , n8071 );
not ( n8073 , n8072 );
buf ( n8074 , n8073 );
not ( n8075 , n8074 );
or ( n8076 , n8032 , n8075 );
or ( n8077 , n8074 , n8031 );
nand ( n8078 , n8076 , n8077 );
not ( n8079 , n8078 );
and ( n8080 , n7980 , n8079 );
not ( n8081 , n7980 );
and ( n8082 , n8081 , n8078 );
nor ( n8083 , n8080 , n8082 );
not ( n8084 , n8083 );
or ( n8085 , n7803 , n8084 );
or ( n8086 , n8083 , n7802 );
nand ( n8087 , n8085 , n8086 );
xnor ( n8088 , n7536 , n8087 );
not ( n8089 , n8088 );
or ( n8090 , n6886 , n8089 );
not ( n8091 , n6885 );
xor ( n8092 , n7530 , n7267 );
xnor ( n8093 , n8092 , n8087 );
nand ( n8094 , n8091 , n8093 );
nand ( n8095 , n8090 , n8094 );
buf ( n8096 , n4634 );
nand ( n8097 , n7356 , n8096 );
buf ( n8098 , n4635 );
not ( n8099 , n8098 );
and ( n8100 , n8097 , n8099 );
not ( n8101 , n8097 );
buf ( n8102 , n8098 );
and ( n8103 , n8101 , n8102 );
nor ( n8104 , n8100 , n8103 );
not ( n8105 , n8104 );
buf ( n8106 , n4636 );
buf ( n8107 , n8106 );
not ( n8108 , n8107 );
buf ( n8109 , n4637 );
not ( n8110 , n8109 );
not ( n8111 , n8110 );
or ( n8112 , n8108 , n8111 );
not ( n8113 , n8106 );
buf ( n8114 , n8109 );
nand ( n8115 , n8113 , n8114 );
nand ( n8116 , n8112 , n8115 );
buf ( n8117 , n4638 );
buf ( n8118 , n8117 );
and ( n8119 , n8116 , n8118 );
not ( n8120 , n8116 );
not ( n8121 , n8117 );
and ( n8122 , n8120 , n8121 );
nor ( n8123 , n8119 , n8122 );
buf ( n8124 , n4639 );
nand ( n8125 , n7471 , n8124 );
buf ( n8126 , n4640 );
buf ( n8127 , n8126 );
and ( n8128 , n8125 , n8127 );
not ( n8129 , n8125 );
not ( n8130 , n8126 );
and ( n8131 , n8129 , n8130 );
nor ( n8132 , n8128 , n8131 );
xor ( n8133 , n8123 , n8132 );
buf ( n8134 , n6659 );
buf ( n8135 , n8134 );
buf ( n8136 , n4641 );
nand ( n8137 , n8135 , n8136 );
buf ( n8138 , n4642 );
not ( n8139 , n8138 );
and ( n8140 , n8137 , n8139 );
not ( n8141 , n8137 );
buf ( n8142 , n8138 );
and ( n8143 , n8141 , n8142 );
nor ( n8144 , n8140 , n8143 );
xor ( n8145 , n8133 , n8144 );
not ( n8146 , n8145 );
or ( n8147 , n8105 , n8146 );
not ( n8148 , n8104 );
xor ( n8149 , n8123 , n8132 );
xnor ( n8150 , n8149 , n8144 );
nand ( n8151 , n8148 , n8150 );
nand ( n8152 , n8147 , n8151 );
not ( n8153 , n8152 );
buf ( n8154 , n4643 );
buf ( n8155 , n8154 );
not ( n8156 , n8155 );
buf ( n8157 , n4644 );
not ( n8158 , n8157 );
not ( n8159 , n8158 );
or ( n8160 , n8156 , n8159 );
not ( n8161 , n8154 );
buf ( n8162 , n8157 );
nand ( n8163 , n8161 , n8162 );
nand ( n8164 , n8160 , n8163 );
not ( n8165 , n8164 );
buf ( n8166 , n4645 );
buf ( n8167 , n4646 );
nand ( n8168 , n6760 , n8167 );
buf ( n8169 , n4647 );
buf ( n8170 , n8169 );
and ( n8171 , n8168 , n8170 );
not ( n8172 , n8168 );
not ( n8173 , n8169 );
and ( n8174 , n8172 , n8173 );
nor ( n8175 , n8171 , n8174 );
xor ( n8176 , n8166 , n8175 );
buf ( n8177 , n4648 );
nand ( n8178 , n6934 , n8177 );
buf ( n8179 , n4649 );
buf ( n8180 , n8179 );
and ( n8181 , n8178 , n8180 );
not ( n8182 , n8178 );
not ( n8183 , n8179 );
and ( n8184 , n8182 , n8183 );
nor ( n8185 , n8181 , n8184 );
xnor ( n8186 , n8176 , n8185 );
not ( n8187 , n8186 );
or ( n8188 , n8165 , n8187 );
not ( n8189 , n8186 );
not ( n8190 , n8164 );
nand ( n8191 , n8189 , n8190 );
nand ( n8192 , n8188 , n8191 );
not ( n8193 , n8192 );
not ( n8194 , n8193 );
or ( n8195 , n8153 , n8194 );
or ( n8196 , n8193 , n8152 );
nand ( n8197 , n8195 , n8196 );
buf ( n8198 , n4650 );
not ( n8199 , n8198 );
buf ( n8200 , n4651 );
buf ( n8201 , n8200 );
not ( n8202 , n8201 );
buf ( n8203 , n4652 );
not ( n8204 , n8203 );
not ( n8205 , n8204 );
or ( n8206 , n8202 , n8205 );
not ( n8207 , n8200 );
buf ( n8208 , n8203 );
nand ( n8209 , n8207 , n8208 );
nand ( n8210 , n8206 , n8209 );
not ( n8211 , n8210 );
xor ( n8212 , n8199 , n8211 );
buf ( n8213 , n4653 );
nand ( n8214 , n7412 , n8213 );
buf ( n8215 , n4654 );
buf ( n8216 , n8215 );
and ( n8217 , n8214 , n8216 );
not ( n8218 , n8214 );
not ( n8219 , n8215 );
and ( n8220 , n8218 , n8219 );
nor ( n8221 , n8217 , n8220 );
not ( n8222 , n8221 );
buf ( n8223 , n6659 );
buf ( n8224 , n4655 );
nand ( n8225 , n8223 , n8224 );
buf ( n8226 , n4656 );
not ( n8227 , n8226 );
and ( n8228 , n8225 , n8227 );
not ( n8229 , n8225 );
buf ( n8230 , n8226 );
and ( n8231 , n8229 , n8230 );
nor ( n8232 , n8228 , n8231 );
not ( n8233 , n8232 );
or ( n8234 , n8222 , n8233 );
or ( n8235 , n8221 , n8232 );
nand ( n8236 , n8234 , n8235 );
xnor ( n8237 , n8212 , n8236 );
buf ( n8238 , n8237 );
not ( n8239 , n8238 );
buf ( n8240 , n4657 );
buf ( n8241 , n8240 );
not ( n8242 , n8241 );
buf ( n8243 , n4658 );
buf ( n8244 , n8243 );
not ( n8245 , n8244 );
not ( n8246 , n6887 );
not ( n8247 , n8246 );
or ( n8248 , n8245 , n8247 );
not ( n8249 , n8243 );
nand ( n8250 , n8249 , n6888 );
nand ( n8251 , n8248 , n8250 );
buf ( n8252 , n4659 );
buf ( n8253 , n8252 );
and ( n8254 , n8251 , n8253 );
not ( n8255 , n8251 );
not ( n8256 , n8252 );
and ( n8257 , n8255 , n8256 );
nor ( n8258 , n8254 , n8257 );
buf ( n8259 , n4660 );
nand ( n8260 , n7909 , n8259 );
buf ( n8261 , n4661 );
buf ( n8262 , n8261 );
and ( n8263 , n8260 , n8262 );
not ( n8264 , n8260 );
not ( n8265 , n8261 );
and ( n8266 , n8264 , n8265 );
nor ( n8267 , n8263 , n8266 );
xor ( n8268 , n8258 , n8267 );
buf ( n8269 , n7909 );
buf ( n8270 , n4662 );
nand ( n8271 , n8269 , n8270 );
buf ( n8272 , n4663 );
not ( n8273 , n8272 );
and ( n8274 , n8271 , n8273 );
not ( n8275 , n8271 );
buf ( n8276 , n8272 );
and ( n8277 , n8275 , n8276 );
nor ( n8278 , n8274 , n8277 );
xnor ( n8279 , n8268 , n8278 );
not ( n8280 , n8279 );
not ( n8281 , n8280 );
or ( n8282 , n8242 , n8281 );
or ( n8283 , n8280 , n8241 );
nand ( n8284 , n8282 , n8283 );
not ( n8285 , n8284 );
and ( n8286 , n8239 , n8285 );
not ( n8287 , n8237 );
not ( n8288 , n8287 );
and ( n8289 , n8288 , n8284 );
nor ( n8290 , n8286 , n8289 );
nand ( n8291 , n8197 , n8290 );
not ( n8292 , n8291 );
buf ( n8293 , n6828 );
not ( n8294 , n8293 );
buf ( n8295 , n4664 );
buf ( n8296 , n8295 );
not ( n8297 , n8296 );
buf ( n8298 , n4665 );
not ( n8299 , n8298 );
buf ( n8300 , n4666 );
buf ( n8301 , n8300 );
not ( n8302 , n8301 );
buf ( n8303 , n4667 );
not ( n8304 , n8303 );
not ( n8305 , n8304 );
or ( n8306 , n8302 , n8305 );
not ( n8307 , n8300 );
buf ( n8308 , n8303 );
nand ( n8309 , n8307 , n8308 );
nand ( n8310 , n8306 , n8309 );
xor ( n8311 , n8299 , n8310 );
buf ( n8312 , n4668 );
not ( n8313 , n8312 );
not ( n8314 , n8313 );
buf ( n8315 , n4669 );
nand ( n8316 , n7401 , n8315 );
buf ( n8317 , n4670 );
not ( n8318 , n8317 );
and ( n8319 , n8316 , n8318 );
not ( n8320 , n8316 );
buf ( n8321 , n8317 );
and ( n8322 , n8320 , n8321 );
nor ( n8323 , n8319 , n8322 );
not ( n8324 , n8323 );
or ( n8325 , n8314 , n8324 );
or ( n8326 , n8323 , n8313 );
nand ( n8327 , n8325 , n8326 );
xnor ( n8328 , n8311 , n8327 );
not ( n8329 , n8328 );
not ( n8330 , n8329 );
or ( n8331 , n8297 , n8330 );
or ( n8332 , n8329 , n8296 );
nand ( n8333 , n8331 , n8332 );
not ( n8334 , n8333 );
or ( n8335 , n8294 , n8334 );
or ( n8336 , n8333 , n8293 );
nand ( n8337 , n8335 , n8336 );
not ( n8338 , n8337 );
and ( n8339 , n8292 , n8338 );
and ( n8340 , n8291 , n8337 );
nor ( n8341 , n8339 , n8340 );
not ( n8342 , n8341 );
buf ( n8343 , n6620 );
buf ( n8344 , n8343 );
buf ( n8345 , n4671 );
nand ( n8346 , n8344 , n8345 );
buf ( n8347 , n4672 );
buf ( n8348 , n8347 );
and ( n8349 , n8346 , n8348 );
not ( n8350 , n8346 );
not ( n8351 , n8347 );
and ( n8352 , n8350 , n8351 );
nor ( n8353 , n8349 , n8352 );
buf ( n8354 , n8353 );
not ( n8355 , n8354 );
buf ( n8356 , n4673 );
buf ( n8357 , n4674 );
not ( n8358 , n8357 );
buf ( n8359 , n4675 );
buf ( n8360 , n8359 );
and ( n8361 , n8358 , n8360 );
not ( n8362 , n8358 );
not ( n8363 , n8359 );
and ( n8364 , n8362 , n8363 );
nor ( n8365 , n8361 , n8364 );
xor ( n8366 , n8356 , n8365 );
buf ( n8367 , n4676 );
not ( n8368 , n8367 );
buf ( n8369 , n4677 );
nand ( n8370 , n6905 , n8369 );
buf ( n8371 , n4678 );
buf ( n8372 , n8371 );
and ( n8373 , n8370 , n8372 );
not ( n8374 , n8370 );
not ( n8375 , n8371 );
and ( n8376 , n8374 , n8375 );
nor ( n8377 , n8373 , n8376 );
not ( n8378 , n8377 );
or ( n8379 , n8368 , n8378 );
or ( n8380 , n8377 , n8367 );
nand ( n8381 , n8379 , n8380 );
xnor ( n8382 , n8366 , n8381 );
not ( n8383 , n8382 );
or ( n8384 , n8355 , n8383 );
or ( n8385 , n8382 , n8354 );
nand ( n8386 , n8384 , n8385 );
buf ( n8387 , n7125 );
buf ( n8388 , n4679 );
nand ( n8389 , n8387 , n8388 );
buf ( n8390 , n4680 );
buf ( n8391 , n8390 );
and ( n8392 , n8389 , n8391 );
not ( n8393 , n8389 );
not ( n8394 , n8390 );
and ( n8395 , n8393 , n8394 );
nor ( n8396 , n8392 , n8395 );
not ( n8397 , n8396 );
buf ( n8398 , n4681 );
nand ( n8399 , n7299 , n8398 );
buf ( n8400 , n4682 );
not ( n8401 , n8400 );
and ( n8402 , n8399 , n8401 );
not ( n8403 , n8399 );
buf ( n8404 , n8400 );
and ( n8405 , n8403 , n8404 );
nor ( n8406 , n8402 , n8405 );
not ( n8407 , n8406 );
or ( n8408 , n8397 , n8407 );
or ( n8409 , n8396 , n8406 );
nand ( n8410 , n8408 , n8409 );
buf ( n8411 , n4683 );
buf ( n8412 , n8411 );
not ( n8413 , n8412 );
buf ( n8414 , n4684 );
not ( n8415 , n8414 );
not ( n8416 , n8415 );
or ( n8417 , n8413 , n8416 );
not ( n8418 , n8411 );
buf ( n8419 , n8414 );
nand ( n8420 , n8418 , n8419 );
nand ( n8421 , n8417 , n8420 );
buf ( n8422 , n4685 );
not ( n8423 , n8422 );
and ( n8424 , n8421 , n8423 );
not ( n8425 , n8421 );
buf ( n8426 , n8422 );
and ( n8427 , n8425 , n8426 );
nor ( n8428 , n8424 , n8427 );
not ( n8429 , n8428 );
and ( n8430 , n8410 , n8429 );
not ( n8431 , n8410 );
and ( n8432 , n8431 , n8428 );
nor ( n8433 , n8430 , n8432 );
buf ( n8434 , n8433 );
and ( n8435 , n8386 , n8434 );
not ( n8436 , n8386 );
buf ( n8437 , n8396 );
xor ( n8438 , n8428 , n8437 );
buf ( n8439 , n8406 );
xnor ( n8440 , n8438 , n8439 );
buf ( n8441 , n8440 );
and ( n8442 , n8436 , n8441 );
nor ( n8443 , n8435 , n8442 );
buf ( n8444 , n4686 );
not ( n8445 , n8444 );
buf ( n8446 , n4687 );
buf ( n8447 , n8446 );
not ( n8448 , n8447 );
buf ( n8449 , n4688 );
not ( n8450 , n8449 );
not ( n8451 , n8450 );
or ( n8452 , n8448 , n8451 );
not ( n8453 , n8446 );
buf ( n8454 , n8449 );
nand ( n8455 , n8453 , n8454 );
nand ( n8456 , n8452 , n8455 );
buf ( n8457 , n4689 );
buf ( n8458 , n8457 );
and ( n8459 , n8456 , n8458 );
not ( n8460 , n8456 );
not ( n8461 , n8457 );
and ( n8462 , n8460 , n8461 );
nor ( n8463 , n8459 , n8462 );
buf ( n8464 , n4690 );
nand ( n8465 , n7909 , n8464 );
buf ( n8466 , n4691 );
buf ( n8467 , n8466 );
and ( n8468 , n8465 , n8467 );
not ( n8469 , n8465 );
not ( n8470 , n8466 );
and ( n8471 , n8469 , n8470 );
nor ( n8472 , n8468 , n8471 );
xor ( n8473 , n8463 , n8472 );
buf ( n8474 , n4692 );
nand ( n8475 , n7750 , n8474 );
buf ( n8476 , n4693 );
not ( n8477 , n8476 );
and ( n8478 , n8475 , n8477 );
not ( n8479 , n8475 );
buf ( n8480 , n8476 );
and ( n8481 , n8479 , n8480 );
nor ( n8482 , n8478 , n8481 );
xor ( n8483 , n8473 , n8482 );
not ( n8484 , n8483 );
or ( n8485 , n8445 , n8484 );
not ( n8486 , n8444 );
xor ( n8487 , n8463 , n8472 );
xnor ( n8488 , n8487 , n8482 );
nand ( n8489 , n8486 , n8488 );
nand ( n8490 , n8485 , n8489 );
buf ( n8491 , n4694 );
buf ( n8492 , n8491 );
not ( n8493 , n8492 );
buf ( n8494 , n4695 );
not ( n8495 , n8494 );
not ( n8496 , n8495 );
or ( n8497 , n8493 , n8496 );
not ( n8498 , n8491 );
buf ( n8499 , n8494 );
nand ( n8500 , n8498 , n8499 );
nand ( n8501 , n8497 , n8500 );
buf ( n8502 , n4696 );
buf ( n8503 , n8502 );
and ( n8504 , n8501 , n8503 );
not ( n8505 , n8501 );
not ( n8506 , n8502 );
and ( n8507 , n8505 , n8506 );
nor ( n8508 , n8504 , n8507 );
buf ( n8509 , n4697 );
nand ( n8510 , n7955 , n8509 );
buf ( n8511 , n4698 );
not ( n8512 , n8511 );
and ( n8513 , n8510 , n8512 );
not ( n8514 , n8510 );
buf ( n8515 , n8511 );
and ( n8516 , n8514 , n8515 );
nor ( n8517 , n8513 , n8516 );
xor ( n8518 , n8508 , n8517 );
buf ( n8519 , n8343 );
buf ( n8520 , n8519 );
buf ( n8521 , n4699 );
nand ( n8522 , n8520 , n8521 );
buf ( n8523 , n4700 );
not ( n8524 , n8523 );
and ( n8525 , n8522 , n8524 );
not ( n8526 , n8522 );
buf ( n8527 , n8523 );
and ( n8528 , n8526 , n8527 );
nor ( n8529 , n8525 , n8528 );
xnor ( n8530 , n8518 , n8529 );
not ( n8531 , n8530 );
buf ( n8532 , n8531 );
not ( n8533 , n8532 );
and ( n8534 , n8490 , n8533 );
not ( n8535 , n8490 );
not ( n8536 , n8531 );
not ( n8537 , n8536 );
and ( n8538 , n8535 , n8537 );
nor ( n8539 , n8534 , n8538 );
nand ( n8540 , n8443 , n8539 );
buf ( n8541 , n4701 );
buf ( n8542 , n8541 );
buf ( n8543 , n4702 );
buf ( n8544 , n8543 );
not ( n8545 , n8544 );
buf ( n8546 , n4703 );
not ( n8547 , n8546 );
not ( n8548 , n8547 );
or ( n8549 , n8545 , n8548 );
not ( n8550 , n8543 );
buf ( n8551 , n8546 );
nand ( n8552 , n8550 , n8551 );
nand ( n8553 , n8549 , n8552 );
buf ( n8554 , n4704 );
not ( n8555 , n8554 );
and ( n8556 , n8553 , n8555 );
not ( n8557 , n8553 );
buf ( n8558 , n8554 );
and ( n8559 , n8557 , n8558 );
nor ( n8560 , n8556 , n8559 );
buf ( n8561 , n4705 );
nand ( n8562 , n7471 , n8561 );
buf ( n8563 , n4706 );
not ( n8564 , n8563 );
and ( n8565 , n8562 , n8564 );
not ( n8566 , n8562 );
buf ( n8567 , n8563 );
and ( n8568 , n8566 , n8567 );
nor ( n8569 , n8565 , n8568 );
xor ( n8570 , n8560 , n8569 );
buf ( n8571 , n4707 );
nand ( n8572 , n7477 , n8571 );
buf ( n8573 , n4708 );
buf ( n8574 , n8573 );
and ( n8575 , n8572 , n8574 );
not ( n8576 , n8572 );
not ( n8577 , n8573 );
and ( n8578 , n8576 , n8577 );
nor ( n8579 , n8575 , n8578 );
xor ( n8580 , n8570 , n8579 );
not ( n8581 , n8580 );
xor ( n8582 , n8542 , n8581 );
not ( n8583 , n8582 );
buf ( n8584 , n4709 );
not ( n8585 , n8584 );
buf ( n8586 , n4710 );
buf ( n8587 , n8586 );
and ( n8588 , n8585 , n8587 );
not ( n8589 , n8585 );
not ( n8590 , n8586 );
and ( n8591 , n8589 , n8590 );
nor ( n8592 , n8588 , n8591 );
not ( n8593 , n8592 );
buf ( n8594 , n4711 );
buf ( n8595 , n4712 );
not ( n8596 , n8595 );
xor ( n8597 , n8594 , n8596 );
buf ( n8598 , n4713 );
nand ( n8599 , n7442 , n8598 );
buf ( n8600 , n4714 );
not ( n8601 , n8600 );
and ( n8602 , n8599 , n8601 );
not ( n8603 , n8599 );
buf ( n8604 , n8600 );
and ( n8605 , n8603 , n8604 );
nor ( n8606 , n8602 , n8605 );
xnor ( n8607 , n8597 , n8606 );
not ( n8608 , n8607 );
or ( n8609 , n8593 , n8608 );
or ( n8610 , n8607 , n8592 );
nand ( n8611 , n8609 , n8610 );
buf ( n8612 , n8611 );
not ( n8613 , n8612 );
or ( n8614 , n8583 , n8613 );
or ( n8615 , n8612 , n8582 );
nand ( n8616 , n8614 , n8615 );
not ( n8617 , n8616 );
and ( n8618 , n8540 , n8617 );
not ( n8619 , n8540 );
and ( n8620 , n8619 , n8616 );
nor ( n8621 , n8618 , n8620 );
not ( n8622 , n8621 );
or ( n8623 , n8342 , n8622 );
or ( n8624 , n8621 , n8341 );
nand ( n8625 , n8623 , n8624 );
buf ( n8626 , n4715 );
buf ( n8627 , n8626 );
buf ( n8628 , n4716 );
buf ( n8629 , n8628 );
not ( n8630 , n8629 );
buf ( n8631 , n4717 );
not ( n8632 , n8631 );
not ( n8633 , n8632 );
or ( n8634 , n8630 , n8633 );
not ( n8635 , n8628 );
buf ( n8636 , n8631 );
nand ( n8637 , n8635 , n8636 );
nand ( n8638 , n8634 , n8637 );
buf ( n8639 , n4718 );
not ( n8640 , n8639 );
and ( n8641 , n8638 , n8640 );
not ( n8642 , n8638 );
buf ( n8643 , n8639 );
and ( n8644 , n8642 , n8643 );
nor ( n8645 , n8641 , n8644 );
buf ( n8646 , n4719 );
nand ( n8647 , n7750 , n8646 );
buf ( n8648 , n4720 );
buf ( n8649 , n8648 );
and ( n8650 , n8647 , n8649 );
not ( n8651 , n8647 );
not ( n8652 , n8648 );
and ( n8653 , n8651 , n8652 );
nor ( n8654 , n8650 , n8653 );
xor ( n8655 , n8645 , n8654 );
buf ( n8656 , n4721 );
nand ( n8657 , n7196 , n8656 );
buf ( n8658 , n4722 );
buf ( n8659 , n8658 );
and ( n8660 , n8657 , n8659 );
not ( n8661 , n8657 );
not ( n8662 , n8658 );
and ( n8663 , n8661 , n8662 );
nor ( n8664 , n8660 , n8663 );
xor ( n8665 , n8655 , n8664 );
not ( n8666 , n8665 );
xor ( n8667 , n8627 , n8666 );
buf ( n8668 , n4723 );
buf ( n8669 , n8668 );
not ( n8670 , n8669 );
buf ( n8671 , n4724 );
not ( n8672 , n8671 );
not ( n8673 , n8672 );
or ( n8674 , n8670 , n8673 );
not ( n8675 , n8668 );
buf ( n8676 , n8671 );
nand ( n8677 , n8675 , n8676 );
nand ( n8678 , n8674 , n8677 );
not ( n8679 , n8678 );
buf ( n8680 , n4725 );
buf ( n8681 , n8680 );
buf ( n8682 , n4726 );
nand ( n8683 , n8387 , n8682 );
buf ( n8684 , n4727 );
buf ( n8685 , n8684 );
and ( n8686 , n8683 , n8685 );
not ( n8687 , n8683 );
not ( n8688 , n8684 );
and ( n8689 , n8687 , n8688 );
nor ( n8690 , n8686 , n8689 );
xor ( n8691 , n8681 , n8690 );
buf ( n8692 , n4728 );
nand ( n8693 , n6945 , n8692 );
buf ( n8694 , n4729 );
not ( n8695 , n8694 );
and ( n8696 , n8693 , n8695 );
not ( n8697 , n8693 );
buf ( n8698 , n8694 );
and ( n8699 , n8697 , n8698 );
nor ( n8700 , n8696 , n8699 );
xnor ( n8701 , n8691 , n8700 );
not ( n8702 , n8701 );
not ( n8703 , n8702 );
or ( n8704 , n8679 , n8703 );
not ( n8705 , n8678 );
nand ( n8706 , n8705 , n8701 );
nand ( n8707 , n8704 , n8706 );
not ( n8708 , n8707 );
xnor ( n8709 , n8667 , n8708 );
not ( n8710 , n8709 );
buf ( n8711 , n4730 );
nand ( n8712 , n7955 , n8711 );
buf ( n8713 , n4731 );
buf ( n8714 , n8713 );
and ( n8715 , n8712 , n8714 );
not ( n8716 , n8712 );
not ( n8717 , n8713 );
and ( n8718 , n8716 , n8717 );
nor ( n8719 , n8715 , n8718 );
not ( n8720 , n8719 );
not ( n8721 , n8720 );
buf ( n8722 , n4732 );
buf ( n8723 , n8722 );
not ( n8724 , n8723 );
buf ( n8725 , n4733 );
not ( n8726 , n8725 );
not ( n8727 , n8726 );
or ( n8728 , n8724 , n8727 );
not ( n8729 , n8722 );
buf ( n8730 , n8725 );
nand ( n8731 , n8729 , n8730 );
nand ( n8732 , n8728 , n8731 );
buf ( n8733 , n4734 );
buf ( n8734 , n8733 );
and ( n8735 , n8732 , n8734 );
not ( n8736 , n8732 );
not ( n8737 , n8733 );
and ( n8738 , n8736 , n8737 );
nor ( n8739 , n8735 , n8738 );
buf ( n8740 , n8343 );
buf ( n8741 , n4735 );
nand ( n8742 , n8740 , n8741 );
buf ( n8743 , n4736 );
buf ( n8744 , n8743 );
and ( n8745 , n8742 , n8744 );
not ( n8746 , n8742 );
not ( n8747 , n8743 );
and ( n8748 , n8746 , n8747 );
nor ( n8749 , n8745 , n8748 );
xor ( n8750 , n8739 , n8749 );
buf ( n8751 , n4737 );
nand ( n8752 , n7126 , n8751 );
buf ( n8753 , n4738 );
buf ( n8754 , n8753 );
and ( n8755 , n8752 , n8754 );
not ( n8756 , n8752 );
not ( n8757 , n8753 );
and ( n8758 , n8756 , n8757 );
nor ( n8759 , n8755 , n8758 );
xnor ( n8760 , n8750 , n8759 );
not ( n8761 , n8760 );
or ( n8762 , n8721 , n8761 );
not ( n8763 , n8720 );
not ( n8764 , n8760 );
nand ( n8765 , n8763 , n8764 );
nand ( n8766 , n8762 , n8765 );
not ( n8767 , n8766 );
buf ( n8768 , n4739 );
buf ( n8769 , n4740 );
buf ( n8770 , n8769 );
not ( n8771 , n8770 );
buf ( n8772 , n4741 );
not ( n8773 , n8772 );
not ( n8774 , n8773 );
or ( n8775 , n8771 , n8774 );
not ( n8776 , n8769 );
buf ( n8777 , n8772 );
nand ( n8778 , n8776 , n8777 );
nand ( n8779 , n8775 , n8778 );
xor ( n8780 , n8768 , n8779 );
buf ( n8781 , n4742 );
buf ( n8782 , n4743 );
not ( n8783 , n8782 );
xor ( n8784 , n8781 , n8783 );
buf ( n8785 , n7477 );
buf ( n8786 , n4744 );
nand ( n8787 , n8785 , n8786 );
xnor ( n8788 , n8784 , n8787 );
xnor ( n8789 , n8780 , n8788 );
not ( n8790 , n8789 );
not ( n8791 , n8790 );
not ( n8792 , n8791 );
not ( n8793 , n8792 );
and ( n8794 , n8767 , n8793 );
and ( n8795 , n8790 , n8766 );
nor ( n8796 , n8794 , n8795 );
not ( n8797 , n8796 );
nand ( n8798 , n8710 , n8797 );
not ( n8799 , n8798 );
buf ( n8800 , n4745 );
buf ( n8801 , n8800 );
not ( n8802 , n8801 );
buf ( n8803 , n4746 );
buf ( n8804 , n8803 );
not ( n8805 , n8804 );
buf ( n8806 , n4747 );
not ( n8807 , n8806 );
not ( n8808 , n8807 );
or ( n8809 , n8805 , n8808 );
not ( n8810 , n8803 );
buf ( n8811 , n8806 );
nand ( n8812 , n8810 , n8811 );
nand ( n8813 , n8809 , n8812 );
buf ( n8814 , n4748 );
not ( n8815 , n8814 );
and ( n8816 , n8813 , n8815 );
not ( n8817 , n8813 );
buf ( n8818 , n8814 );
and ( n8819 , n8817 , n8818 );
nor ( n8820 , n8816 , n8819 );
buf ( n8821 , n6815 );
buf ( n8822 , n4749 );
nand ( n8823 , n8821 , n8822 );
buf ( n8824 , n4750 );
not ( n8825 , n8824 );
and ( n8826 , n8823 , n8825 );
not ( n8827 , n8823 );
buf ( n8828 , n8824 );
and ( n8829 , n8827 , n8828 );
nor ( n8830 , n8826 , n8829 );
xor ( n8831 , n8820 , n8830 );
buf ( n8832 , n4751 );
nand ( n8833 , n6996 , n8832 );
buf ( n8834 , n4752 );
not ( n8835 , n8834 );
and ( n8836 , n8833 , n8835 );
not ( n8837 , n8833 );
buf ( n8838 , n8834 );
and ( n8839 , n8837 , n8838 );
nor ( n8840 , n8836 , n8839 );
xnor ( n8841 , n8831 , n8840 );
not ( n8842 , n8841 );
not ( n8843 , n8842 );
or ( n8844 , n8802 , n8843 );
xor ( n8845 , n8820 , n8830 );
xnor ( n8846 , n8845 , n8840 );
not ( n8847 , n8846 );
or ( n8848 , n8847 , n8801 );
nand ( n8849 , n8844 , n8848 );
buf ( n8850 , n4753 );
buf ( n8851 , n8850 );
not ( n8852 , n8851 );
buf ( n8853 , n4754 );
not ( n8854 , n8853 );
not ( n8855 , n8854 );
or ( n8856 , n8852 , n8855 );
not ( n8857 , n8850 );
buf ( n8858 , n8853 );
nand ( n8859 , n8857 , n8858 );
nand ( n8860 , n8856 , n8859 );
buf ( n8861 , n4755 );
buf ( n8862 , n8861 );
and ( n8863 , n8860 , n8862 );
not ( n8864 , n8860 );
not ( n8865 , n8861 );
and ( n8866 , n8864 , n8865 );
nor ( n8867 , n8863 , n8866 );
buf ( n8868 , n4756 );
nand ( n8869 , n8821 , n8868 );
buf ( n8870 , n4757 );
not ( n8871 , n8870 );
and ( n8872 , n8869 , n8871 );
not ( n8873 , n8869 );
buf ( n8874 , n8870 );
and ( n8875 , n8873 , n8874 );
nor ( n8876 , n8872 , n8875 );
xor ( n8877 , n8867 , n8876 );
buf ( n8878 , n4758 );
nand ( n8879 , n8135 , n8878 );
buf ( n8880 , n4759 );
not ( n8881 , n8880 );
and ( n8882 , n8879 , n8881 );
not ( n8883 , n8879 );
buf ( n8884 , n8880 );
and ( n8885 , n8883 , n8884 );
nor ( n8886 , n8882 , n8885 );
xnor ( n8887 , n8877 , n8886 );
not ( n8888 , n8887 );
buf ( n8889 , n8888 );
xnor ( n8890 , n8849 , n8889 );
buf ( n8891 , n8890 );
not ( n8892 , n8891 );
not ( n8893 , n8892 );
and ( n8894 , n8799 , n8893 );
and ( n8895 , n8798 , n8892 );
nor ( n8896 , n8894 , n8895 );
not ( n8897 , n8896 );
and ( n8898 , n8625 , n8897 );
not ( n8899 , n8625 );
and ( n8900 , n8899 , n8896 );
nor ( n8901 , n8898 , n8900 );
buf ( n8902 , n4760 );
buf ( n8903 , n8902 );
not ( n8904 , n8903 );
buf ( n8905 , n4761 );
buf ( n8906 , n8905 );
not ( n8907 , n8906 );
buf ( n8908 , n4762 );
not ( n8909 , n8908 );
not ( n8910 , n8909 );
or ( n8911 , n8907 , n8910 );
not ( n8912 , n8905 );
buf ( n8913 , n8908 );
nand ( n8914 , n8912 , n8913 );
nand ( n8915 , n8911 , n8914 );
buf ( n8916 , n4763 );
buf ( n8917 , n8916 );
and ( n8918 , n8915 , n8917 );
not ( n8919 , n8915 );
not ( n8920 , n8916 );
and ( n8921 , n8919 , n8920 );
nor ( n8922 , n8918 , n8921 );
buf ( n8923 , n6621 );
buf ( n8924 , n4764 );
nand ( n8925 , n8923 , n8924 );
buf ( n8926 , n4765 );
not ( n8927 , n8926 );
and ( n8928 , n8925 , n8927 );
not ( n8929 , n8925 );
buf ( n8930 , n8926 );
and ( n8931 , n8929 , n8930 );
nor ( n8932 , n8928 , n8931 );
xor ( n8933 , n8922 , n8932 );
buf ( n8934 , n7981 );
buf ( n8935 , n4766 );
nand ( n8936 , n8934 , n8935 );
buf ( n8937 , n4767 );
not ( n8938 , n8937 );
and ( n8939 , n8936 , n8938 );
not ( n8940 , n8936 );
buf ( n8941 , n8937 );
and ( n8942 , n8940 , n8941 );
nor ( n8943 , n8939 , n8942 );
xnor ( n8944 , n8933 , n8943 );
not ( n8945 , n8944 );
buf ( n8946 , n8945 );
not ( n8947 , n8946 );
not ( n8948 , n8947 );
or ( n8949 , n8904 , n8948 );
not ( n8950 , n8945 );
buf ( n8951 , n8950 );
or ( n8952 , n8951 , n8903 );
nand ( n8953 , n8949 , n8952 );
buf ( n8954 , n4768 );
buf ( n8955 , n4769 );
buf ( n8956 , n8955 );
not ( n8957 , n8956 );
buf ( n8958 , n4770 );
not ( n8959 , n8958 );
not ( n8960 , n8959 );
or ( n8961 , n8957 , n8960 );
not ( n8962 , n8955 );
buf ( n8963 , n8958 );
nand ( n8964 , n8962 , n8963 );
nand ( n8965 , n8961 , n8964 );
xor ( n8966 , n8954 , n8965 );
buf ( n8967 , n4771 );
buf ( n8968 , n4772 );
not ( n8969 , n8968 );
xor ( n8970 , n8967 , n8969 );
buf ( n8971 , n7865 );
buf ( n8972 , n4773 );
nand ( n8973 , n8971 , n8972 );
xnor ( n8974 , n8970 , n8973 );
xnor ( n8975 , n8966 , n8974 );
not ( n8976 , n8975 );
buf ( n8977 , n8976 );
and ( n8978 , n8953 , n8977 );
not ( n8979 , n8953 );
not ( n8980 , n8977 );
and ( n8981 , n8979 , n8980 );
nor ( n8982 , n8978 , n8981 );
buf ( n8983 , n4774 );
nand ( n8984 , n8135 , n8983 );
buf ( n8985 , n8984 );
buf ( n8986 , n4775 );
not ( n8987 , n8986 );
and ( n8988 , n8985 , n8987 );
not ( n8989 , n8985 );
buf ( n8990 , n8986 );
and ( n8991 , n8989 , n8990 );
or ( n8992 , n8988 , n8991 );
not ( n8993 , n8992 );
buf ( n8994 , n4776 );
buf ( n8995 , n8994 );
not ( n8996 , n8995 );
buf ( n8997 , n4777 );
not ( n8998 , n8997 );
not ( n8999 , n8998 );
or ( n9000 , n8996 , n8999 );
not ( n9001 , n8994 );
buf ( n9002 , n8997 );
nand ( n9003 , n9001 , n9002 );
nand ( n9004 , n9000 , n9003 );
buf ( n9005 , n4778 );
buf ( n9006 , n9005 );
and ( n9007 , n9004 , n9006 );
not ( n9008 , n9004 );
not ( n9009 , n9005 );
and ( n9010 , n9008 , n9009 );
nor ( n9011 , n9007 , n9010 );
buf ( n9012 , n4779 );
nand ( n9013 , n7412 , n9012 );
buf ( n9014 , n4780 );
buf ( n9015 , n9014 );
and ( n9016 , n9013 , n9015 );
not ( n9017 , n9013 );
not ( n9018 , n9014 );
and ( n9019 , n9017 , n9018 );
nor ( n9020 , n9016 , n9019 );
xor ( n9021 , n9011 , n9020 );
buf ( n9022 , n4781 );
nand ( n9023 , n6945 , n9022 );
buf ( n9024 , n4782 );
not ( n9025 , n9024 );
and ( n9026 , n9023 , n9025 );
not ( n9027 , n9023 );
buf ( n9028 , n9024 );
and ( n9029 , n9027 , n9028 );
nor ( n9030 , n9026 , n9029 );
xnor ( n9031 , n9021 , n9030 );
buf ( n9032 , n9031 );
not ( n9033 , n9032 );
or ( n9034 , n8993 , n9033 );
or ( n9035 , n9032 , n8992 );
nand ( n9036 , n9034 , n9035 );
buf ( n9037 , n4783 );
buf ( n9038 , n9037 );
not ( n9039 , n9038 );
buf ( n9040 , n4784 );
not ( n9041 , n9040 );
not ( n9042 , n9041 );
or ( n9043 , n9039 , n9042 );
not ( n9044 , n9037 );
buf ( n9045 , n9040 );
nand ( n9046 , n9044 , n9045 );
nand ( n9047 , n9043 , n9046 );
buf ( n9048 , n4785 );
buf ( n9049 , n9048 );
and ( n9050 , n9047 , n9049 );
not ( n9051 , n9047 );
not ( n9052 , n9048 );
and ( n9053 , n9051 , n9052 );
nor ( n9054 , n9050 , n9053 );
buf ( n9055 , n4786 );
nand ( n9056 , n7477 , n9055 );
buf ( n9057 , n4787 );
buf ( n9058 , n9057 );
and ( n9059 , n9056 , n9058 );
not ( n9060 , n9056 );
not ( n9061 , n9057 );
and ( n9062 , n9060 , n9061 );
nor ( n9063 , n9059 , n9062 );
xor ( n9064 , n9054 , n9063 );
buf ( n9065 , n4788 );
nand ( n9066 , n7094 , n9065 );
buf ( n9067 , n4789 );
not ( n9068 , n9067 );
and ( n9069 , n9066 , n9068 );
not ( n9070 , n9066 );
buf ( n9071 , n9067 );
and ( n9072 , n9070 , n9071 );
nor ( n9073 , n9069 , n9072 );
xnor ( n9074 , n9064 , n9073 );
buf ( n9075 , n9074 );
not ( n9076 , n9075 );
and ( n9077 , n9036 , n9076 );
not ( n9078 , n9036 );
and ( n9079 , n9078 , n9075 );
or ( n9080 , n9077 , n9079 );
nand ( n9081 , n8982 , n9080 );
not ( n9082 , n9081 );
buf ( n9083 , n4790 );
buf ( n9084 , n9083 );
not ( n9085 , n9084 );
buf ( n9086 , n4791 );
buf ( n9087 , n9086 );
not ( n9088 , n9087 );
buf ( n9089 , n4792 );
not ( n9090 , n9089 );
not ( n9091 , n9090 );
or ( n9092 , n9088 , n9091 );
not ( n9093 , n9086 );
buf ( n9094 , n9089 );
nand ( n9095 , n9093 , n9094 );
nand ( n9096 , n9092 , n9095 );
buf ( n9097 , n4793 );
buf ( n9098 , n9097 );
and ( n9099 , n9096 , n9098 );
not ( n9100 , n9096 );
not ( n9101 , n9097 );
and ( n9102 , n9100 , n9101 );
nor ( n9103 , n9099 , n9102 );
buf ( n9104 , n4794 );
nand ( n9105 , n6933 , n9104 );
buf ( n9106 , n4795 );
buf ( n9107 , n9106 );
and ( n9108 , n9105 , n9107 );
not ( n9109 , n9105 );
not ( n9110 , n9106 );
and ( n9111 , n9109 , n9110 );
nor ( n9112 , n9108 , n9111 );
xor ( n9113 , n9103 , n9112 );
buf ( n9114 , n4796 );
nand ( n9115 , n6804 , n9114 );
buf ( n9116 , n4797 );
not ( n9117 , n9116 );
and ( n9118 , n9115 , n9117 );
not ( n9119 , n9115 );
buf ( n9120 , n9116 );
and ( n9121 , n9119 , n9120 );
nor ( n9122 , n9118 , n9121 );
xnor ( n9123 , n9113 , n9122 );
not ( n9124 , n9123 );
not ( n9125 , n9124 );
or ( n9126 , n9085 , n9125 );
not ( n9127 , n9124 );
not ( n9128 , n9083 );
nand ( n9129 , n9127 , n9128 );
nand ( n9130 , n9126 , n9129 );
buf ( n9131 , n4798 );
buf ( n9132 , n9131 );
not ( n9133 , n9132 );
buf ( n9134 , n4799 );
not ( n9135 , n9134 );
not ( n9136 , n9135 );
or ( n9137 , n9133 , n9136 );
not ( n9138 , n9131 );
buf ( n9139 , n9134 );
nand ( n9140 , n9138 , n9139 );
nand ( n9141 , n9137 , n9140 );
buf ( n9142 , n4800 );
not ( n9143 , n9142 );
and ( n9144 , n9141 , n9143 );
not ( n9145 , n9141 );
buf ( n9146 , n9142 );
and ( n9147 , n9145 , n9146 );
nor ( n9148 , n9144 , n9147 );
buf ( n9149 , n4801 );
nand ( n9150 , n7093 , n9149 );
buf ( n9151 , n4802 );
buf ( n9152 , n9151 );
and ( n9153 , n9150 , n9152 );
not ( n9154 , n9150 );
not ( n9155 , n9151 );
and ( n9156 , n9154 , n9155 );
nor ( n9157 , n9153 , n9156 );
xor ( n9158 , n9148 , n9157 );
buf ( n9159 , n7412 );
buf ( n9160 , n4803 );
nand ( n9161 , n9159 , n9160 );
buf ( n9162 , n4804 );
not ( n9163 , n9162 );
and ( n9164 , n9161 , n9163 );
not ( n9165 , n9161 );
buf ( n9166 , n9162 );
and ( n9167 , n9165 , n9166 );
nor ( n9168 , n9164 , n9167 );
xnor ( n9169 , n9158 , n9168 );
buf ( n9170 , n9169 );
not ( n9171 , n9170 );
and ( n9172 , n9130 , n9171 );
not ( n9173 , n9130 );
and ( n9174 , n9173 , n9170 );
nor ( n9175 , n9172 , n9174 );
not ( n9176 , n9175 );
and ( n9177 , n9082 , n9176 );
and ( n9178 , n9081 , n9175 );
nor ( n9179 , n9177 , n9178 );
buf ( n9180 , n4805 );
buf ( n9181 , n9180 );
buf ( n9182 , n4806 );
buf ( n9183 , n9182 );
not ( n9184 , n9183 );
buf ( n9185 , n4807 );
not ( n9186 , n9185 );
not ( n9187 , n9186 );
or ( n9188 , n9184 , n9187 );
not ( n9189 , n9182 );
buf ( n9190 , n9185 );
nand ( n9191 , n9189 , n9190 );
nand ( n9192 , n9188 , n9191 );
buf ( n9193 , n4808 );
not ( n9194 , n9193 );
and ( n9195 , n9192 , n9194 );
not ( n9196 , n9192 );
buf ( n9197 , n9193 );
and ( n9198 , n9196 , n9197 );
nor ( n9199 , n9195 , n9198 );
buf ( n9200 , n4809 );
nand ( n9201 , n7195 , n9200 );
buf ( n9202 , n4810 );
buf ( n9203 , n9202 );
and ( n9204 , n9201 , n9203 );
not ( n9205 , n9201 );
not ( n9206 , n9202 );
and ( n9207 , n9205 , n9206 );
nor ( n9208 , n9204 , n9207 );
xor ( n9209 , n9199 , n9208 );
buf ( n9210 , n4811 );
nand ( n9211 , n7094 , n9210 );
buf ( n9212 , n4812 );
not ( n9213 , n9212 );
and ( n9214 , n9211 , n9213 );
not ( n9215 , n9211 );
buf ( n9216 , n9212 );
and ( n9217 , n9215 , n9216 );
nor ( n9218 , n9214 , n9217 );
xnor ( n9219 , n9209 , n9218 );
not ( n9220 , n9219 );
not ( n9221 , n9220 );
xor ( n9222 , n9181 , n9221 );
buf ( n9223 , n4813 );
buf ( n9224 , n9223 );
buf ( n9225 , n4814 );
buf ( n9226 , n9225 );
not ( n9227 , n9226 );
buf ( n9228 , n4815 );
not ( n9229 , n9228 );
not ( n9230 , n9229 );
or ( n9231 , n9227 , n9230 );
not ( n9232 , n9225 );
buf ( n9233 , n9228 );
nand ( n9234 , n9232 , n9233 );
nand ( n9235 , n9231 , n9234 );
xor ( n9236 , n9224 , n9235 );
buf ( n9237 , n4816 );
buf ( n9238 , n4817 );
xor ( n9239 , n9237 , n9238 );
buf ( n9240 , n4818 );
nand ( n9241 , n8520 , n9240 );
xnor ( n9242 , n9239 , n9241 );
xnor ( n9243 , n9236 , n9242 );
buf ( n9244 , n9243 );
xnor ( n9245 , n9222 , n9244 );
not ( n9246 , n8439 );
buf ( n9247 , n4819 );
nand ( n9248 , n8821 , n9247 );
buf ( n9249 , n4820 );
buf ( n9250 , n9249 );
and ( n9251 , n9248 , n9250 );
not ( n9252 , n9248 );
not ( n9253 , n9249 );
and ( n9254 , n9252 , n9253 );
nor ( n9255 , n9251 , n9254 );
not ( n9256 , n9255 );
buf ( n9257 , n8134 );
buf ( n9258 , n4821 );
nand ( n9259 , n9257 , n9258 );
buf ( n9260 , n4822 );
not ( n9261 , n9260 );
and ( n9262 , n9259 , n9261 );
not ( n9263 , n9259 );
buf ( n9264 , n9260 );
and ( n9265 , n9263 , n9264 );
nor ( n9266 , n9262 , n9265 );
not ( n9267 , n9266 );
or ( n9268 , n9256 , n9267 );
or ( n9269 , n9255 , n9266 );
nand ( n9270 , n9268 , n9269 );
buf ( n9271 , n4823 );
buf ( n9272 , n9271 );
not ( n9273 , n9272 );
buf ( n9274 , n4824 );
not ( n9275 , n9274 );
not ( n9276 , n9275 );
or ( n9277 , n9273 , n9276 );
not ( n9278 , n9271 );
buf ( n9279 , n9274 );
nand ( n9280 , n9278 , n9279 );
nand ( n9281 , n9277 , n9280 );
buf ( n9282 , n4825 );
not ( n9283 , n9282 );
and ( n9284 , n9281 , n9283 );
not ( n9285 , n9281 );
buf ( n9286 , n9282 );
and ( n9287 , n9285 , n9286 );
nor ( n9288 , n9284 , n9287 );
and ( n9289 , n9270 , n9288 );
not ( n9290 , n9270 );
not ( n9291 , n9288 );
and ( n9292 , n9290 , n9291 );
nor ( n9293 , n9289 , n9292 );
buf ( n9294 , n9293 );
not ( n9295 , n9294 );
or ( n9296 , n9246 , n9295 );
not ( n9297 , n8439 );
not ( n9298 , n9255 );
xor ( n9299 , n9288 , n9298 );
buf ( n9300 , n9266 );
xnor ( n9301 , n9299 , n9300 );
buf ( n9302 , n9301 );
nand ( n9303 , n9297 , n9302 );
nand ( n9304 , n9296 , n9303 );
buf ( n9305 , n4826 );
buf ( n9306 , n9305 );
not ( n9307 , n9306 );
buf ( n9308 , n4827 );
not ( n9309 , n9308 );
not ( n9310 , n9309 );
or ( n9311 , n9307 , n9310 );
not ( n9312 , n9305 );
buf ( n9313 , n9308 );
nand ( n9314 , n9312 , n9313 );
nand ( n9315 , n9311 , n9314 );
buf ( n9316 , n4828 );
not ( n9317 , n9316 );
and ( n9318 , n9315 , n9317 );
not ( n9319 , n9315 );
buf ( n9320 , n9316 );
and ( n9321 , n9319 , n9320 );
nor ( n9322 , n9318 , n9321 );
buf ( n9323 , n4829 );
nand ( n9324 , n7195 , n9323 );
buf ( n9325 , n4830 );
buf ( n9326 , n9325 );
and ( n9327 , n9324 , n9326 );
not ( n9328 , n9324 );
not ( n9329 , n9325 );
and ( n9330 , n9328 , n9329 );
nor ( n9331 , n9327 , n9330 );
xor ( n9332 , n9322 , n9331 );
buf ( n9333 , n4831 );
nand ( n9334 , n6985 , n9333 );
buf ( n9335 , n4832 );
buf ( n9336 , n9335 );
and ( n9337 , n9334 , n9336 );
not ( n9338 , n9334 );
not ( n9339 , n9335 );
and ( n9340 , n9338 , n9339 );
nor ( n9341 , n9337 , n9340 );
xnor ( n9342 , n9332 , n9341 );
not ( n9343 , n9342 );
not ( n9344 , n9343 );
and ( n9345 , n9304 , n9344 );
not ( n9346 , n9304 );
buf ( n9347 , n9342 );
not ( n9348 , n9347 );
and ( n9349 , n9346 , n9348 );
nor ( n9350 , n9345 , n9349 );
nand ( n9351 , n9245 , n9350 );
buf ( n9352 , n4833 );
buf ( n9353 , n9352 );
not ( n9354 , n9353 );
buf ( n9355 , n4834 );
buf ( n9356 , n9355 );
not ( n9357 , n9356 );
buf ( n9358 , n4835 );
not ( n9359 , n9358 );
not ( n9360 , n9359 );
or ( n9361 , n9357 , n9360 );
not ( n9362 , n9355 );
buf ( n9363 , n9358 );
nand ( n9364 , n9362 , n9363 );
nand ( n9365 , n9361 , n9364 );
buf ( n9366 , n4836 );
not ( n9367 , n9366 );
and ( n9368 , n9365 , n9367 );
not ( n9369 , n9365 );
buf ( n9370 , n9366 );
and ( n9371 , n9369 , n9370 );
nor ( n9372 , n9368 , n9371 );
buf ( n9373 , n4837 );
nand ( n9374 , n7401 , n9373 );
buf ( n9375 , n4838 );
buf ( n9376 , n9375 );
and ( n9377 , n9374 , n9376 );
not ( n9378 , n9374 );
not ( n9379 , n9375 );
and ( n9380 , n9378 , n9379 );
nor ( n9381 , n9377 , n9380 );
xor ( n9382 , n9372 , n9381 );
buf ( n9383 , n4839 );
nand ( n9384 , n7442 , n9383 );
buf ( n9385 , n4840 );
not ( n9386 , n9385 );
and ( n9387 , n9384 , n9386 );
not ( n9388 , n9384 );
buf ( n9389 , n9385 );
and ( n9390 , n9388 , n9389 );
nor ( n9391 , n9387 , n9390 );
xnor ( n9392 , n9382 , n9391 );
not ( n9393 , n9392 );
not ( n9394 , n9393 );
not ( n9395 , n9394 );
or ( n9396 , n9354 , n9395 );
not ( n9397 , n9392 );
not ( n9398 , n9352 );
nand ( n9399 , n9397 , n9398 );
nand ( n9400 , n9396 , n9399 );
not ( n9401 , n7660 );
xor ( n9402 , n7651 , n9401 );
xnor ( n9403 , n9402 , n7670 );
not ( n9404 , n9403 );
not ( n9405 , n9404 );
and ( n9406 , n9400 , n9405 );
not ( n9407 , n9400 );
and ( n9408 , n9407 , n7672 );
nor ( n9409 , n9406 , n9408 );
not ( n9410 , n9409 );
and ( n9411 , n9351 , n9410 );
not ( n9412 , n9351 );
and ( n9413 , n9412 , n9409 );
nor ( n9414 , n9411 , n9413 );
xor ( n9415 , n9179 , n9414 );
and ( n9416 , n8901 , n9415 );
not ( n9417 , n8901 );
not ( n9418 , n9415 );
and ( n9419 , n9417 , n9418 );
nor ( n9420 , n9416 , n9419 );
not ( n9421 , n9420 );
not ( n9422 , n9421 );
not ( n9423 , n9422 );
and ( n9424 , n8095 , n9423 );
not ( n9425 , n8095 );
not ( n9426 , n9420 );
buf ( n9427 , n9426 );
not ( n9428 , n9427 );
and ( n9429 , n9425 , n9428 );
nor ( n9430 , n9424 , n9429 );
not ( n9431 , n8801 );
buf ( n9432 , n4841 );
not ( n9433 , n9432 );
not ( n9434 , n9433 );
or ( n9435 , n9431 , n9434 );
not ( n9436 , n8800 );
buf ( n9437 , n9432 );
nand ( n9438 , n9436 , n9437 );
nand ( n9439 , n9435 , n9438 );
buf ( n9440 , n4842 );
buf ( n9441 , n9440 );
and ( n9442 , n9439 , n9441 );
not ( n9443 , n9439 );
not ( n9444 , n9440 );
and ( n9445 , n9443 , n9444 );
nor ( n9446 , n9442 , n9445 );
not ( n9447 , n9446 );
buf ( n9448 , n4843 );
nand ( n9449 , n7412 , n9448 );
buf ( n9450 , n4844 );
buf ( n9451 , n9450 );
and ( n9452 , n9449 , n9451 );
not ( n9453 , n9449 );
not ( n9454 , n9450 );
and ( n9455 , n9453 , n9454 );
nor ( n9456 , n9452 , n9455 );
xor ( n9457 , n9447 , n9456 );
buf ( n9458 , n4845 );
nand ( n9459 , n7134 , n9458 );
buf ( n9460 , n4846 );
buf ( n9461 , n9460 );
and ( n9462 , n9459 , n9461 );
not ( n9463 , n9459 );
not ( n9464 , n9460 );
and ( n9465 , n9463 , n9464 );
nor ( n9466 , n9462 , n9465 );
xnor ( n9467 , n9457 , n9466 );
buf ( n9468 , n9467 );
xor ( n9469 , n6968 , n9468 );
buf ( n9470 , n4847 );
not ( n9471 , n9470 );
buf ( n9472 , n4848 );
not ( n9473 , n9472 );
buf ( n9474 , n4849 );
buf ( n9475 , n9474 );
and ( n9476 , n9473 , n9475 );
not ( n9477 , n9473 );
not ( n9478 , n9474 );
and ( n9479 , n9477 , n9478 );
nor ( n9480 , n9476 , n9479 );
xor ( n9481 , n9471 , n9480 );
buf ( n9482 , n4850 );
buf ( n9483 , n4851 );
xor ( n9484 , n9482 , n9483 );
buf ( n9485 , n4852 );
nand ( n9486 , n8971 , n9485 );
xnor ( n9487 , n9484 , n9486 );
xnor ( n9488 , n9481 , n9487 );
buf ( n9489 , n9488 );
xnor ( n9490 , n9469 , n9489 );
buf ( n9491 , n4853 );
buf ( n9492 , n9491 );
not ( n9493 , n9492 );
buf ( n9494 , n4854 );
buf ( n9495 , n9494 );
not ( n9496 , n9495 );
buf ( n9497 , n4855 );
not ( n9498 , n9497 );
not ( n9499 , n9498 );
or ( n9500 , n9496 , n9499 );
not ( n9501 , n9494 );
buf ( n9502 , n9497 );
nand ( n9503 , n9501 , n9502 );
nand ( n9504 , n9500 , n9503 );
buf ( n9505 , n4856 );
not ( n9506 , n9505 );
and ( n9507 , n9504 , n9506 );
not ( n9508 , n9504 );
buf ( n9509 , n9505 );
and ( n9510 , n9508 , n9509 );
nor ( n9511 , n9507 , n9510 );
buf ( n9512 , n4857 );
nand ( n9513 , n7515 , n9512 );
buf ( n9514 , n4858 );
buf ( n9515 , n9514 );
and ( n9516 , n9513 , n9515 );
not ( n9517 , n9513 );
not ( n9518 , n9514 );
and ( n9519 , n9517 , n9518 );
nor ( n9520 , n9516 , n9519 );
xor ( n9521 , n9511 , n9520 );
buf ( n9522 , n4859 );
nand ( n9523 , n7617 , n9522 );
buf ( n9524 , n4860 );
buf ( n9525 , n9524 );
and ( n9526 , n9523 , n9525 );
not ( n9527 , n9523 );
not ( n9528 , n9524 );
and ( n9529 , n9527 , n9528 );
nor ( n9530 , n9526 , n9529 );
xnor ( n9531 , n9521 , n9530 );
not ( n9532 , n9531 );
not ( n9533 , n9532 );
or ( n9534 , n9493 , n9533 );
or ( n9535 , n9492 , n9532 );
nand ( n9536 , n9534 , n9535 );
not ( n9537 , n7207 );
not ( n9538 , n9537 );
and ( n9539 , n9536 , n9538 );
not ( n9540 , n9536 );
xor ( n9541 , n7181 , n7205 );
not ( n9542 , n7193 );
xnor ( n9543 , n9541 , n9542 );
buf ( n9544 , n9543 );
and ( n9545 , n9540 , n9544 );
nor ( n9546 , n9539 , n9545 );
not ( n9547 , n9546 );
nand ( n9548 , n9490 , n9547 );
buf ( n9549 , n4861 );
nand ( n9550 , n8134 , n9549 );
buf ( n9551 , n4862 );
buf ( n9552 , n9551 );
and ( n9553 , n9550 , n9552 );
not ( n9554 , n9550 );
not ( n9555 , n9551 );
and ( n9556 , n9554 , n9555 );
nor ( n9557 , n9553 , n9556 );
buf ( n9558 , n9557 );
not ( n9559 , n9558 );
buf ( n9560 , n4863 );
buf ( n9561 , n9560 );
not ( n9562 , n9561 );
buf ( n9563 , n4864 );
not ( n9564 , n9563 );
not ( n9565 , n9564 );
or ( n9566 , n9562 , n9565 );
not ( n9567 , n9560 );
buf ( n9568 , n9563 );
nand ( n9569 , n9567 , n9568 );
nand ( n9570 , n9566 , n9569 );
buf ( n9571 , n4865 );
not ( n9572 , n9571 );
and ( n9573 , n9570 , n9572 );
not ( n9574 , n9570 );
buf ( n9575 , n9571 );
and ( n9576 , n9574 , n9575 );
nor ( n9577 , n9573 , n9576 );
buf ( n9578 , n4866 );
nand ( n9579 , n7043 , n9578 );
buf ( n9580 , n4867 );
buf ( n9581 , n9580 );
and ( n9582 , n9579 , n9581 );
not ( n9583 , n9579 );
not ( n9584 , n9580 );
and ( n9585 , n9583 , n9584 );
nor ( n9586 , n9582 , n9585 );
xor ( n9587 , n9577 , n9586 );
buf ( n9588 , n4868 );
nand ( n9589 , n7471 , n9588 );
buf ( n9590 , n4869 );
buf ( n9591 , n9590 );
and ( n9592 , n9589 , n9591 );
not ( n9593 , n9589 );
not ( n9594 , n9590 );
and ( n9595 , n9593 , n9594 );
nor ( n9596 , n9592 , n9595 );
xnor ( n9597 , n9587 , n9596 );
not ( n9598 , n9597 );
or ( n9599 , n9559 , n9598 );
or ( n9600 , n9597 , n9558 );
nand ( n9601 , n9599 , n9600 );
not ( n9602 , n9601 );
not ( n9603 , n9602 );
buf ( n9604 , n4870 );
buf ( n9605 , n9604 );
buf ( n9606 , n4871 );
not ( n9607 , n9606 );
buf ( n9608 , n4872 );
buf ( n9609 , n9608 );
and ( n9610 , n9607 , n9609 );
not ( n9611 , n9607 );
not ( n9612 , n9608 );
and ( n9613 , n9611 , n9612 );
nor ( n9614 , n9610 , n9613 );
xor ( n9615 , n9605 , n9614 );
buf ( n9616 , n4873 );
buf ( n9617 , n4874 );
xor ( n9618 , n9616 , n9617 );
buf ( n9619 , n8387 );
buf ( n9620 , n4875 );
nand ( n9621 , n9619 , n9620 );
xnor ( n9622 , n9618 , n9621 );
xnor ( n9623 , n9615 , n9622 );
buf ( n9624 , n9623 );
not ( n9625 , n9624 );
or ( n9626 , n9603 , n9625 );
not ( n9627 , n9604 );
xor ( n9628 , n9627 , n9614 );
xnor ( n9629 , n9628 , n9622 );
buf ( n9630 , n9629 );
nand ( n9631 , n9630 , n9601 );
nand ( n9632 , n9626 , n9631 );
not ( n9633 , n9632 );
and ( n9634 , n9548 , n9633 );
not ( n9635 , n9548 );
and ( n9636 , n9635 , n9632 );
nor ( n9637 , n9634 , n9636 );
not ( n9638 , n9637 );
nand ( n9639 , n9633 , n9546 );
not ( n9640 , n9639 );
buf ( n9641 , n4876 );
nand ( n9642 , n7909 , n9641 );
buf ( n9643 , n4877 );
xor ( n9644 , n9642 , n9643 );
not ( n9645 , n9644 );
not ( n9646 , n8433 );
or ( n9647 , n9645 , n9646 );
or ( n9648 , n8433 , n9644 );
nand ( n9649 , n9647 , n9648 );
buf ( n9650 , n4878 );
buf ( n9651 , n9650 );
not ( n9652 , n9651 );
buf ( n9653 , n4879 );
not ( n9654 , n9653 );
not ( n9655 , n9654 );
or ( n9656 , n9652 , n9655 );
not ( n9657 , n9650 );
buf ( n9658 , n9653 );
nand ( n9659 , n9657 , n9658 );
nand ( n9660 , n9656 , n9659 );
buf ( n9661 , n4880 );
buf ( n9662 , n9661 );
and ( n9663 , n9660 , n9662 );
not ( n9664 , n9660 );
not ( n9665 , n9661 );
and ( n9666 , n9664 , n9665 );
nor ( n9667 , n9663 , n9666 );
buf ( n9668 , n4881 );
nand ( n9669 , n8223 , n9668 );
buf ( n9670 , n4882 );
buf ( n9671 , n9670 );
and ( n9672 , n9669 , n9671 );
not ( n9673 , n9669 );
not ( n9674 , n9670 );
and ( n9675 , n9673 , n9674 );
nor ( n9676 , n9672 , n9675 );
xor ( n9677 , n9667 , n9676 );
buf ( n9678 , n4883 );
nand ( n9679 , n6934 , n9678 );
buf ( n9680 , n4884 );
buf ( n9681 , n9680 );
and ( n9682 , n9679 , n9681 );
not ( n9683 , n9679 );
not ( n9684 , n9680 );
and ( n9685 , n9683 , n9684 );
nor ( n9686 , n9682 , n9685 );
xnor ( n9687 , n9677 , n9686 );
not ( n9688 , n9687 );
not ( n9689 , n9688 );
and ( n9690 , n9649 , n9689 );
not ( n9691 , n9649 );
and ( n9692 , n9691 , n9688 );
nor ( n9693 , n9690 , n9692 );
not ( n9694 , n9693 );
not ( n9695 , n9694 );
and ( n9696 , n9640 , n9695 );
and ( n9697 , n9639 , n9694 );
nor ( n9698 , n9696 , n9697 );
not ( n9699 , n9698 );
buf ( n9700 , n4885 );
xor ( n9701 , n9700 , n7990 );
buf ( n9702 , n4886 );
nand ( n9703 , n7184 , n9702 );
buf ( n9704 , n4887 );
not ( n9705 , n9704 );
and ( n9706 , n9703 , n9705 );
not ( n9707 , n9703 );
buf ( n9708 , n9704 );
and ( n9709 , n9707 , n9708 );
nor ( n9710 , n9706 , n9709 );
xnor ( n9711 , n9701 , n9710 );
not ( n9712 , n9711 );
buf ( n9713 , n4888 );
not ( n9714 , n9713 );
not ( n9715 , n9714 );
buf ( n9716 , n4889 );
not ( n9717 , n9716 );
and ( n9718 , n9715 , n9717 );
and ( n9719 , n9716 , n9714 );
nor ( n9720 , n9718 , n9719 );
not ( n9721 , n9720 );
and ( n9722 , n9712 , n9721 );
and ( n9723 , n9711 , n9720 );
nor ( n9724 , n9722 , n9723 );
buf ( n9725 , n9724 );
not ( n9726 , n9725 );
buf ( n9727 , n4890 );
nand ( n9728 , n8821 , n9727 );
buf ( n9729 , n4891 );
buf ( n9730 , n9729 );
and ( n9731 , n9728 , n9730 );
not ( n9732 , n9728 );
not ( n9733 , n9729 );
and ( n9734 , n9732 , n9733 );
nor ( n9735 , n9731 , n9734 );
not ( n9736 , n9735 );
not ( n9737 , n9736 );
buf ( n9738 , n4892 );
buf ( n9739 , n9738 );
not ( n9740 , n9739 );
buf ( n9741 , n4893 );
not ( n9742 , n9741 );
not ( n9743 , n9742 );
or ( n9744 , n9740 , n9743 );
not ( n9745 , n9738 );
buf ( n9746 , n9741 );
nand ( n9747 , n9745 , n9746 );
nand ( n9748 , n9744 , n9747 );
buf ( n9749 , n4894 );
not ( n9750 , n9749 );
and ( n9751 , n9748 , n9750 );
not ( n9752 , n9748 );
buf ( n9753 , n9749 );
and ( n9754 , n9752 , n9753 );
nor ( n9755 , n9751 , n9754 );
buf ( n9756 , n4895 );
nand ( n9757 , n7043 , n9756 );
buf ( n9758 , n4896 );
buf ( n9759 , n9758 );
and ( n9760 , n9757 , n9759 );
not ( n9761 , n9757 );
not ( n9762 , n9758 );
and ( n9763 , n9761 , n9762 );
nor ( n9764 , n9760 , n9763 );
xor ( n9765 , n9755 , n9764 );
buf ( n9766 , n4897 );
nand ( n9767 , n7785 , n9766 );
buf ( n9768 , n4898 );
buf ( n9769 , n9768 );
and ( n9770 , n9767 , n9769 );
not ( n9771 , n9767 );
not ( n9772 , n9768 );
and ( n9773 , n9771 , n9772 );
nor ( n9774 , n9770 , n9773 );
xnor ( n9775 , n9765 , n9774 );
not ( n9776 , n9775 );
not ( n9777 , n9776 );
or ( n9778 , n9737 , n9777 );
not ( n9779 , n9736 );
buf ( n9780 , n9775 );
nand ( n9781 , n9779 , n9780 );
nand ( n9782 , n9778 , n9781 );
not ( n9783 , n9782 );
and ( n9784 , n9726 , n9783 );
and ( n9785 , n9725 , n9782 );
nor ( n9786 , n9784 , n9785 );
not ( n9787 , n9786 );
not ( n9788 , n9787 );
not ( n9789 , n8792 );
buf ( n9790 , n4899 );
buf ( n9791 , n9790 );
not ( n9792 , n9791 );
not ( n9793 , n8760 );
or ( n9794 , n9792 , n9793 );
not ( n9795 , n9791 );
nand ( n9796 , n9795 , n8764 );
nand ( n9797 , n9794 , n9796 );
not ( n9798 , n9797 );
or ( n9799 , n9789 , n9798 );
not ( n9800 , n8789 );
or ( n9801 , n9800 , n9797 );
nand ( n9802 , n9799 , n9801 );
buf ( n9803 , n4900 );
nand ( n9804 , n7477 , n9803 );
buf ( n9805 , n4901 );
buf ( n9806 , n9805 );
and ( n9807 , n9804 , n9806 );
not ( n9808 , n9804 );
not ( n9809 , n9805 );
and ( n9810 , n9808 , n9809 );
nor ( n9811 , n9807 , n9810 );
buf ( n9812 , n9811 );
not ( n9813 , n9812 );
not ( n9814 , n9813 );
buf ( n9815 , n4902 );
buf ( n9816 , n9815 );
not ( n9817 , n9816 );
not ( n9818 , n7631 );
not ( n9819 , n9818 );
or ( n9820 , n9817 , n9819 );
not ( n9821 , n9815 );
nand ( n9822 , n9821 , n7632 );
nand ( n9823 , n9820 , n9822 );
buf ( n9824 , n4903 );
buf ( n9825 , n9824 );
and ( n9826 , n9823 , n9825 );
not ( n9827 , n9823 );
not ( n9828 , n9824 );
and ( n9829 , n9827 , n9828 );
nor ( n9830 , n9826 , n9829 );
buf ( n9831 , n4904 );
nand ( n9832 , n7288 , n9831 );
buf ( n9833 , n4905 );
buf ( n9834 , n9833 );
and ( n9835 , n9832 , n9834 );
not ( n9836 , n9832 );
not ( n9837 , n9833 );
and ( n9838 , n9836 , n9837 );
nor ( n9839 , n9835 , n9838 );
xor ( n9840 , n9830 , n9839 );
buf ( n9841 , n4906 );
nand ( n9842 , n6816 , n9841 );
buf ( n9843 , n4907 );
buf ( n9844 , n9843 );
and ( n9845 , n9842 , n9844 );
not ( n9846 , n9842 );
not ( n9847 , n9843 );
and ( n9848 , n9846 , n9847 );
nor ( n9849 , n9845 , n9848 );
xnor ( n9850 , n9840 , n9849 );
not ( n9851 , n9850 );
or ( n9852 , n9814 , n9851 );
xor ( n9853 , n9830 , n9849 );
not ( n9854 , n9839 );
xnor ( n9855 , n9853 , n9854 );
nand ( n9856 , n9855 , n9812 );
nand ( n9857 , n9852 , n9856 );
not ( n9858 , n9857 );
buf ( n9859 , n4908 );
buf ( n9860 , n9859 );
not ( n9861 , n9860 );
buf ( n9862 , n4909 );
not ( n9863 , n9862 );
not ( n9864 , n9863 );
or ( n9865 , n9861 , n9864 );
not ( n9866 , n9859 );
buf ( n9867 , n9862 );
nand ( n9868 , n9866 , n9867 );
nand ( n9869 , n9865 , n9868 );
buf ( n9870 , n4910 );
not ( n9871 , n9870 );
and ( n9872 , n9869 , n9871 );
not ( n9873 , n9869 );
buf ( n9874 , n9870 );
and ( n9875 , n9873 , n9874 );
nor ( n9876 , n9872 , n9875 );
buf ( n9877 , n4911 );
nand ( n9878 , n6934 , n9877 );
buf ( n9879 , n4912 );
buf ( n9880 , n9879 );
and ( n9881 , n9878 , n9880 );
not ( n9882 , n9878 );
not ( n9883 , n9879 );
and ( n9884 , n9882 , n9883 );
nor ( n9885 , n9881 , n9884 );
xor ( n9886 , n9876 , n9885 );
buf ( n9887 , n4913 );
nand ( n9888 , n9159 , n9887 );
buf ( n9889 , n4914 );
buf ( n9890 , n9889 );
and ( n9891 , n9888 , n9890 );
not ( n9892 , n9888 );
not ( n9893 , n9889 );
and ( n9894 , n9892 , n9893 );
nor ( n9895 , n9891 , n9894 );
xnor ( n9896 , n9886 , n9895 );
not ( n9897 , n9896 );
not ( n9898 , n9897 );
and ( n9899 , n9858 , n9898 );
and ( n9900 , n9857 , n9897 );
nor ( n9901 , n9899 , n9900 );
nand ( n9902 , n9802 , n9901 );
not ( n9903 , n9902 );
or ( n9904 , n9788 , n9903 );
or ( n9905 , n9787 , n9902 );
nand ( n9906 , n9904 , n9905 );
not ( n9907 , n9906 );
or ( n9908 , n9699 , n9907 );
or ( n9909 , n9906 , n9698 );
nand ( n9910 , n9908 , n9909 );
buf ( n9911 , n4915 );
buf ( n9912 , n9911 );
not ( n9913 , n9912 );
buf ( n9914 , n4916 );
not ( n9915 , n9914 );
not ( n9916 , n9915 );
or ( n9917 , n9913 , n9916 );
not ( n9918 , n9911 );
buf ( n9919 , n9914 );
nand ( n9920 , n9918 , n9919 );
nand ( n9921 , n9917 , n9920 );
buf ( n9922 , n4917 );
buf ( n9923 , n9922 );
and ( n9924 , n9921 , n9923 );
not ( n9925 , n9921 );
not ( n9926 , n9922 );
and ( n9927 , n9925 , n9926 );
nor ( n9928 , n9924 , n9927 );
buf ( n9929 , n4918 );
nand ( n9930 , n6863 , n9929 );
buf ( n9931 , n4919 );
buf ( n9932 , n9931 );
and ( n9933 , n9930 , n9932 );
not ( n9934 , n9930 );
not ( n9935 , n9931 );
and ( n9936 , n9934 , n9935 );
nor ( n9937 , n9933 , n9936 );
xor ( n9938 , n9928 , n9937 );
buf ( n9939 , n4920 );
nand ( n9940 , n7750 , n9939 );
buf ( n9941 , n4921 );
not ( n9942 , n9941 );
and ( n9943 , n9940 , n9942 );
not ( n9944 , n9940 );
buf ( n9945 , n9941 );
and ( n9946 , n9944 , n9945 );
nor ( n9947 , n9943 , n9946 );
xnor ( n9948 , n9938 , n9947 );
not ( n9949 , n9948 );
not ( n9950 , n9949 );
xor ( n9951 , n7375 , n9950 );
buf ( n9952 , n4922 );
buf ( n9953 , n4923 );
buf ( n9954 , n9953 );
not ( n9955 , n9954 );
buf ( n9956 , n4924 );
not ( n9957 , n9956 );
not ( n9958 , n9957 );
or ( n9959 , n9955 , n9958 );
not ( n9960 , n9953 );
buf ( n9961 , n9956 );
nand ( n9962 , n9960 , n9961 );
nand ( n9963 , n9959 , n9962 );
xor ( n9964 , n9952 , n9963 );
buf ( n9965 , n4925 );
buf ( n9966 , n4926 );
not ( n9967 , n9966 );
xor ( n9968 , n9965 , n9967 );
buf ( n9969 , n4927 );
nand ( n9970 , n7617 , n9969 );
xnor ( n9971 , n9968 , n9970 );
xnor ( n9972 , n9964 , n9971 );
not ( n9973 , n9972 );
not ( n9974 , n9973 );
xnor ( n9975 , n9951 , n9974 );
not ( n9976 , n9975 );
buf ( n9977 , n4928 );
buf ( n9978 , n9977 );
not ( n9979 , n9978 );
buf ( n9980 , n4929 );
buf ( n9981 , n9980 );
not ( n9982 , n9981 );
buf ( n9983 , n4930 );
not ( n9984 , n9983 );
not ( n9985 , n9984 );
or ( n9986 , n9982 , n9985 );
not ( n9987 , n9980 );
buf ( n9988 , n9983 );
nand ( n9989 , n9987 , n9988 );
nand ( n9990 , n9986 , n9989 );
buf ( n9991 , n4931 );
not ( n9992 , n9991 );
and ( n9993 , n9990 , n9992 );
not ( n9994 , n9990 );
buf ( n9995 , n9991 );
and ( n9996 , n9994 , n9995 );
nor ( n9997 , n9993 , n9996 );
buf ( n9998 , n4932 );
nand ( n9999 , n6934 , n9998 );
buf ( n10000 , n4933 );
buf ( n10001 , n10000 );
and ( n10002 , n9999 , n10001 );
not ( n10003 , n9999 );
not ( n10004 , n10000 );
and ( n10005 , n10003 , n10004 );
nor ( n10006 , n10002 , n10005 );
xor ( n10007 , n9997 , n10006 );
buf ( n10008 , n4934 );
nand ( n10009 , n7516 , n10008 );
buf ( n10010 , n4935 );
not ( n10011 , n10010 );
and ( n10012 , n10009 , n10011 );
not ( n10013 , n10009 );
buf ( n10014 , n10010 );
and ( n10015 , n10013 , n10014 );
nor ( n10016 , n10012 , n10015 );
xnor ( n10017 , n10007 , n10016 );
buf ( n10018 , n10017 );
not ( n10019 , n10018 );
or ( n10020 , n9979 , n10019 );
buf ( n10021 , n10018 );
or ( n10022 , n10021 , n9978 );
nand ( n10023 , n10020 , n10022 );
not ( n10024 , n10023 );
buf ( n10025 , n4936 );
buf ( n10026 , n10025 );
not ( n10027 , n10026 );
not ( n10028 , n7585 );
or ( n10029 , n10027 , n10028 );
not ( n10030 , n10025 );
nand ( n10031 , n10030 , n7538 );
nand ( n10032 , n10029 , n10031 );
buf ( n10033 , n4937 );
not ( n10034 , n10033 );
and ( n10035 , n10032 , n10034 );
not ( n10036 , n10032 );
buf ( n10037 , n10033 );
and ( n10038 , n10036 , n10037 );
nor ( n10039 , n10035 , n10038 );
buf ( n10040 , n4938 );
nand ( n10041 , n8134 , n10040 );
buf ( n10042 , n4939 );
buf ( n10043 , n10042 );
and ( n10044 , n10041 , n10043 );
not ( n10045 , n10041 );
not ( n10046 , n10042 );
and ( n10047 , n10045 , n10046 );
nor ( n10048 , n10044 , n10047 );
xor ( n10049 , n10039 , n10048 );
buf ( n10050 , n4940 );
nand ( n10051 , n6934 , n10050 );
buf ( n10052 , n4941 );
not ( n10053 , n10052 );
and ( n10054 , n10051 , n10053 );
not ( n10055 , n10051 );
buf ( n10056 , n10052 );
and ( n10057 , n10055 , n10056 );
nor ( n10058 , n10054 , n10057 );
xnor ( n10059 , n10049 , n10058 );
buf ( n10060 , n10059 );
buf ( n10061 , n10060 );
not ( n10062 , n10061 );
and ( n10063 , n10024 , n10062 );
and ( n10064 , n10023 , n10061 );
nor ( n10065 , n10063 , n10064 );
not ( n10066 , n10065 );
nand ( n10067 , n9976 , n10066 );
not ( n10068 , n10067 );
buf ( n10069 , n4942 );
nand ( n10070 , n7134 , n10069 );
buf ( n10071 , n10070 );
not ( n10072 , n10071 );
buf ( n10073 , n4943 );
not ( n10074 , n10073 );
and ( n10075 , n10072 , n10074 );
and ( n10076 , n10071 , n10073 );
nor ( n10077 , n10075 , n10076 );
not ( n10078 , n10077 );
buf ( n10079 , n4944 );
buf ( n10080 , n10079 );
not ( n10081 , n10080 );
buf ( n10082 , n4945 );
not ( n10083 , n10082 );
not ( n10084 , n10083 );
or ( n10085 , n10081 , n10084 );
not ( n10086 , n10079 );
buf ( n10087 , n10082 );
nand ( n10088 , n10086 , n10087 );
nand ( n10089 , n10085 , n10088 );
buf ( n10090 , n4946 );
buf ( n10091 , n10090 );
and ( n10092 , n10089 , n10091 );
not ( n10093 , n10089 );
not ( n10094 , n10090 );
and ( n10095 , n10093 , n10094 );
nor ( n10096 , n10092 , n10095 );
buf ( n10097 , n4947 );
nand ( n10098 , n7288 , n10097 );
buf ( n10099 , n4948 );
buf ( n10100 , n10099 );
and ( n10101 , n10098 , n10100 );
not ( n10102 , n10098 );
not ( n10103 , n10099 );
and ( n10104 , n10102 , n10103 );
nor ( n10105 , n10101 , n10104 );
xor ( n10106 , n10096 , n10105 );
buf ( n10107 , n6803 );
buf ( n10108 , n4949 );
nand ( n10109 , n10107 , n10108 );
buf ( n10110 , n4950 );
buf ( n10111 , n10110 );
and ( n10112 , n10109 , n10111 );
not ( n10113 , n10109 );
not ( n10114 , n10110 );
and ( n10115 , n10113 , n10114 );
nor ( n10116 , n10112 , n10115 );
xor ( n10117 , n10106 , n10116 );
not ( n10118 , n10117 );
or ( n10119 , n10078 , n10118 );
or ( n10120 , n10117 , n10077 );
nand ( n10121 , n10119 , n10120 );
not ( n10122 , n10121 );
buf ( n10123 , n4951 );
nand ( n10124 , n6905 , n10123 );
buf ( n10125 , n4952 );
buf ( n10126 , n10125 );
and ( n10127 , n10124 , n10126 );
not ( n10128 , n10124 );
not ( n10129 , n10125 );
and ( n10130 , n10128 , n10129 );
nor ( n10131 , n10127 , n10130 );
not ( n10132 , n10131 );
buf ( n10133 , n4953 );
nand ( n10134 , n7955 , n10133 );
buf ( n10135 , n4954 );
not ( n10136 , n10135 );
and ( n10137 , n10134 , n10136 );
not ( n10138 , n10134 );
buf ( n10139 , n10135 );
and ( n10140 , n10138 , n10139 );
nor ( n10141 , n10137 , n10140 );
not ( n10142 , n10141 );
or ( n10143 , n10132 , n10142 );
or ( n10144 , n10131 , n10141 );
nand ( n10145 , n10143 , n10144 );
buf ( n10146 , n4955 );
buf ( n10147 , n10146 );
not ( n10148 , n10147 );
buf ( n10149 , n4956 );
not ( n10150 , n10149 );
not ( n10151 , n10150 );
or ( n10152 , n10148 , n10151 );
not ( n10153 , n10146 );
buf ( n10154 , n10149 );
nand ( n10155 , n10153 , n10154 );
nand ( n10156 , n10152 , n10155 );
buf ( n10157 , n4957 );
buf ( n10158 , n10157 );
and ( n10159 , n10156 , n10158 );
not ( n10160 , n10156 );
not ( n10161 , n10157 );
and ( n10162 , n10160 , n10161 );
nor ( n10163 , n10159 , n10162 );
not ( n10164 , n10163 );
and ( n10165 , n10145 , n10164 );
not ( n10166 , n10145 );
and ( n10167 , n10166 , n10163 );
nor ( n10168 , n10165 , n10167 );
buf ( n10169 , n10168 );
buf ( n10170 , n10169 );
not ( n10171 , n10170 );
and ( n10172 , n10122 , n10171 );
and ( n10173 , n10121 , n10169 );
nor ( n10174 , n10172 , n10173 );
not ( n10175 , n10174 );
not ( n10176 , n10175 );
and ( n10177 , n10068 , n10176 );
and ( n10178 , n10067 , n10175 );
nor ( n10179 , n10177 , n10178 );
and ( n10180 , n9910 , n10179 );
not ( n10181 , n9910 );
not ( n10182 , n10179 );
and ( n10183 , n10181 , n10182 );
nor ( n10184 , n10180 , n10183 );
not ( n10185 , n10184 );
buf ( n10186 , n4958 );
not ( n10187 , n10186 );
buf ( n10188 , n4959 );
not ( n10189 , n10188 );
buf ( n10190 , n4960 );
not ( n10191 , n10190 );
and ( n10192 , n10187 , n10189 , n10191 );
buf ( n10193 , n4961 );
not ( n10194 , n10193 );
and ( n10195 , n10192 , n10194 );
buf ( n10196 , n4962 );
not ( n10197 , n10196 );
buf ( n10198 , n4963 );
not ( n10199 , n10198 );
and ( n10200 , n10197 , n10199 );
buf ( n10201 , n4964 );
not ( n10202 , n10201 );
and ( n10203 , n10195 , n10200 , n10202 );
buf ( n10204 , n6815 );
buf ( n10205 , n4965 );
nand ( n10206 , n10204 , n10205 );
buf ( n10207 , n4966 );
not ( n10208 , n10207 );
and ( n10209 , n10206 , n10208 );
not ( n10210 , n10206 );
buf ( n10211 , n10207 );
and ( n10212 , n10210 , n10211 );
nor ( n10213 , n10209 , n10212 );
buf ( n10214 , n10213 );
not ( n10215 , n10214 );
buf ( n10216 , n4967 );
buf ( n10217 , n4968 );
buf ( n10218 , n10217 );
not ( n10219 , n10218 );
buf ( n10220 , n4969 );
not ( n10221 , n10220 );
not ( n10222 , n10221 );
or ( n10223 , n10219 , n10222 );
not ( n10224 , n10217 );
buf ( n10225 , n10220 );
nand ( n10226 , n10224 , n10225 );
nand ( n10227 , n10223 , n10226 );
xor ( n10228 , n10216 , n10227 );
buf ( n10229 , n4970 );
buf ( n10230 , n4971 );
not ( n10231 , n10230 );
xor ( n10232 , n10229 , n10231 );
buf ( n10233 , n4972 );
nand ( n10234 , n8740 , n10233 );
xnor ( n10235 , n10232 , n10234 );
xnor ( n10236 , n10228 , n10235 );
not ( n10237 , n10236 );
not ( n10238 , n10237 );
or ( n10239 , n10215 , n10238 );
not ( n10240 , n10214 );
nand ( n10241 , n10240 , n10236 );
nand ( n10242 , n10239 , n10241 );
buf ( n10243 , n4973 );
buf ( n10244 , n10243 );
not ( n10245 , n10244 );
buf ( n10246 , n4974 );
not ( n10247 , n10246 );
not ( n10248 , n10247 );
or ( n10249 , n10245 , n10248 );
not ( n10250 , n10243 );
buf ( n10251 , n10246 );
nand ( n10252 , n10250 , n10251 );
nand ( n10253 , n10249 , n10252 );
buf ( n10254 , n4975 );
buf ( n10255 , n10254 );
and ( n10256 , n10253 , n10255 );
not ( n10257 , n10253 );
not ( n10258 , n10254 );
and ( n10259 , n10257 , n10258 );
nor ( n10260 , n10256 , n10259 );
xor ( n10261 , n10260 , n9735 );
buf ( n10262 , n4976 );
nand ( n10263 , n7288 , n10262 );
buf ( n10264 , n4977 );
buf ( n10265 , n10264 );
and ( n10266 , n10263 , n10265 );
not ( n10267 , n10263 );
not ( n10268 , n10264 );
and ( n10269 , n10267 , n10268 );
nor ( n10270 , n10266 , n10269 );
not ( n10271 , n10270 );
xnor ( n10272 , n10261 , n10271 );
not ( n10273 , n10272 );
not ( n10274 , n10273 );
and ( n10275 , n10242 , n10274 );
not ( n10276 , n10242 );
xor ( n10277 , n10260 , n10270 );
xor ( n10278 , n10277 , n9736 );
buf ( n10279 , n10278 );
and ( n10280 , n10276 , n10279 );
nor ( n10281 , n10275 , n10280 );
xor ( n10282 , n10203 , n10281 );
buf ( n10283 , n4978 );
nand ( n10284 , n7921 , n10283 );
buf ( n10285 , n4979 );
not ( n10286 , n10285 );
and ( n10287 , n10284 , n10286 );
not ( n10288 , n10284 );
buf ( n10289 , n10285 );
and ( n10290 , n10288 , n10289 );
nor ( n10291 , n10287 , n10290 );
not ( n10292 , n10291 );
buf ( n10293 , n4980 );
buf ( n10294 , n10293 );
not ( n10295 , n10294 );
buf ( n10296 , n4981 );
not ( n10297 , n10296 );
not ( n10298 , n10297 );
or ( n10299 , n10295 , n10298 );
not ( n10300 , n10293 );
buf ( n10301 , n10296 );
nand ( n10302 , n10300 , n10301 );
nand ( n10303 , n10299 , n10302 );
buf ( n10304 , n4982 );
not ( n10305 , n10304 );
and ( n10306 , n10303 , n10305 );
not ( n10307 , n10303 );
buf ( n10308 , n10304 );
and ( n10309 , n10307 , n10308 );
nor ( n10310 , n10306 , n10309 );
buf ( n10311 , n4983 );
nand ( n10312 , n7133 , n10311 );
buf ( n10313 , n4984 );
buf ( n10314 , n10313 );
and ( n10315 , n10312 , n10314 );
not ( n10316 , n10312 );
not ( n10317 , n10313 );
and ( n10318 , n10316 , n10317 );
nor ( n10319 , n10315 , n10318 );
xor ( n10320 , n10310 , n10319 );
buf ( n10321 , n4985 );
nand ( n10322 , n7750 , n10321 );
buf ( n10323 , n4986 );
not ( n10324 , n10323 );
and ( n10325 , n10322 , n10324 );
not ( n10326 , n10322 );
buf ( n10327 , n10323 );
and ( n10328 , n10326 , n10327 );
nor ( n10329 , n10325 , n10328 );
xor ( n10330 , n10320 , n10329 );
not ( n10331 , n10330 );
not ( n10332 , n10331 );
or ( n10333 , n10292 , n10332 );
not ( n10334 , n10291 );
nand ( n10335 , n10334 , n10330 );
nand ( n10336 , n10333 , n10335 );
buf ( n10337 , n4987 );
buf ( n10338 , n10337 );
not ( n10339 , n10338 );
buf ( n10340 , n4988 );
not ( n10341 , n10340 );
not ( n10342 , n10341 );
or ( n10343 , n10339 , n10342 );
not ( n10344 , n10337 );
buf ( n10345 , n10340 );
nand ( n10346 , n10344 , n10345 );
nand ( n10347 , n10343 , n10346 );
buf ( n10348 , n4989 );
buf ( n10349 , n10348 );
and ( n10350 , n10347 , n10349 );
not ( n10351 , n10347 );
not ( n10352 , n10348 );
and ( n10353 , n10351 , n10352 );
nor ( n10354 , n10350 , n10353 );
buf ( n10355 , n4990 );
nand ( n10356 , n6863 , n10355 );
buf ( n10357 , n4991 );
buf ( n10358 , n10357 );
and ( n10359 , n10356 , n10358 );
not ( n10360 , n10356 );
not ( n10361 , n10357 );
and ( n10362 , n10360 , n10361 );
nor ( n10363 , n10359 , n10362 );
xor ( n10364 , n10354 , n10363 );
buf ( n10365 , n4992 );
nand ( n10366 , n9257 , n10365 );
buf ( n10367 , n4993 );
not ( n10368 , n10367 );
and ( n10369 , n10366 , n10368 );
not ( n10370 , n10366 );
buf ( n10371 , n10367 );
and ( n10372 , n10370 , n10371 );
nor ( n10373 , n10369 , n10372 );
xnor ( n10374 , n10364 , n10373 );
not ( n10375 , n10374 );
buf ( n10376 , n10375 );
not ( n10377 , n10376 );
and ( n10378 , n10336 , n10377 );
not ( n10379 , n10336 );
and ( n10380 , n10379 , n10376 );
nor ( n10381 , n10378 , n10380 );
not ( n10382 , n8858 );
buf ( n10383 , n4994 );
not ( n10384 , n10383 );
not ( n10385 , n10384 );
buf ( n10386 , n4995 );
not ( n10387 , n10386 );
and ( n10388 , n10385 , n10387 );
and ( n10389 , n10386 , n10384 );
nor ( n10390 , n10388 , n10389 );
not ( n10391 , n10390 );
or ( n10392 , n10382 , n10391 );
or ( n10393 , n10390 , n8858 );
nand ( n10394 , n10392 , n10393 );
not ( n10395 , n10394 );
buf ( n10396 , n4996 );
not ( n10397 , n10396 );
buf ( n10398 , n4997 );
nand ( n10399 , n7133 , n10398 );
buf ( n10400 , n4998 );
buf ( n10401 , n10400 );
and ( n10402 , n10399 , n10401 );
not ( n10403 , n10399 );
not ( n10404 , n10400 );
and ( n10405 , n10403 , n10404 );
nor ( n10406 , n10402 , n10405 );
xor ( n10407 , n10397 , n10406 );
buf ( n10408 , n4999 );
nand ( n10409 , n7955 , n10408 );
buf ( n10410 , n5000 );
buf ( n10411 , n10410 );
and ( n10412 , n10409 , n10411 );
not ( n10413 , n10409 );
not ( n10414 , n10410 );
and ( n10415 , n10413 , n10414 );
nor ( n10416 , n10412 , n10415 );
xnor ( n10417 , n10407 , n10416 );
not ( n10418 , n10417 );
not ( n10419 , n10418 );
or ( n10420 , n10395 , n10419 );
or ( n10421 , n10418 , n10394 );
nand ( n10422 , n10420 , n10421 );
not ( n10423 , n10422 );
buf ( n10424 , n5001 );
buf ( n10425 , n10424 );
not ( n10426 , n10425 );
buf ( n10427 , n5002 );
not ( n10428 , n10427 );
not ( n10429 , n10428 );
or ( n10430 , n10426 , n10429 );
not ( n10431 , n10424 );
buf ( n10432 , n10427 );
nand ( n10433 , n10431 , n10432 );
nand ( n10434 , n10430 , n10433 );
buf ( n10435 , n5003 );
not ( n10436 , n10435 );
and ( n10437 , n10434 , n10436 );
not ( n10438 , n10434 );
buf ( n10439 , n10435 );
and ( n10440 , n10438 , n10439 );
nor ( n10441 , n10437 , n10440 );
not ( n10442 , n10441 );
buf ( n10443 , n5004 );
nand ( n10444 , n6660 , n10443 );
buf ( n10445 , n5005 );
buf ( n10446 , n10445 );
and ( n10447 , n10444 , n10446 );
not ( n10448 , n10444 );
not ( n10449 , n10445 );
and ( n10450 , n10448 , n10449 );
nor ( n10451 , n10447 , n10450 );
xor ( n10452 , n10442 , n10451 );
buf ( n10453 , n5006 );
nand ( n10454 , n7617 , n10453 );
buf ( n10455 , n5007 );
buf ( n10456 , n10455 );
and ( n10457 , n10454 , n10456 );
not ( n10458 , n10454 );
not ( n10459 , n10455 );
and ( n10460 , n10458 , n10459 );
nor ( n10461 , n10457 , n10460 );
xnor ( n10462 , n10452 , n10461 );
buf ( n10463 , n10462 );
not ( n10464 , n10463 );
and ( n10465 , n10423 , n10464 );
and ( n10466 , n10422 , n10463 );
nor ( n10467 , n10465 , n10466 );
nor ( n10468 , n10381 , n10467 );
xnor ( n10469 , n10282 , n10468 );
not ( n10470 , n10469 );
buf ( n10471 , n5008 );
not ( n10472 , n10471 );
not ( n10473 , n10472 );
buf ( n10474 , n5009 );
buf ( n10475 , n5010 );
buf ( n10476 , n10475 );
not ( n10477 , n10476 );
buf ( n10478 , n5011 );
not ( n10479 , n10478 );
not ( n10480 , n10479 );
or ( n10481 , n10477 , n10480 );
not ( n10482 , n10475 );
buf ( n10483 , n10478 );
nand ( n10484 , n10482 , n10483 );
nand ( n10485 , n10481 , n10484 );
not ( n10486 , n10485 );
xor ( n10487 , n10474 , n10486 );
buf ( n10488 , n5012 );
buf ( n10489 , n5013 );
xor ( n10490 , n10488 , n10489 );
buf ( n10491 , n5014 );
nand ( n10492 , n8821 , n10491 );
xnor ( n10493 , n10490 , n10492 );
xnor ( n10494 , n10487 , n10493 );
not ( n10495 , n10494 );
or ( n10496 , n10473 , n10495 );
not ( n10497 , n10472 );
not ( n10498 , n10494 );
nand ( n10499 , n10497 , n10498 );
nand ( n10500 , n10496 , n10499 );
buf ( n10501 , n5015 );
buf ( n10502 , n10501 );
not ( n10503 , n10502 );
buf ( n10504 , n5016 );
not ( n10505 , n10504 );
not ( n10506 , n10505 );
or ( n10507 , n10503 , n10506 );
not ( n10508 , n10501 );
buf ( n10509 , n10504 );
nand ( n10510 , n10508 , n10509 );
nand ( n10511 , n10507 , n10510 );
buf ( n10512 , n5017 );
not ( n10513 , n10512 );
and ( n10514 , n10511 , n10513 );
not ( n10515 , n10511 );
buf ( n10516 , n10512 );
and ( n10517 , n10515 , n10516 );
nor ( n10518 , n10514 , n10517 );
buf ( n10519 , n5018 );
nand ( n10520 , n7126 , n10519 );
buf ( n10521 , n5019 );
buf ( n10522 , n10521 );
and ( n10523 , n10520 , n10522 );
not ( n10524 , n10520 );
not ( n10525 , n10521 );
and ( n10526 , n10524 , n10525 );
nor ( n10527 , n10523 , n10526 );
xor ( n10528 , n10518 , n10527 );
buf ( n10529 , n5020 );
nand ( n10530 , n8135 , n10529 );
buf ( n10531 , n5021 );
not ( n10532 , n10531 );
and ( n10533 , n10530 , n10532 );
not ( n10534 , n10530 );
buf ( n10535 , n10531 );
and ( n10536 , n10534 , n10535 );
nor ( n10537 , n10533 , n10536 );
xnor ( n10538 , n10528 , n10537 );
buf ( n10539 , n10538 );
buf ( n10540 , n10539 );
and ( n10541 , n10500 , n10540 );
not ( n10542 , n10500 );
not ( n10543 , n10539 );
and ( n10544 , n10542 , n10543 );
nor ( n10545 , n10541 , n10544 );
not ( n10546 , n10545 );
buf ( n10547 , n5022 );
not ( n10548 , n10547 );
buf ( n10549 , n5023 );
buf ( n10550 , n10549 );
not ( n10551 , n10550 );
buf ( n10552 , n5024 );
not ( n10553 , n10552 );
not ( n10554 , n10553 );
or ( n10555 , n10551 , n10554 );
not ( n10556 , n10549 );
buf ( n10557 , n10552 );
nand ( n10558 , n10556 , n10557 );
nand ( n10559 , n10555 , n10558 );
buf ( n10560 , n5025 );
not ( n10561 , n10560 );
and ( n10562 , n10559 , n10561 );
not ( n10563 , n10559 );
buf ( n10564 , n10560 );
and ( n10565 , n10563 , n10564 );
nor ( n10566 , n10562 , n10565 );
buf ( n10567 , n5026 );
nand ( n10568 , n7471 , n10567 );
buf ( n10569 , n5027 );
buf ( n10570 , n10569 );
and ( n10571 , n10568 , n10570 );
not ( n10572 , n10568 );
not ( n10573 , n10569 );
and ( n10574 , n10572 , n10573 );
nor ( n10575 , n10571 , n10574 );
xor ( n10576 , n10566 , n10575 );
buf ( n10577 , n6803 );
buf ( n10578 , n5028 );
nand ( n10579 , n10577 , n10578 );
buf ( n10580 , n5029 );
not ( n10581 , n10580 );
and ( n10582 , n10579 , n10581 );
not ( n10583 , n10579 );
buf ( n10584 , n10580 );
and ( n10585 , n10583 , n10584 );
nor ( n10586 , n10582 , n10585 );
xnor ( n10587 , n10576 , n10586 );
not ( n10588 , n10587 );
not ( n10589 , n10588 );
not ( n10590 , n10589 );
or ( n10591 , n10548 , n10590 );
not ( n10592 , n10547 );
nand ( n10593 , n10592 , n10588 );
nand ( n10594 , n10591 , n10593 );
buf ( n10595 , n5030 );
nand ( n10596 , n8923 , n10595 );
buf ( n10597 , n5031 );
buf ( n10598 , n10597 );
and ( n10599 , n10596 , n10598 );
not ( n10600 , n10596 );
not ( n10601 , n10597 );
and ( n10602 , n10600 , n10601 );
nor ( n10603 , n10599 , n10602 );
not ( n10604 , n10603 );
buf ( n10605 , n5032 );
nand ( n10606 , n7477 , n10605 );
buf ( n10607 , n5033 );
not ( n10608 , n10607 );
and ( n10609 , n10606 , n10608 );
not ( n10610 , n10606 );
buf ( n10611 , n10607 );
and ( n10612 , n10610 , n10611 );
nor ( n10613 , n10609 , n10612 );
not ( n10614 , n10613 );
or ( n10615 , n10604 , n10614 );
or ( n10616 , n10603 , n10613 );
nand ( n10617 , n10615 , n10616 );
buf ( n10618 , n5034 );
buf ( n10619 , n10618 );
not ( n10620 , n10619 );
buf ( n10621 , n5035 );
not ( n10622 , n10621 );
not ( n10623 , n10622 );
or ( n10624 , n10620 , n10623 );
not ( n10625 , n10618 );
buf ( n10626 , n10621 );
nand ( n10627 , n10625 , n10626 );
nand ( n10628 , n10624 , n10627 );
buf ( n10629 , n5036 );
not ( n10630 , n10629 );
and ( n10631 , n10628 , n10630 );
not ( n10632 , n10628 );
buf ( n10633 , n10629 );
and ( n10634 , n10632 , n10633 );
nor ( n10635 , n10631 , n10634 );
not ( n10636 , n10635 );
and ( n10637 , n10617 , n10636 );
not ( n10638 , n10617 );
and ( n10639 , n10638 , n10635 );
nor ( n10640 , n10637 , n10639 );
not ( n10641 , n10640 );
and ( n10642 , n10594 , n10641 );
not ( n10643 , n10594 );
not ( n10644 , n10641 );
and ( n10645 , n10643 , n10644 );
nor ( n10646 , n10642 , n10645 );
nand ( n10647 , n10546 , n10646 );
not ( n10648 , n10647 );
buf ( n10649 , n5037 );
nand ( n10650 , n7413 , n10649 );
buf ( n10651 , n5038 );
buf ( n10652 , n10651 );
and ( n10653 , n10650 , n10652 );
not ( n10654 , n10650 );
not ( n10655 , n10651 );
and ( n10656 , n10654 , n10655 );
nor ( n10657 , n10653 , n10656 );
not ( n10658 , n10657 );
buf ( n10659 , n5039 );
buf ( n10660 , n10659 );
not ( n10661 , n10660 );
buf ( n10662 , n5040 );
not ( n10663 , n10662 );
not ( n10664 , n10663 );
or ( n10665 , n10661 , n10664 );
not ( n10666 , n10659 );
buf ( n10667 , n10662 );
nand ( n10668 , n10666 , n10667 );
nand ( n10669 , n10665 , n10668 );
buf ( n10670 , n5041 );
buf ( n10671 , n10670 );
and ( n10672 , n10669 , n10671 );
not ( n10673 , n10669 );
not ( n10674 , n10670 );
and ( n10675 , n10673 , n10674 );
nor ( n10676 , n10672 , n10675 );
buf ( n10677 , n5042 );
nand ( n10678 , n7183 , n10677 );
buf ( n10679 , n5043 );
not ( n10680 , n10679 );
and ( n10681 , n10678 , n10680 );
not ( n10682 , n10678 );
buf ( n10683 , n10679 );
and ( n10684 , n10682 , n10683 );
nor ( n10685 , n10681 , n10684 );
xor ( n10686 , n10676 , n10685 );
buf ( n10687 , n5044 );
nand ( n10688 , n6608 , n10687 );
buf ( n10689 , n5045 );
not ( n10690 , n10689 );
and ( n10691 , n10688 , n10690 );
not ( n10692 , n10688 );
buf ( n10693 , n10689 );
and ( n10694 , n10692 , n10693 );
nor ( n10695 , n10691 , n10694 );
xnor ( n10696 , n10686 , n10695 );
not ( n10697 , n10696 );
not ( n10698 , n10697 );
or ( n10699 , n10658 , n10698 );
or ( n10700 , n10697 , n10657 );
nand ( n10701 , n10699 , n10700 );
not ( n10702 , n10701 );
not ( n10703 , n10702 );
buf ( n10704 , n5046 );
not ( n10705 , n10704 );
buf ( n10706 , n5047 );
buf ( n10707 , n10706 );
not ( n10708 , n10707 );
buf ( n10709 , n5048 );
not ( n10710 , n10709 );
not ( n10711 , n10710 );
or ( n10712 , n10708 , n10711 );
not ( n10713 , n10706 );
buf ( n10714 , n10709 );
nand ( n10715 , n10713 , n10714 );
nand ( n10716 , n10712 , n10715 );
xor ( n10717 , n10705 , n10716 );
buf ( n10718 , n5049 );
not ( n10719 , n10718 );
buf ( n10720 , n5050 );
nand ( n10721 , n6660 , n10720 );
buf ( n10722 , n5051 );
buf ( n10723 , n10722 );
and ( n10724 , n10721 , n10723 );
not ( n10725 , n10721 );
not ( n10726 , n10722 );
and ( n10727 , n10725 , n10726 );
nor ( n10728 , n10724 , n10727 );
not ( n10729 , n10728 );
or ( n10730 , n10719 , n10729 );
or ( n10731 , n10728 , n10718 );
nand ( n10732 , n10730 , n10731 );
xnor ( n10733 , n10717 , n10732 );
buf ( n10734 , n10733 );
not ( n10735 , n10734 );
or ( n10736 , n10703 , n10735 );
buf ( n10737 , n10704 );
xor ( n10738 , n10737 , n10716 );
xnor ( n10739 , n10738 , n10732 );
nand ( n10740 , n10739 , n10701 );
nand ( n10741 , n10736 , n10740 );
buf ( n10742 , n10741 );
not ( n10743 , n10742 );
and ( n10744 , n10648 , n10743 );
and ( n10745 , n10647 , n10742 );
nor ( n10746 , n10744 , n10745 );
not ( n10747 , n10746 );
and ( n10748 , n10470 , n10747 );
and ( n10749 , n10469 , n10746 );
nor ( n10750 , n10748 , n10749 );
and ( n10751 , n10185 , n10750 );
not ( n10752 , n10185 );
not ( n10753 , n10750 );
and ( n10754 , n10752 , n10753 );
nor ( n10755 , n10751 , n10754 );
not ( n10756 , n10755 );
or ( n10757 , n9638 , n10756 );
not ( n10758 , n9637 );
not ( n10759 , n10750 );
not ( n10760 , n10184 );
not ( n10761 , n10760 );
or ( n10762 , n10759 , n10761 );
not ( n10763 , n10750 );
nand ( n10764 , n10763 , n10184 );
nand ( n10765 , n10762 , n10764 );
nand ( n10766 , n10758 , n10765 );
nand ( n10767 , n10757 , n10766 );
buf ( n10768 , n5052 );
buf ( n10769 , n10768 );
not ( n10770 , n10769 );
buf ( n10771 , n5053 );
buf ( n10772 , n10771 );
not ( n10773 , n10772 );
buf ( n10774 , n5054 );
not ( n10775 , n10774 );
not ( n10776 , n10775 );
or ( n10777 , n10773 , n10776 );
not ( n10778 , n10771 );
buf ( n10779 , n10774 );
nand ( n10780 , n10778 , n10779 );
nand ( n10781 , n10777 , n10780 );
buf ( n10782 , n5055 );
buf ( n10783 , n10782 );
and ( n10784 , n10781 , n10783 );
not ( n10785 , n10781 );
not ( n10786 , n10782 );
and ( n10787 , n10785 , n10786 );
nor ( n10788 , n10784 , n10787 );
buf ( n10789 , n5056 );
nand ( n10790 , n8923 , n10789 );
buf ( n10791 , n5057 );
buf ( n10792 , n10791 );
and ( n10793 , n10790 , n10792 );
not ( n10794 , n10790 );
not ( n10795 , n10791 );
and ( n10796 , n10794 , n10795 );
nor ( n10797 , n10793 , n10796 );
xor ( n10798 , n10788 , n10797 );
buf ( n10799 , n5058 );
nand ( n10800 , n7184 , n10799 );
buf ( n10801 , n5059 );
not ( n10802 , n10801 );
and ( n10803 , n10800 , n10802 );
not ( n10804 , n10800 );
buf ( n10805 , n10801 );
and ( n10806 , n10804 , n10805 );
nor ( n10807 , n10803 , n10806 );
xnor ( n10808 , n10798 , n10807 );
buf ( n10809 , n10808 );
not ( n10810 , n10809 );
not ( n10811 , n10810 );
or ( n10812 , n10770 , n10811 );
or ( n10813 , n10810 , n10769 );
nand ( n10814 , n10812 , n10813 );
buf ( n10815 , n5060 );
buf ( n10816 , n10815 );
buf ( n10817 , n5061 );
buf ( n10818 , n10817 );
not ( n10819 , n10818 );
buf ( n10820 , n5062 );
not ( n10821 , n10820 );
not ( n10822 , n10821 );
or ( n10823 , n10819 , n10822 );
not ( n10824 , n10817 );
buf ( n10825 , n10820 );
nand ( n10826 , n10824 , n10825 );
nand ( n10827 , n10823 , n10826 );
xor ( n10828 , n10816 , n10827 );
buf ( n10829 , n5063 );
nand ( n10830 , n8387 , n10829 );
buf ( n10831 , n5064 );
buf ( n10832 , n10831 );
and ( n10833 , n10830 , n10832 );
not ( n10834 , n10830 );
not ( n10835 , n10831 );
and ( n10836 , n10834 , n10835 );
nor ( n10837 , n10833 , n10836 );
not ( n10838 , n10837 );
buf ( n10839 , n5065 );
not ( n10840 , n10839 );
and ( n10841 , n10838 , n10840 );
and ( n10842 , n10837 , n10839 );
nor ( n10843 , n10841 , n10842 );
xnor ( n10844 , n10828 , n10843 );
not ( n10845 , n10844 );
not ( n10846 , n10845 );
and ( n10847 , n10814 , n10846 );
not ( n10848 , n10814 );
and ( n10849 , n10848 , n10845 );
nor ( n10850 , n10847 , n10849 );
buf ( n10851 , n5066 );
buf ( n10852 , n10851 );
not ( n10853 , n10852 );
buf ( n10854 , n9219 );
not ( n10855 , n10854 );
or ( n10856 , n10853 , n10855 );
or ( n10857 , n9221 , n10852 );
nand ( n10858 , n10856 , n10857 );
not ( n10859 , n6581 );
buf ( n10860 , n5067 );
not ( n10861 , n10860 );
not ( n10862 , n10861 );
or ( n10863 , n10859 , n10862 );
not ( n10864 , n6580 );
buf ( n10865 , n10860 );
nand ( n10866 , n10864 , n10865 );
nand ( n10867 , n10863 , n10866 );
buf ( n10868 , n5068 );
not ( n10869 , n10868 );
and ( n10870 , n10867 , n10869 );
not ( n10871 , n10867 );
buf ( n10872 , n10868 );
and ( n10873 , n10871 , n10872 );
nor ( n10874 , n10870 , n10873 );
buf ( n10875 , n5069 );
nand ( n10876 , n7230 , n10875 );
buf ( n10877 , n5070 );
buf ( n10878 , n10877 );
and ( n10879 , n10876 , n10878 );
not ( n10880 , n10876 );
not ( n10881 , n10877 );
and ( n10882 , n10880 , n10881 );
nor ( n10883 , n10879 , n10882 );
xor ( n10884 , n10874 , n10883 );
buf ( n10885 , n5071 );
nand ( n10886 , n7356 , n10885 );
buf ( n10887 , n5072 );
buf ( n10888 , n10887 );
and ( n10889 , n10886 , n10888 );
not ( n10890 , n10886 );
not ( n10891 , n10887 );
and ( n10892 , n10890 , n10891 );
nor ( n10893 , n10889 , n10892 );
xnor ( n10894 , n10884 , n10893 );
not ( n10895 , n10894 );
buf ( n10896 , n10895 );
xor ( n10897 , n10858 , n10896 );
nand ( n10898 , n10850 , n10897 );
not ( n10899 , n10898 );
not ( n10900 , n7548 );
not ( n10901 , n6772 );
or ( n10902 , n10900 , n10901 );
not ( n10903 , n6773 );
nand ( n10904 , n10903 , n7544 );
nand ( n10905 , n10902 , n10904 );
not ( n10906 , n10905 );
buf ( n10907 , n5073 );
buf ( n10908 , n10907 );
not ( n10909 , n10908 );
not ( n10910 , n9128 );
or ( n10911 , n10909 , n10910 );
not ( n10912 , n10907 );
nand ( n10913 , n10912 , n9084 );
nand ( n10914 , n10911 , n10913 );
buf ( n10915 , n5074 );
not ( n10916 , n10915 );
and ( n10917 , n10914 , n10916 );
not ( n10918 , n10914 );
buf ( n10919 , n10915 );
and ( n10920 , n10918 , n10919 );
nor ( n10921 , n10917 , n10920 );
buf ( n10922 , n5075 );
nand ( n10923 , n7471 , n10922 );
buf ( n10924 , n5076 );
buf ( n10925 , n10924 );
and ( n10926 , n10923 , n10925 );
not ( n10927 , n10923 );
not ( n10928 , n10924 );
and ( n10929 , n10927 , n10928 );
nor ( n10930 , n10926 , n10929 );
xor ( n10931 , n10921 , n10930 );
buf ( n10932 , n5077 );
nand ( n10933 , n7196 , n10932 );
buf ( n10934 , n5078 );
buf ( n10935 , n10934 );
and ( n10936 , n10933 , n10935 );
not ( n10937 , n10933 );
not ( n10938 , n10934 );
and ( n10939 , n10937 , n10938 );
nor ( n10940 , n10936 , n10939 );
xnor ( n10941 , n10931 , n10940 );
buf ( n10942 , n10941 );
not ( n10943 , n10942 );
not ( n10944 , n10943 );
and ( n10945 , n10906 , n10944 );
and ( n10946 , n10905 , n10943 );
nor ( n10947 , n10945 , n10946 );
not ( n10948 , n10947 );
not ( n10949 , n10948 );
and ( n10950 , n10899 , n10949 );
and ( n10951 , n10898 , n10948 );
nor ( n10952 , n10950 , n10951 );
not ( n10953 , n10952 );
buf ( n10954 , n5079 );
buf ( n10955 , n10954 );
not ( n10956 , n10955 );
buf ( n10957 , n5080 );
buf ( n10958 , n10957 );
not ( n10959 , n10958 );
buf ( n10960 , n5081 );
not ( n10961 , n10960 );
not ( n10962 , n10961 );
or ( n10963 , n10959 , n10962 );
not ( n10964 , n10957 );
buf ( n10965 , n10960 );
nand ( n10966 , n10964 , n10965 );
nand ( n10967 , n10963 , n10966 );
buf ( n10968 , n5082 );
not ( n10969 , n10968 );
and ( n10970 , n10967 , n10969 );
not ( n10971 , n10967 );
buf ( n10972 , n10968 );
and ( n10973 , n10971 , n10972 );
nor ( n10974 , n10970 , n10973 );
buf ( n10975 , n5083 );
nand ( n10976 , n7126 , n10975 );
buf ( n10977 , n5084 );
buf ( n10978 , n10977 );
and ( n10979 , n10976 , n10978 );
not ( n10980 , n10976 );
not ( n10981 , n10977 );
and ( n10982 , n10980 , n10981 );
nor ( n10983 , n10979 , n10982 );
xor ( n10984 , n10974 , n10983 );
buf ( n10985 , n5085 );
nand ( n10986 , n7082 , n10985 );
buf ( n10987 , n5086 );
not ( n10988 , n10987 );
and ( n10989 , n10986 , n10988 );
not ( n10990 , n10986 );
buf ( n10991 , n10987 );
and ( n10992 , n10990 , n10991 );
nor ( n10993 , n10989 , n10992 );
xnor ( n10994 , n10984 , n10993 );
buf ( n10995 , n10994 );
not ( n10996 , n10995 );
or ( n10997 , n10956 , n10996 );
not ( n10998 , n10983 );
not ( n10999 , n10993 );
or ( n11000 , n10998 , n10999 );
or ( n11001 , n10983 , n10993 );
nand ( n11002 , n11000 , n11001 );
not ( n11003 , n10974 );
and ( n11004 , n11002 , n11003 );
not ( n11005 , n11002 );
and ( n11006 , n11005 , n10974 );
nor ( n11007 , n11004 , n11006 );
not ( n11008 , n11007 );
not ( n11009 , n11008 );
not ( n11010 , n10954 );
nand ( n11011 , n11009 , n11010 );
nand ( n11012 , n10997 , n11011 );
not ( n11013 , n10021 );
and ( n11014 , n11012 , n11013 );
not ( n11015 , n11012 );
and ( n11016 , n11015 , n10021 );
nor ( n11017 , n11014 , n11016 );
not ( n11018 , n11017 );
buf ( n11019 , n5087 );
buf ( n11020 , n11019 );
buf ( n11021 , n5088 );
buf ( n11022 , n11021 );
not ( n11023 , n11022 );
buf ( n11024 , n5089 );
not ( n11025 , n11024 );
not ( n11026 , n11025 );
or ( n11027 , n11023 , n11026 );
not ( n11028 , n11021 );
buf ( n11029 , n11024 );
nand ( n11030 , n11028 , n11029 );
nand ( n11031 , n11027 , n11030 );
buf ( n11032 , n5090 );
buf ( n11033 , n11032 );
and ( n11034 , n11031 , n11033 );
not ( n11035 , n11031 );
not ( n11036 , n11032 );
and ( n11037 , n11035 , n11036 );
nor ( n11038 , n11034 , n11037 );
buf ( n11039 , n5091 );
nand ( n11040 , n6607 , n11039 );
buf ( n11041 , n5092 );
buf ( n11042 , n11041 );
and ( n11043 , n11040 , n11042 );
not ( n11044 , n11040 );
not ( n11045 , n11041 );
and ( n11046 , n11044 , n11045 );
nor ( n11047 , n11043 , n11046 );
xor ( n11048 , n11038 , n11047 );
buf ( n11049 , n5093 );
nand ( n11050 , n7442 , n11049 );
buf ( n11051 , n5094 );
not ( n11052 , n11051 );
and ( n11053 , n11050 , n11052 );
not ( n11054 , n11050 );
buf ( n11055 , n11051 );
and ( n11056 , n11054 , n11055 );
nor ( n11057 , n11053 , n11056 );
xnor ( n11058 , n11048 , n11057 );
buf ( n11059 , n11058 );
xor ( n11060 , n11020 , n11059 );
not ( n11061 , n8612 );
xnor ( n11062 , n11060 , n11061 );
nand ( n11063 , n11018 , n11062 );
buf ( n11064 , n5095 );
buf ( n11065 , n11064 );
not ( n11066 , n11065 );
buf ( n11067 , n5096 );
buf ( n11068 , n11067 );
not ( n11069 , n11068 );
buf ( n11070 , n5097 );
not ( n11071 , n11070 );
not ( n11072 , n11071 );
or ( n11073 , n11069 , n11072 );
not ( n11074 , n11067 );
buf ( n11075 , n11070 );
nand ( n11076 , n11074 , n11075 );
nand ( n11077 , n11073 , n11076 );
buf ( n11078 , n5098 );
not ( n11079 , n11078 );
and ( n11080 , n11077 , n11079 );
not ( n11081 , n11077 );
buf ( n11082 , n11078 );
and ( n11083 , n11081 , n11082 );
nor ( n11084 , n11080 , n11083 );
buf ( n11085 , n5099 );
nand ( n11086 , n6803 , n11085 );
buf ( n11087 , n5100 );
buf ( n11088 , n11087 );
and ( n11089 , n11086 , n11088 );
not ( n11090 , n11086 );
not ( n11091 , n11087 );
and ( n11092 , n11090 , n11091 );
nor ( n11093 , n11089 , n11092 );
xor ( n11094 , n11084 , n11093 );
buf ( n11095 , n5101 );
nand ( n11096 , n7184 , n11095 );
buf ( n11097 , n5102 );
not ( n11098 , n11097 );
and ( n11099 , n11096 , n11098 );
not ( n11100 , n11096 );
buf ( n11101 , n11097 );
and ( n11102 , n11100 , n11101 );
nor ( n11103 , n11099 , n11102 );
xnor ( n11104 , n11094 , n11103 );
not ( n11105 , n11104 );
or ( n11106 , n11066 , n11105 );
not ( n11107 , n11084 );
xor ( n11108 , n11107 , n11093 );
xnor ( n11109 , n11108 , n11103 );
not ( n11110 , n11064 );
nand ( n11111 , n11109 , n11110 );
nand ( n11112 , n11106 , n11111 );
not ( n11113 , n11112 );
buf ( n11114 , n5103 );
not ( n11115 , n11114 );
buf ( n11116 , n5104 );
not ( n11117 , n11116 );
buf ( n11118 , n5105 );
buf ( n11119 , n11118 );
nand ( n11120 , n11117 , n11119 );
not ( n11121 , n11118 );
buf ( n11122 , n11116 );
nand ( n11123 , n11121 , n11122 );
and ( n11124 , n11120 , n11123 );
xor ( n11125 , n11115 , n11124 );
buf ( n11126 , n5106 );
xor ( n11127 , n11126 , n10073 );
xnor ( n11128 , n11127 , n10070 );
xnor ( n11129 , n11125 , n11128 );
buf ( n11130 , n11129 );
not ( n11131 , n11130 );
or ( n11132 , n11113 , n11131 );
or ( n11133 , n11130 , n11112 );
nand ( n11134 , n11132 , n11133 );
not ( n11135 , n11134 );
and ( n11136 , n11063 , n11135 );
not ( n11137 , n11063 );
and ( n11138 , n11137 , n11134 );
nor ( n11139 , n11136 , n11138 );
not ( n11140 , n11139 );
or ( n11141 , n10953 , n11140 );
or ( n11142 , n11139 , n10952 );
nand ( n11143 , n11141 , n11142 );
not ( n11144 , n11143 );
not ( n11145 , n8810 );
buf ( n11146 , n5107 );
buf ( n11147 , n5108 );
not ( n11148 , n11147 );
buf ( n11149 , n5109 );
buf ( n11150 , n11149 );
and ( n11151 , n11148 , n11150 );
not ( n11152 , n11148 );
not ( n11153 , n11149 );
and ( n11154 , n11152 , n11153 );
nor ( n11155 , n11151 , n11154 );
xor ( n11156 , n11146 , n11155 );
buf ( n11157 , n5110 );
nand ( n11158 , n7477 , n11157 );
not ( n11159 , n11158 );
buf ( n11160 , n5111 );
not ( n11161 , n11160 );
and ( n11162 , n11159 , n11161 );
nand ( n11163 , n7082 , n11157 );
and ( n11164 , n11163 , n11160 );
nor ( n11165 , n11162 , n11164 );
not ( n11166 , n11165 );
buf ( n11167 , n5112 );
not ( n11168 , n11167 );
and ( n11169 , n11166 , n11168 );
and ( n11170 , n11165 , n11167 );
nor ( n11171 , n11169 , n11170 );
xnor ( n11172 , n11156 , n11171 );
not ( n11173 , n11172 );
not ( n11174 , n11173 );
or ( n11175 , n11145 , n11174 );
buf ( n11176 , n11172 );
not ( n11177 , n11176 );
or ( n11178 , n11177 , n8810 );
nand ( n11179 , n11175 , n11178 );
not ( n11180 , n10390 );
not ( n11181 , n11180 );
not ( n11182 , n10418 );
or ( n11183 , n11181 , n11182 );
nand ( n11184 , n10417 , n10390 );
nand ( n11185 , n11183 , n11184 );
buf ( n11186 , n11185 );
not ( n11187 , n11186 );
and ( n11188 , n11179 , n11187 );
not ( n11189 , n11179 );
and ( n11190 , n11189 , n11186 );
nor ( n11191 , n11188 , n11190 );
buf ( n11192 , n5113 );
buf ( n11193 , n5114 );
buf ( n11194 , n11193 );
not ( n11195 , n11194 );
buf ( n11196 , n5115 );
not ( n11197 , n11196 );
not ( n11198 , n11197 );
or ( n11199 , n11195 , n11198 );
not ( n11200 , n11193 );
buf ( n11201 , n11196 );
nand ( n11202 , n11200 , n11201 );
nand ( n11203 , n11199 , n11202 );
xor ( n11204 , n11192 , n11203 );
buf ( n11205 , n5116 );
nand ( n11206 , n7093 , n11205 );
buf ( n11207 , n5117 );
buf ( n11208 , n11207 );
and ( n11209 , n11206 , n11208 );
not ( n11210 , n11206 );
not ( n11211 , n11207 );
and ( n11212 , n11210 , n11211 );
nor ( n11213 , n11209 , n11212 );
not ( n11214 , n11213 );
buf ( n11215 , n5118 );
nand ( n11216 , n6760 , n11215 );
buf ( n11217 , n5119 );
not ( n11218 , n11217 );
and ( n11219 , n11216 , n11218 );
not ( n11220 , n11216 );
buf ( n11221 , n11217 );
and ( n11222 , n11220 , n11221 );
nor ( n11223 , n11219 , n11222 );
not ( n11224 , n11223 );
or ( n11225 , n11214 , n11224 );
or ( n11226 , n11213 , n11223 );
nand ( n11227 , n11225 , n11226 );
xnor ( n11228 , n11204 , n11227 );
buf ( n11229 , n11228 );
buf ( n11230 , n5120 );
buf ( n11231 , n11230 );
not ( n11232 , n11231 );
not ( n11233 , n10472 );
or ( n11234 , n11232 , n11233 );
not ( n11235 , n11230 );
buf ( n11236 , n10471 );
nand ( n11237 , n11235 , n11236 );
nand ( n11238 , n11234 , n11237 );
buf ( n11239 , n5121 );
buf ( n11240 , n11239 );
and ( n11241 , n11238 , n11240 );
not ( n11242 , n11238 );
not ( n11243 , n11239 );
and ( n11244 , n11242 , n11243 );
nor ( n11245 , n11241 , n11244 );
buf ( n11246 , n5122 );
nand ( n11247 , n6760 , n11246 );
buf ( n11248 , n5123 );
xor ( n11249 , n11247 , n11248 );
xor ( n11250 , n11245 , n11249 );
buf ( n11251 , n5124 );
nand ( n11252 , n7478 , n11251 );
buf ( n11253 , n5125 );
not ( n11254 , n11253 );
and ( n11255 , n11252 , n11254 );
not ( n11256 , n11252 );
buf ( n11257 , n11253 );
and ( n11258 , n11256 , n11257 );
nor ( n11259 , n11255 , n11258 );
xnor ( n11260 , n11250 , n11259 );
not ( n11261 , n11260 );
not ( n11262 , n11261 );
buf ( n11263 , n5126 );
buf ( n11264 , n11263 );
not ( n11265 , n11264 );
and ( n11266 , n11262 , n11265 );
xor ( n11267 , n11245 , n11249 );
xnor ( n11268 , n11267 , n11259 );
not ( n11269 , n11268 );
and ( n11270 , n11269 , n11264 );
nor ( n11271 , n11266 , n11270 );
not ( n11272 , n11271 );
xor ( n11273 , n11229 , n11272 );
not ( n11274 , n11273 );
nand ( n11275 , n11191 , n11274 );
not ( n11276 , n6874 );
buf ( n11277 , n5127 );
buf ( n11278 , n11277 );
not ( n11279 , n11278 );
and ( n11280 , n11276 , n11279 );
not ( n11281 , n6873 );
and ( n11282 , n11281 , n11278 );
nor ( n11283 , n11280 , n11282 );
buf ( n11284 , n7006 );
and ( n11285 , n11283 , n11284 );
not ( n11286 , n11283 );
buf ( n11287 , n7012 );
and ( n11288 , n11286 , n11287 );
nor ( n11289 , n11285 , n11288 );
not ( n11290 , n11289 );
and ( n11291 , n11275 , n11290 );
not ( n11292 , n11275 );
and ( n11293 , n11292 , n11289 );
nor ( n11294 , n11291 , n11293 );
not ( n11295 , n11294 );
not ( n11296 , n11295 );
buf ( n11297 , n5128 );
buf ( n11298 , n11297 );
not ( n11299 , n11298 );
buf ( n11300 , n5129 );
not ( n11301 , n11300 );
not ( n11302 , n7805 );
buf ( n11303 , n5130 );
not ( n11304 , n11303 );
not ( n11305 , n11304 );
or ( n11306 , n11302 , n11305 );
not ( n11307 , n7804 );
buf ( n11308 , n11303 );
nand ( n11309 , n11307 , n11308 );
nand ( n11310 , n11306 , n11309 );
xor ( n11311 , n11301 , n11310 );
buf ( n11312 , n5131 );
buf ( n11313 , n5132 );
xor ( n11314 , n11312 , n11313 );
buf ( n11315 , n5133 );
nand ( n11316 , n6851 , n11315 );
xnor ( n11317 , n11314 , n11316 );
xor ( n11318 , n11311 , n11317 );
not ( n11319 , n11318 );
or ( n11320 , n11299 , n11319 );
or ( n11321 , n11318 , n11298 );
nand ( n11322 , n11320 , n11321 );
not ( n11323 , n11322 );
buf ( n11324 , n5134 );
buf ( n11325 , n11324 );
not ( n11326 , n11325 );
buf ( n11327 , n5135 );
not ( n11328 , n11327 );
not ( n11329 , n11328 );
or ( n11330 , n11326 , n11329 );
not ( n11331 , n11324 );
buf ( n11332 , n11327 );
nand ( n11333 , n11331 , n11332 );
nand ( n11334 , n11330 , n11333 );
buf ( n11335 , n5136 );
buf ( n11336 , n11335 );
and ( n11337 , n11334 , n11336 );
not ( n11338 , n11334 );
not ( n11339 , n11335 );
and ( n11340 , n11338 , n11339 );
nor ( n11341 , n11337 , n11340 );
buf ( n11342 , n5137 );
nand ( n11343 , n6905 , n11342 );
buf ( n11344 , n5138 );
buf ( n11345 , n11344 );
and ( n11346 , n11343 , n11345 );
not ( n11347 , n11343 );
not ( n11348 , n11344 );
and ( n11349 , n11347 , n11348 );
nor ( n11350 , n11346 , n11349 );
xor ( n11351 , n11341 , n11350 );
buf ( n11352 , n5139 );
nand ( n11353 , n7471 , n11352 );
buf ( n11354 , n5140 );
buf ( n11355 , n11354 );
and ( n11356 , n11353 , n11355 );
not ( n11357 , n11353 );
not ( n11358 , n11354 );
and ( n11359 , n11357 , n11358 );
nor ( n11360 , n11356 , n11359 );
xnor ( n11361 , n11351 , n11360 );
not ( n11362 , n11361 );
not ( n11363 , n11362 );
not ( n11364 , n11363 );
and ( n11365 , n11323 , n11364 );
and ( n11366 , n11322 , n11363 );
nor ( n11367 , n11365 , n11366 );
not ( n11368 , n11367 );
not ( n11369 , n11368 );
buf ( n11370 , n5141 );
buf ( n11371 , n11370 );
not ( n11372 , n11371 );
not ( n11373 , n8440 );
or ( n11374 , n11372 , n11373 );
not ( n11375 , n11371 );
nand ( n11376 , n11375 , n8433 );
nand ( n11377 , n11374 , n11376 );
not ( n11378 , n9687 );
buf ( n11379 , n11378 );
and ( n11380 , n11377 , n11379 );
not ( n11381 , n11377 );
and ( n11382 , n11381 , n9689 );
nor ( n11383 , n11380 , n11382 );
buf ( n11384 , n5142 );
buf ( n11385 , n11384 );
not ( n11386 , n11385 );
buf ( n11387 , n5143 );
buf ( n11388 , n11387 );
not ( n11389 , n11388 );
buf ( n11390 , n5144 );
not ( n11391 , n11390 );
not ( n11392 , n11391 );
or ( n11393 , n11389 , n11392 );
not ( n11394 , n11387 );
buf ( n11395 , n11390 );
nand ( n11396 , n11394 , n11395 );
nand ( n11397 , n11393 , n11396 );
buf ( n11398 , n5145 );
buf ( n11399 , n11398 );
and ( n11400 , n11397 , n11399 );
not ( n11401 , n11397 );
not ( n11402 , n11398 );
and ( n11403 , n11401 , n11402 );
nor ( n11404 , n11400 , n11403 );
buf ( n11405 , n5146 );
nand ( n11406 , n7094 , n11405 );
buf ( n11407 , n5147 );
buf ( n11408 , n11407 );
and ( n11409 , n11406 , n11408 );
not ( n11410 , n11406 );
not ( n11411 , n11407 );
and ( n11412 , n11410 , n11411 );
nor ( n11413 , n11409 , n11412 );
xor ( n11414 , n11404 , n11413 );
buf ( n11415 , n5148 );
nand ( n11416 , n8740 , n11415 );
buf ( n11417 , n5149 );
buf ( n11418 , n11417 );
and ( n11419 , n11416 , n11418 );
not ( n11420 , n11416 );
not ( n11421 , n11417 );
and ( n11422 , n11420 , n11421 );
nor ( n11423 , n11419 , n11422 );
buf ( n11424 , n11423 );
xnor ( n11425 , n11414 , n11424 );
not ( n11426 , n11425 );
or ( n11427 , n11386 , n11426 );
or ( n11428 , n11425 , n11385 );
nand ( n11429 , n11427 , n11428 );
buf ( n11430 , n5150 );
buf ( n11431 , n11430 );
not ( n11432 , n11431 );
buf ( n11433 , n5151 );
not ( n11434 , n11433 );
not ( n11435 , n11434 );
or ( n11436 , n11432 , n11435 );
not ( n11437 , n11430 );
buf ( n11438 , n11433 );
nand ( n11439 , n11437 , n11438 );
nand ( n11440 , n11436 , n11439 );
buf ( n11441 , n5152 );
buf ( n11442 , n11441 );
and ( n11443 , n11440 , n11442 );
not ( n11444 , n11440 );
not ( n11445 , n11441 );
and ( n11446 , n11444 , n11445 );
nor ( n11447 , n11443 , n11446 );
buf ( n11448 , n5153 );
nand ( n11449 , n7401 , n11448 );
buf ( n11450 , n5154 );
buf ( n11451 , n11450 );
and ( n11452 , n11449 , n11451 );
not ( n11453 , n11449 );
not ( n11454 , n11450 );
and ( n11455 , n11453 , n11454 );
nor ( n11456 , n11452 , n11455 );
xor ( n11457 , n11447 , n11456 );
buf ( n11458 , n5155 );
nand ( n11459 , n6622 , n11458 );
buf ( n11460 , n5156 );
buf ( n11461 , n11460 );
and ( n11462 , n11459 , n11461 );
not ( n11463 , n11459 );
not ( n11464 , n11460 );
and ( n11465 , n11463 , n11464 );
nor ( n11466 , n11462 , n11465 );
not ( n11467 , n11466 );
xor ( n11468 , n11457 , n11467 );
not ( n11469 , n11468 );
not ( n11470 , n11469 );
and ( n11471 , n11429 , n11470 );
not ( n11472 , n11429 );
buf ( n11473 , n11468 );
not ( n11474 , n11473 );
and ( n11475 , n11472 , n11474 );
nor ( n11476 , n11471 , n11475 );
nand ( n11477 , n11383 , n11476 );
not ( n11478 , n11477 );
or ( n11479 , n11369 , n11478 );
or ( n11480 , n11477 , n11368 );
nand ( n11481 , n11479 , n11480 );
buf ( n11482 , n5157 );
buf ( n11483 , n5158 );
buf ( n11484 , n11483 );
not ( n11485 , n11484 );
buf ( n11486 , n5159 );
not ( n11487 , n11486 );
not ( n11488 , n11487 );
or ( n11489 , n11485 , n11488 );
not ( n11490 , n11483 );
buf ( n11491 , n11486 );
nand ( n11492 , n11490 , n11491 );
nand ( n11493 , n11489 , n11492 );
xor ( n11494 , n11482 , n11493 );
buf ( n11495 , n5160 );
buf ( n11496 , n5161 );
not ( n11497 , n11496 );
xor ( n11498 , n11495 , n11497 );
buf ( n11499 , n5162 );
nand ( n11500 , n7617 , n11499 );
xnor ( n11501 , n11498 , n11500 );
xnor ( n11502 , n11494 , n11501 );
not ( n11503 , n11502 );
not ( n11504 , n11503 );
buf ( n11505 , n5163 );
buf ( n11506 , n11505 );
not ( n11507 , n11506 );
buf ( n11508 , n5164 );
not ( n11509 , n11508 );
not ( n11510 , n11509 );
or ( n11511 , n11507 , n11510 );
not ( n11512 , n11505 );
buf ( n11513 , n11508 );
nand ( n11514 , n11512 , n11513 );
nand ( n11515 , n11511 , n11514 );
buf ( n11516 , n5165 );
buf ( n11517 , n11516 );
and ( n11518 , n11515 , n11517 );
not ( n11519 , n11515 );
not ( n11520 , n11516 );
and ( n11521 , n11519 , n11520 );
nor ( n11522 , n11518 , n11521 );
buf ( n11523 , n5166 );
nand ( n11524 , n7133 , n11523 );
buf ( n11525 , n5167 );
not ( n11526 , n11525 );
and ( n11527 , n11524 , n11526 );
not ( n11528 , n11524 );
buf ( n11529 , n11525 );
and ( n11530 , n11528 , n11529 );
nor ( n11531 , n11527 , n11530 );
xor ( n11532 , n11522 , n11531 );
buf ( n11533 , n5168 );
nand ( n11534 , n8135 , n11533 );
buf ( n11535 , n5169 );
not ( n11536 , n11535 );
and ( n11537 , n11534 , n11536 );
not ( n11538 , n11534 );
buf ( n11539 , n11535 );
and ( n11540 , n11538 , n11539 );
nor ( n11541 , n11537 , n11540 );
xnor ( n11542 , n11532 , n11541 );
not ( n11543 , n11542 );
buf ( n11544 , n5170 );
buf ( n11545 , n11544 );
not ( n11546 , n11545 );
and ( n11547 , n11543 , n11546 );
and ( n11548 , n11542 , n11545 );
nor ( n11549 , n11547 , n11548 );
and ( n11550 , n11504 , n11549 );
not ( n11551 , n11504 );
not ( n11552 , n11549 );
and ( n11553 , n11551 , n11552 );
nor ( n11554 , n11550 , n11553 );
buf ( n11555 , n5171 );
buf ( n11556 , n11555 );
not ( n11557 , n11556 );
buf ( n11558 , n5172 );
not ( n11559 , n11558 );
not ( n11560 , n11559 );
or ( n11561 , n11557 , n11560 );
not ( n11562 , n11555 );
buf ( n11563 , n11558 );
nand ( n11564 , n11562 , n11563 );
nand ( n11565 , n11561 , n11564 );
buf ( n11566 , n5173 );
buf ( n11567 , n11566 );
and ( n11568 , n11565 , n11567 );
not ( n11569 , n11565 );
not ( n11570 , n11566 );
and ( n11571 , n11569 , n11570 );
nor ( n11572 , n11568 , n11571 );
buf ( n11573 , n5174 );
nand ( n11574 , n8923 , n11573 );
buf ( n11575 , n5175 );
buf ( n11576 , n11575 );
and ( n11577 , n11574 , n11576 );
not ( n11578 , n11574 );
not ( n11579 , n11575 );
and ( n11580 , n11578 , n11579 );
nor ( n11581 , n11577 , n11580 );
xor ( n11582 , n11572 , n11581 );
buf ( n11583 , n5176 );
nand ( n11584 , n8269 , n11583 );
buf ( n11585 , n5177 );
not ( n11586 , n11585 );
and ( n11587 , n11584 , n11586 );
not ( n11588 , n11584 );
buf ( n11589 , n11585 );
and ( n11590 , n11588 , n11589 );
nor ( n11591 , n11587 , n11590 );
xnor ( n11592 , n11582 , n11591 );
not ( n11593 , n11592 );
not ( n11594 , n11593 );
not ( n11595 , n9223 );
not ( n11596 , n11595 );
buf ( n11597 , n5178 );
buf ( n11598 , n11597 );
not ( n11599 , n11598 );
buf ( n11600 , n5179 );
not ( n11601 , n11600 );
not ( n11602 , n11601 );
or ( n11603 , n11599 , n11602 );
not ( n11604 , n11597 );
buf ( n11605 , n11600 );
nand ( n11606 , n11604 , n11605 );
nand ( n11607 , n11603 , n11606 );
buf ( n11608 , n5180 );
buf ( n11609 , n11608 );
and ( n11610 , n11607 , n11609 );
not ( n11611 , n11607 );
not ( n11612 , n11608 );
and ( n11613 , n11611 , n11612 );
nor ( n11614 , n11610 , n11613 );
buf ( n11615 , n5181 );
nand ( n11616 , n6660 , n11615 );
buf ( n11617 , n5182 );
xor ( n11618 , n11616 , n11617 );
xor ( n11619 , n11614 , n11618 );
buf ( n11620 , n5183 );
nand ( n11621 , n7134 , n11620 );
buf ( n11622 , n5184 );
buf ( n11623 , n11622 );
and ( n11624 , n11621 , n11623 );
not ( n11625 , n11621 );
not ( n11626 , n11622 );
and ( n11627 , n11625 , n11626 );
nor ( n11628 , n11624 , n11627 );
xor ( n11629 , n11619 , n11628 );
not ( n11630 , n11629 );
or ( n11631 , n11596 , n11630 );
or ( n11632 , n11629 , n11595 );
nand ( n11633 , n11631 , n11632 );
not ( n11634 , n11633 );
or ( n11635 , n11594 , n11634 );
or ( n11636 , n11633 , n11593 );
nand ( n11637 , n11635 , n11636 );
nand ( n11638 , n11554 , n11637 );
not ( n11639 , n11638 );
buf ( n11640 , n5185 );
buf ( n11641 , n11640 );
not ( n11642 , n11641 );
buf ( n11643 , n5186 );
buf ( n11644 , n11643 );
not ( n11645 , n11644 );
buf ( n11646 , n5187 );
not ( n11647 , n11646 );
not ( n11648 , n11647 );
or ( n11649 , n11645 , n11648 );
not ( n11650 , n11643 );
buf ( n11651 , n11646 );
nand ( n11652 , n11650 , n11651 );
nand ( n11653 , n11649 , n11652 );
buf ( n11654 , n5188 );
not ( n11655 , n11654 );
and ( n11656 , n11653 , n11655 );
not ( n11657 , n11653 );
buf ( n11658 , n11654 );
and ( n11659 , n11657 , n11658 );
nor ( n11660 , n11656 , n11659 );
buf ( n11661 , n5189 );
nand ( n11662 , n7183 , n11661 );
buf ( n11663 , n5190 );
buf ( n11664 , n11663 );
and ( n11665 , n11662 , n11664 );
not ( n11666 , n11662 );
not ( n11667 , n11663 );
and ( n11668 , n11666 , n11667 );
nor ( n11669 , n11665 , n11668 );
xor ( n11670 , n11660 , n11669 );
xnor ( n11671 , n11670 , n10291 );
not ( n11672 , n11671 );
not ( n11673 , n11672 );
not ( n11674 , n11673 );
or ( n11675 , n11642 , n11674 );
not ( n11676 , n11641 );
nand ( n11677 , n11676 , n11672 );
nand ( n11678 , n11675 , n11677 );
buf ( n11679 , n5191 );
buf ( n11680 , n11679 );
not ( n11681 , n11680 );
buf ( n11682 , n5192 );
not ( n11683 , n11682 );
not ( n11684 , n11683 );
or ( n11685 , n11681 , n11684 );
not ( n11686 , n11679 );
buf ( n11687 , n11682 );
nand ( n11688 , n11686 , n11687 );
nand ( n11689 , n11685 , n11688 );
buf ( n11690 , n5193 );
buf ( n11691 , n11690 );
and ( n11692 , n11689 , n11691 );
not ( n11693 , n11689 );
not ( n11694 , n11690 );
and ( n11695 , n11693 , n11694 );
nor ( n11696 , n11692 , n11695 );
buf ( n11697 , n5194 );
nand ( n11698 , n7195 , n11697 );
buf ( n11699 , n5195 );
buf ( n11700 , n11699 );
and ( n11701 , n11698 , n11700 );
not ( n11702 , n11698 );
not ( n11703 , n11699 );
and ( n11704 , n11702 , n11703 );
nor ( n11705 , n11701 , n11704 );
xor ( n11706 , n11696 , n11705 );
buf ( n11707 , n5196 );
nand ( n11708 , n10577 , n11707 );
buf ( n11709 , n5197 );
buf ( n11710 , n11709 );
and ( n11711 , n11708 , n11710 );
not ( n11712 , n11708 );
not ( n11713 , n11709 );
and ( n11714 , n11712 , n11713 );
nor ( n11715 , n11711 , n11714 );
xnor ( n11716 , n11706 , n11715 );
buf ( n11717 , n11716 );
and ( n11718 , n11678 , n11717 );
not ( n11719 , n11678 );
not ( n11720 , n11717 );
and ( n11721 , n11719 , n11720 );
nor ( n11722 , n11718 , n11721 );
not ( n11723 , n11722 );
not ( n11724 , n11723 );
and ( n11725 , n11639 , n11724 );
and ( n11726 , n11638 , n11723 );
nor ( n11727 , n11725 , n11726 );
nor ( n11728 , n11481 , n11727 );
not ( n11729 , n11728 );
nand ( n11730 , n11481 , n11727 );
nand ( n11731 , n11729 , n11730 );
not ( n11732 , n11731 );
and ( n11733 , n11296 , n11732 );
and ( n11734 , n11295 , n11731 );
nor ( n11735 , n11733 , n11734 );
not ( n11736 , n11735 );
and ( n11737 , n11144 , n11736 );
and ( n11738 , n11143 , n11735 );
nor ( n11739 , n11737 , n11738 );
not ( n11740 , n11739 );
not ( n11741 , n11740 );
and ( n11742 , n10767 , n11741 );
not ( n11743 , n10767 );
not ( n11744 , n11735 );
not ( n11745 , n11744 );
not ( n11746 , n11143 );
not ( n11747 , n11746 );
or ( n11748 , n11745 , n11747 );
nand ( n11749 , n11735 , n11143 );
nand ( n11750 , n11748 , n11749 );
buf ( n11751 , n11750 );
and ( n11752 , n11743 , n11751 );
nor ( n11753 , n11742 , n11752 );
nand ( n11754 , n9430 , n11753 );
buf ( n11755 , n6758 );
buf ( n11756 , n9123 );
xor ( n11757 , n11755 , n11756 );
buf ( n11758 , n5198 );
buf ( n11759 , n11758 );
not ( n11760 , n11759 );
buf ( n11761 , n5199 );
not ( n11762 , n11761 );
not ( n11763 , n11762 );
or ( n11764 , n11760 , n11763 );
not ( n11765 , n11758 );
buf ( n11766 , n11761 );
nand ( n11767 , n11765 , n11766 );
nand ( n11768 , n11764 , n11767 );
not ( n11769 , n11768 );
xor ( n11770 , n8444 , n11769 );
buf ( n11771 , n5200 );
buf ( n11772 , n5201 );
xor ( n11773 , n11771 , n11772 );
buf ( n11774 , n5202 );
nand ( n11775 , n6906 , n11774 );
xnor ( n11776 , n11773 , n11775 );
xnor ( n11777 , n11770 , n11776 );
buf ( n11778 , n11777 );
xnor ( n11779 , n11757 , n11778 );
not ( n11780 , n11779 );
buf ( n11781 , n5203 );
buf ( n11782 , n11781 );
not ( n11783 , n11782 );
buf ( n11784 , n5204 );
buf ( n11785 , n11784 );
not ( n11786 , n11785 );
buf ( n11787 , n5205 );
not ( n11788 , n11787 );
not ( n11789 , n11788 );
or ( n11790 , n11786 , n11789 );
not ( n11791 , n11784 );
buf ( n11792 , n11787 );
nand ( n11793 , n11791 , n11792 );
nand ( n11794 , n11790 , n11793 );
buf ( n11795 , n5206 );
buf ( n11796 , n11795 );
and ( n11797 , n11794 , n11796 );
not ( n11798 , n11794 );
not ( n11799 , n11795 );
and ( n11800 , n11798 , n11799 );
nor ( n11801 , n11797 , n11800 );
buf ( n11802 , n5207 );
nand ( n11803 , n6804 , n11802 );
buf ( n11804 , n5208 );
not ( n11805 , n11804 );
and ( n11806 , n11803 , n11805 );
not ( n11807 , n11803 );
buf ( n11808 , n11804 );
and ( n11809 , n11807 , n11808 );
nor ( n11810 , n11806 , n11809 );
xor ( n11811 , n11801 , n11810 );
buf ( n11812 , n5209 );
nand ( n11813 , n9159 , n11812 );
buf ( n11814 , n5210 );
not ( n11815 , n11814 );
and ( n11816 , n11813 , n11815 );
not ( n11817 , n11813 );
buf ( n11818 , n11814 );
and ( n11819 , n11817 , n11818 );
nor ( n11820 , n11816 , n11819 );
xnor ( n11821 , n11811 , n11820 );
not ( n11822 , n11821 );
not ( n11823 , n11822 );
not ( n11824 , n11823 );
or ( n11825 , n11783 , n11824 );
not ( n11826 , n11781 );
nand ( n11827 , n11822 , n11826 );
nand ( n11828 , n11825 , n11827 );
not ( n11829 , n11828 );
buf ( n11830 , n5211 );
buf ( n11831 , n11830 );
not ( n11832 , n11831 );
buf ( n11833 , n5212 );
not ( n11834 , n11833 );
not ( n11835 , n11834 );
or ( n11836 , n11832 , n11835 );
not ( n11837 , n11830 );
buf ( n11838 , n11833 );
nand ( n11839 , n11837 , n11838 );
nand ( n11840 , n11836 , n11839 );
buf ( n11841 , n5213 );
buf ( n11842 , n11841 );
and ( n11843 , n11840 , n11842 );
not ( n11844 , n11840 );
not ( n11845 , n11841 );
and ( n11846 , n11844 , n11845 );
nor ( n11847 , n11843 , n11846 );
buf ( n11848 , n5214 );
nand ( n11849 , n7133 , n11848 );
buf ( n11850 , n5215 );
buf ( n11851 , n11850 );
and ( n11852 , n11849 , n11851 );
not ( n11853 , n11849 );
not ( n11854 , n11850 );
and ( n11855 , n11853 , n11854 );
nor ( n11856 , n11852 , n11855 );
xor ( n11857 , n11847 , n11856 );
buf ( n11858 , n5216 );
nand ( n11859 , n7617 , n11858 );
buf ( n11860 , n5217 );
not ( n11861 , n11860 );
and ( n11862 , n11859 , n11861 );
not ( n11863 , n11859 );
buf ( n11864 , n11860 );
and ( n11865 , n11863 , n11864 );
nor ( n11866 , n11862 , n11865 );
xor ( n11867 , n11857 , n11866 );
buf ( n11868 , n11867 );
not ( n11869 , n11868 );
and ( n11870 , n11829 , n11869 );
and ( n11871 , n11828 , n11868 );
nor ( n11872 , n11870 , n11871 );
not ( n11873 , n11872 );
nand ( n11874 , n11780 , n11873 );
buf ( n11875 , n5218 );
nand ( n11876 , n6985 , n11875 );
buf ( n11877 , n5219 );
not ( n11878 , n11877 );
and ( n11879 , n11876 , n11878 );
not ( n11880 , n11876 );
buf ( n11881 , n11877 );
and ( n11882 , n11880 , n11881 );
nor ( n11883 , n11879 , n11882 );
xor ( n11884 , n11883 , n11269 );
buf ( n11885 , n5220 );
buf ( n11886 , n11885 );
not ( n11887 , n11886 );
buf ( n11888 , n5221 );
not ( n11889 , n11888 );
not ( n11890 , n11889 );
or ( n11891 , n11887 , n11890 );
not ( n11892 , n11885 );
buf ( n11893 , n11888 );
nand ( n11894 , n11892 , n11893 );
nand ( n11895 , n11891 , n11894 );
not ( n11896 , n11895 );
buf ( n11897 , n5222 );
buf ( n11898 , n5223 );
nand ( n11899 , n7195 , n11898 );
buf ( n11900 , n5224 );
buf ( n11901 , n11900 );
and ( n11902 , n11899 , n11901 );
not ( n11903 , n11899 );
not ( n11904 , n11900 );
and ( n11905 , n11903 , n11904 );
nor ( n11906 , n11902 , n11905 );
xor ( n11907 , n11897 , n11906 );
buf ( n11908 , n5225 );
nand ( n11909 , n6608 , n11908 );
buf ( n11910 , n5226 );
not ( n11911 , n11910 );
and ( n11912 , n11909 , n11911 );
not ( n11913 , n11909 );
buf ( n11914 , n11910 );
and ( n11915 , n11913 , n11914 );
nor ( n11916 , n11912 , n11915 );
xnor ( n11917 , n11907 , n11916 );
not ( n11918 , n11917 );
not ( n11919 , n11918 );
or ( n11920 , n11896 , n11919 );
not ( n11921 , n11895 );
nand ( n11922 , n11917 , n11921 );
nand ( n11923 , n11920 , n11922 );
not ( n11924 , n11923 );
xnor ( n11925 , n11884 , n11924 );
and ( n11926 , n11874 , n11925 );
not ( n11927 , n11874 );
not ( n11928 , n11925 );
and ( n11929 , n11927 , n11928 );
nor ( n11930 , n11926 , n11929 );
not ( n11931 , n11930 );
not ( n11932 , n11931 );
buf ( n11933 , n5227 );
nand ( n11934 , n7413 , n11933 );
buf ( n11935 , n5228 );
not ( n11936 , n11935 );
and ( n11937 , n11934 , n11936 );
not ( n11938 , n11934 );
buf ( n11939 , n11935 );
and ( n11940 , n11938 , n11939 );
nor ( n11941 , n11937 , n11940 );
not ( n11942 , n11941 );
not ( n11943 , n9937 );
not ( n11944 , n9947 );
or ( n11945 , n11943 , n11944 );
or ( n11946 , n9937 , n9947 );
nand ( n11947 , n11945 , n11946 );
xnor ( n11948 , n11947 , n9928 );
not ( n11949 , n11948 );
or ( n11950 , n11942 , n11949 );
not ( n11951 , n11941 );
nand ( n11952 , n11951 , n9948 );
nand ( n11953 , n11950 , n11952 );
not ( n11954 , n11953 );
buf ( n11955 , n5229 );
buf ( n11956 , n11955 );
not ( n11957 , n11956 );
buf ( n11958 , n5230 );
not ( n11959 , n11958 );
not ( n11960 , n11959 );
or ( n11961 , n11957 , n11960 );
not ( n11962 , n11955 );
buf ( n11963 , n11958 );
nand ( n11964 , n11962 , n11963 );
nand ( n11965 , n11961 , n11964 );
buf ( n11966 , n5231 );
not ( n11967 , n11966 );
and ( n11968 , n11965 , n11967 );
not ( n11969 , n11965 );
buf ( n11970 , n11966 );
and ( n11971 , n11969 , n11970 );
nor ( n11972 , n11968 , n11971 );
buf ( n11973 , n5232 );
nand ( n11974 , n7230 , n11973 );
buf ( n11975 , n5233 );
buf ( n11976 , n11975 );
and ( n11977 , n11974 , n11976 );
not ( n11978 , n11974 );
not ( n11979 , n11975 );
and ( n11980 , n11978 , n11979 );
nor ( n11981 , n11977 , n11980 );
xor ( n11982 , n11972 , n11981 );
buf ( n11983 , n5234 );
nand ( n11984 , n10577 , n11983 );
buf ( n11985 , n5235 );
buf ( n11986 , n11985 );
and ( n11987 , n11984 , n11986 );
not ( n11988 , n11984 );
not ( n11989 , n11985 );
and ( n11990 , n11988 , n11989 );
nor ( n11991 , n11987 , n11990 );
xnor ( n11992 , n11982 , n11991 );
not ( n11993 , n11992 );
not ( n11994 , n11993 );
and ( n11995 , n11954 , n11994 );
buf ( n11996 , n11992 );
not ( n11997 , n11996 );
and ( n11998 , n11953 , n11997 );
nor ( n11999 , n11995 , n11998 );
buf ( n12000 , n5236 );
not ( n12001 , n12000 );
buf ( n12002 , n5237 );
not ( n12003 , n12002 );
buf ( n12004 , n5238 );
buf ( n12005 , n12004 );
and ( n12006 , n12003 , n12005 );
not ( n12007 , n12003 );
not ( n12008 , n12004 );
and ( n12009 , n12007 , n12008 );
nor ( n12010 , n12006 , n12009 );
xor ( n12011 , n12001 , n12010 );
buf ( n12012 , n5239 );
buf ( n12013 , n5240 );
xor ( n12014 , n12012 , n12013 );
buf ( n12015 , n5241 );
nand ( n12016 , n9159 , n12015 );
xnor ( n12017 , n12014 , n12016 );
xnor ( n12018 , n12011 , n12017 );
buf ( n12019 , n12018 );
not ( n12020 , n12019 );
buf ( n12021 , n5242 );
nand ( n12022 , n6660 , n12021 );
buf ( n12023 , n5243 );
buf ( n12024 , n12023 );
and ( n12025 , n12022 , n12024 );
not ( n12026 , n12022 );
not ( n12027 , n12023 );
and ( n12028 , n12026 , n12027 );
nor ( n12029 , n12025 , n12028 );
buf ( n12030 , n12029 );
buf ( n12031 , n5244 );
nand ( n12032 , n6607 , n12031 );
buf ( n12033 , n5245 );
buf ( n12034 , n12033 );
and ( n12035 , n12032 , n12034 );
not ( n12036 , n12032 );
not ( n12037 , n12033 );
and ( n12038 , n12036 , n12037 );
nor ( n12039 , n12035 , n12038 );
not ( n12040 , n12039 );
buf ( n12041 , n5246 );
nand ( n12042 , n7471 , n12041 );
buf ( n12043 , n5247 );
not ( n12044 , n12043 );
and ( n12045 , n12042 , n12044 );
not ( n12046 , n12042 );
buf ( n12047 , n12043 );
and ( n12048 , n12046 , n12047 );
nor ( n12049 , n12045 , n12048 );
not ( n12050 , n12049 );
or ( n12051 , n12040 , n12050 );
or ( n12052 , n12039 , n12049 );
nand ( n12053 , n12051 , n12052 );
buf ( n12054 , n5248 );
buf ( n12055 , n12054 );
not ( n12056 , n12055 );
buf ( n12057 , n5249 );
not ( n12058 , n12057 );
not ( n12059 , n12058 );
or ( n12060 , n12056 , n12059 );
not ( n12061 , n12054 );
buf ( n12062 , n12057 );
nand ( n12063 , n12061 , n12062 );
nand ( n12064 , n12060 , n12063 );
buf ( n12065 , n5250 );
not ( n12066 , n12065 );
and ( n12067 , n12064 , n12066 );
not ( n12068 , n12064 );
buf ( n12069 , n12065 );
and ( n12070 , n12068 , n12069 );
nor ( n12071 , n12067 , n12070 );
not ( n12072 , n12071 );
and ( n12073 , n12053 , n12072 );
not ( n12074 , n12053 );
and ( n12075 , n12074 , n12071 );
nor ( n12076 , n12073 , n12075 );
and ( n12077 , n12030 , n12076 );
not ( n12078 , n12030 );
xor ( n12079 , n12071 , n12039 );
xnor ( n12080 , n12079 , n12049 );
and ( n12081 , n12078 , n12080 );
nor ( n12082 , n12077 , n12081 );
not ( n12083 , n12082 );
not ( n12084 , n12083 );
or ( n12085 , n12020 , n12084 );
buf ( n12086 , n12000 );
xor ( n12087 , n12086 , n12010 );
xnor ( n12088 , n12087 , n12017 );
buf ( n12089 , n12088 );
nand ( n12090 , n12082 , n12089 );
nand ( n12091 , n12085 , n12090 );
nand ( n12092 , n11999 , n12091 );
not ( n12093 , n12092 );
buf ( n12094 , n5251 );
buf ( n12095 , n12094 );
not ( n12096 , n12095 );
not ( n12097 , n7006 );
or ( n12098 , n12096 , n12097 );
or ( n12099 , n7006 , n12095 );
nand ( n12100 , n12098 , n12099 );
and ( n12101 , n12100 , n7055 );
not ( n12102 , n12100 );
and ( n12103 , n12102 , n7054 );
nor ( n12104 , n12101 , n12103 );
not ( n12105 , n12104 );
not ( n12106 , n12105 );
and ( n12107 , n12093 , n12106 );
and ( n12108 , n12092 , n12105 );
nor ( n12109 , n12107 , n12108 );
not ( n12110 , n12109 );
buf ( n12111 , n5252 );
nand ( n12112 , n6863 , n12111 );
buf ( n12113 , n5253 );
buf ( n12114 , n12113 );
and ( n12115 , n12112 , n12114 );
not ( n12116 , n12112 );
not ( n12117 , n12113 );
and ( n12118 , n12116 , n12117 );
nor ( n12119 , n12115 , n12118 );
buf ( n12120 , n12119 );
not ( n12121 , n12120 );
buf ( n12122 , n5254 );
buf ( n12123 , n12122 );
not ( n12124 , n12123 );
buf ( n12125 , n5255 );
not ( n12126 , n12125 );
not ( n12127 , n12126 );
or ( n12128 , n12124 , n12127 );
not ( n12129 , n12122 );
buf ( n12130 , n12125 );
nand ( n12131 , n12129 , n12130 );
nand ( n12132 , n12128 , n12131 );
and ( n12133 , n12132 , n11020 );
not ( n12134 , n12132 );
not ( n12135 , n11019 );
and ( n12136 , n12134 , n12135 );
nor ( n12137 , n12133 , n12136 );
buf ( n12138 , n5256 );
nand ( n12139 , n7288 , n12138 );
buf ( n12140 , n5257 );
buf ( n12141 , n12140 );
and ( n12142 , n12139 , n12141 );
not ( n12143 , n12139 );
not ( n12144 , n12140 );
and ( n12145 , n12143 , n12144 );
nor ( n12146 , n12142 , n12145 );
xor ( n12147 , n12137 , n12146 );
buf ( n12148 , n5258 );
nand ( n12149 , n7471 , n12148 );
buf ( n12150 , n5259 );
buf ( n12151 , n12150 );
and ( n12152 , n12149 , n12151 );
not ( n12153 , n12149 );
not ( n12154 , n12150 );
and ( n12155 , n12153 , n12154 );
nor ( n12156 , n12152 , n12155 );
xor ( n12157 , n12147 , n12156 );
not ( n12158 , n12157 );
or ( n12159 , n12121 , n12158 );
or ( n12160 , n12157 , n12120 );
nand ( n12161 , n12159 , n12160 );
buf ( n12162 , n5260 );
buf ( n12163 , n12162 );
not ( n12164 , n12163 );
buf ( n12165 , n5261 );
not ( n12166 , n12165 );
not ( n12167 , n12166 );
or ( n12168 , n12164 , n12167 );
not ( n12169 , n12162 );
buf ( n12170 , n12165 );
nand ( n12171 , n12169 , n12170 );
nand ( n12172 , n12168 , n12171 );
buf ( n12173 , n5262 );
buf ( n12174 , n12173 );
and ( n12175 , n12172 , n12174 );
not ( n12176 , n12172 );
not ( n12177 , n12173 );
and ( n12178 , n12176 , n12177 );
nor ( n12179 , n12175 , n12178 );
buf ( n12180 , n5263 );
nand ( n12181 , n10204 , n12180 );
buf ( n12182 , n5264 );
buf ( n12183 , n12182 );
and ( n12184 , n12181 , n12183 );
not ( n12185 , n12181 );
not ( n12186 , n12182 );
and ( n12187 , n12185 , n12186 );
nor ( n12188 , n12184 , n12187 );
xor ( n12189 , n12179 , n12188 );
buf ( n12190 , n5265 );
nand ( n12191 , n7750 , n12190 );
buf ( n12192 , n5266 );
buf ( n12193 , n12192 );
and ( n12194 , n12191 , n12193 );
not ( n12195 , n12191 );
not ( n12196 , n12192 );
and ( n12197 , n12195 , n12196 );
nor ( n12198 , n12194 , n12197 );
xnor ( n12199 , n12189 , n12198 );
buf ( n12200 , n12199 );
buf ( n12201 , n12200 );
and ( n12202 , n12161 , n12201 );
not ( n12203 , n12161 );
not ( n12204 , n12199 );
buf ( n12205 , n12204 );
and ( n12206 , n12203 , n12205 );
nor ( n12207 , n12202 , n12206 );
not ( n12208 , n12207 );
buf ( n12209 , n5267 );
nand ( n12210 , n7126 , n12209 );
buf ( n12211 , n5268 );
not ( n12212 , n12211 );
and ( n12213 , n12210 , n12212 );
not ( n12214 , n12210 );
buf ( n12215 , n12211 );
and ( n12216 , n12214 , n12215 );
nor ( n12217 , n12213 , n12216 );
buf ( n12218 , n12217 );
not ( n12219 , n12218 );
buf ( n12220 , n5269 );
buf ( n12221 , n12220 );
buf ( n12222 , n5270 );
not ( n12223 , n12222 );
nand ( n12224 , n12223 , n9492 );
not ( n12225 , n9491 );
buf ( n12226 , n12222 );
nand ( n12227 , n12225 , n12226 );
and ( n12228 , n12224 , n12227 );
xor ( n12229 , n12221 , n12228 );
buf ( n12230 , n5271 );
buf ( n12231 , n5272 );
xor ( n12232 , n12230 , n12231 );
buf ( n12233 , n5273 );
nand ( n12234 , n6985 , n12233 );
xnor ( n12235 , n12232 , n12234 );
xor ( n12236 , n12229 , n12235 );
not ( n12237 , n12236 );
or ( n12238 , n12219 , n12237 );
or ( n12239 , n12236 , n12218 );
nand ( n12240 , n12238 , n12239 );
buf ( n12241 , n5274 );
buf ( n12242 , n12241 );
not ( n12243 , n12242 );
buf ( n12244 , n5275 );
not ( n12245 , n12244 );
not ( n12246 , n12245 );
or ( n12247 , n12243 , n12246 );
not ( n12248 , n12241 );
buf ( n12249 , n12244 );
nand ( n12250 , n12248 , n12249 );
nand ( n12251 , n12247 , n12250 );
buf ( n12252 , n5276 );
not ( n12253 , n12252 );
and ( n12254 , n12251 , n12253 );
not ( n12255 , n12251 );
buf ( n12256 , n12252 );
and ( n12257 , n12255 , n12256 );
nor ( n12258 , n12254 , n12257 );
buf ( n12259 , n5277 );
nand ( n12260 , n8519 , n12259 );
buf ( n12261 , n5278 );
buf ( n12262 , n12261 );
and ( n12263 , n12260 , n12262 );
not ( n12264 , n12260 );
not ( n12265 , n12261 );
and ( n12266 , n12264 , n12265 );
nor ( n12267 , n12263 , n12266 );
xor ( n12268 , n12258 , n12267 );
not ( n12269 , n7161 );
xnor ( n12270 , n12268 , n12269 );
buf ( n12271 , n12270 );
and ( n12272 , n12240 , n12271 );
not ( n12273 , n12240 );
xor ( n12274 , n12258 , n7161 );
buf ( n12275 , n12267 );
xnor ( n12276 , n12274 , n12275 );
buf ( n12277 , n12276 );
and ( n12278 , n12273 , n12277 );
nor ( n12279 , n12272 , n12278 );
nand ( n12280 , n12208 , n12279 );
buf ( n12281 , n5279 );
not ( n12282 , n12281 );
buf ( n12283 , n5280 );
buf ( n12284 , n12283 );
not ( n12285 , n12284 );
buf ( n12286 , n5281 );
not ( n12287 , n12286 );
not ( n12288 , n12287 );
or ( n12289 , n12285 , n12288 );
not ( n12290 , n12283 );
buf ( n12291 , n12286 );
nand ( n12292 , n12290 , n12291 );
nand ( n12293 , n12289 , n12292 );
not ( n12294 , n8902 );
and ( n12295 , n12293 , n12294 );
not ( n12296 , n12293 );
and ( n12297 , n12296 , n8903 );
nor ( n12298 , n12295 , n12297 );
buf ( n12299 , n5282 );
nand ( n12300 , n7955 , n12299 );
buf ( n12301 , n5283 );
buf ( n12302 , n12301 );
and ( n12303 , n12300 , n12302 );
not ( n12304 , n12300 );
not ( n12305 , n12301 );
and ( n12306 , n12304 , n12305 );
nor ( n12307 , n12303 , n12306 );
xor ( n12308 , n12298 , n12307 );
buf ( n12309 , n5284 );
nand ( n12310 , n7288 , n12309 );
buf ( n12311 , n5285 );
buf ( n12312 , n12311 );
and ( n12313 , n12310 , n12312 );
not ( n12314 , n12310 );
not ( n12315 , n12311 );
and ( n12316 , n12314 , n12315 );
nor ( n12317 , n12313 , n12316 );
xor ( n12318 , n12308 , n12317 );
not ( n12319 , n12318 );
or ( n12320 , n12282 , n12319 );
not ( n12321 , n12281 );
xor ( n12322 , n12298 , n12317 );
buf ( n12323 , n12307 );
xnor ( n12324 , n12322 , n12323 );
nand ( n12325 , n12321 , n12324 );
nand ( n12326 , n12320 , n12325 );
buf ( n12327 , n5286 );
buf ( n12328 , n12327 );
not ( n12329 , n12328 );
buf ( n12330 , n5287 );
not ( n12331 , n12330 );
not ( n12332 , n12331 );
or ( n12333 , n12329 , n12332 );
not ( n12334 , n12327 );
buf ( n12335 , n12330 );
nand ( n12336 , n12334 , n12335 );
nand ( n12337 , n12333 , n12336 );
buf ( n12338 , n5288 );
buf ( n12339 , n12338 );
and ( n12340 , n12337 , n12339 );
not ( n12341 , n12337 );
not ( n12342 , n12338 );
and ( n12343 , n12341 , n12342 );
nor ( n12344 , n12340 , n12343 );
buf ( n12345 , n5289 );
nand ( n12346 , n7133 , n12345 );
buf ( n12347 , n5290 );
not ( n12348 , n12347 );
and ( n12349 , n12346 , n12348 );
not ( n12350 , n12346 );
buf ( n12351 , n12347 );
and ( n12352 , n12350 , n12351 );
nor ( n12353 , n12349 , n12352 );
xor ( n12354 , n12344 , n12353 );
buf ( n12355 , n5291 );
nand ( n12356 , n7196 , n12355 );
buf ( n12357 , n5292 );
not ( n12358 , n12357 );
and ( n12359 , n12356 , n12358 );
not ( n12360 , n12356 );
buf ( n12361 , n12357 );
and ( n12362 , n12360 , n12361 );
nor ( n12363 , n12359 , n12362 );
xnor ( n12364 , n12354 , n12363 );
not ( n12365 , n12364 );
not ( n12366 , n12365 );
and ( n12367 , n12326 , n12366 );
not ( n12368 , n12326 );
buf ( n12369 , n12364 );
not ( n12370 , n12369 );
and ( n12371 , n12368 , n12370 );
nor ( n12372 , n12367 , n12371 );
and ( n12373 , n12280 , n12372 );
not ( n12374 , n12280 );
not ( n12375 , n12372 );
and ( n12376 , n12374 , n12375 );
nor ( n12377 , n12373 , n12376 );
not ( n12378 , n12377 );
or ( n12379 , n12110 , n12378 );
or ( n12380 , n12377 , n12109 );
nand ( n12381 , n12379 , n12380 );
buf ( n12382 , n10373 );
not ( n12383 , n12382 );
buf ( n12384 , n5293 );
buf ( n12385 , n5294 );
nand ( n12386 , n7920 , n12385 );
not ( n12387 , n12386 );
buf ( n12388 , n5295 );
not ( n12389 , n12388 );
and ( n12390 , n12387 , n12389 );
nand ( n12391 , n6803 , n12385 );
and ( n12392 , n12391 , n12388 );
nor ( n12393 , n12390 , n12392 );
xor ( n12394 , n12384 , n12393 );
buf ( n12395 , n5296 );
not ( n12396 , n12395 );
buf ( n12397 , n5297 );
nand ( n12398 , n7750 , n12397 );
not ( n12399 , n12398 );
or ( n12400 , n12396 , n12399 );
buf ( n12401 , n7920 );
nand ( n12402 , n12401 , n12397 );
or ( n12403 , n12402 , n12395 );
nand ( n12404 , n12400 , n12403 );
xnor ( n12405 , n12394 , n12404 );
not ( n12406 , n12405 );
buf ( n12407 , n5298 );
buf ( n12408 , n12407 );
not ( n12409 , n12408 );
buf ( n12410 , n5299 );
not ( n12411 , n12410 );
not ( n12412 , n12411 );
or ( n12413 , n12409 , n12412 );
not ( n12414 , n12407 );
buf ( n12415 , n12410 );
nand ( n12416 , n12414 , n12415 );
nand ( n12417 , n12413 , n12416 );
not ( n12418 , n12417 );
not ( n12419 , n12418 );
and ( n12420 , n12406 , n12419 );
and ( n12421 , n12405 , n12418 );
nor ( n12422 , n12420 , n12421 );
not ( n12423 , n12422 );
or ( n12424 , n12383 , n12423 );
or ( n12425 , n12422 , n12382 );
nand ( n12426 , n12424 , n12425 );
buf ( n12427 , n5300 );
buf ( n12428 , n12427 );
not ( n12429 , n12428 );
buf ( n12430 , n5301 );
not ( n12431 , n12430 );
not ( n12432 , n12431 );
or ( n12433 , n12429 , n12432 );
not ( n12434 , n12427 );
buf ( n12435 , n12430 );
nand ( n12436 , n12434 , n12435 );
nand ( n12437 , n12433 , n12436 );
buf ( n12438 , n5302 );
not ( n12439 , n12438 );
and ( n12440 , n12437 , n12439 );
not ( n12441 , n12437 );
buf ( n12442 , n12438 );
and ( n12443 , n12441 , n12442 );
nor ( n12444 , n12440 , n12443 );
buf ( n12445 , n5303 );
nand ( n12446 , n7477 , n12445 );
buf ( n12447 , n5304 );
buf ( n12448 , n12447 );
and ( n12449 , n12446 , n12448 );
not ( n12450 , n12446 );
not ( n12451 , n12447 );
and ( n12452 , n12450 , n12451 );
nor ( n12453 , n12449 , n12452 );
xor ( n12454 , n12444 , n12453 );
buf ( n12455 , n5305 );
nand ( n12456 , n7356 , n12455 );
buf ( n12457 , n5306 );
not ( n12458 , n12457 );
and ( n12459 , n12456 , n12458 );
not ( n12460 , n12456 );
buf ( n12461 , n12457 );
and ( n12462 , n12460 , n12461 );
nor ( n12463 , n12459 , n12462 );
xnor ( n12464 , n12454 , n12463 );
buf ( n12465 , n12464 );
and ( n12466 , n12426 , n12465 );
not ( n12467 , n12426 );
not ( n12468 , n12465 );
and ( n12469 , n12467 , n12468 );
nor ( n12470 , n12466 , n12469 );
not ( n12471 , n12470 );
not ( n12472 , n12275 );
not ( n12473 , n12472 );
not ( n12474 , n9544 );
or ( n12475 , n12473 , n12474 );
nand ( n12476 , n9538 , n12275 );
nand ( n12477 , n12475 , n12476 );
buf ( n12478 , n7255 );
not ( n12479 , n12478 );
and ( n12480 , n12477 , n12479 );
not ( n12481 , n12477 );
and ( n12482 , n12481 , n12478 );
nor ( n12483 , n12480 , n12482 );
nand ( n12484 , n12471 , n12483 );
not ( n12485 , n12484 );
buf ( n12486 , n5307 );
not ( n12487 , n12486 );
buf ( n12488 , n5308 );
buf ( n12489 , n12488 );
not ( n12490 , n12489 );
buf ( n12491 , n5309 );
not ( n12492 , n12491 );
not ( n12493 , n12492 );
or ( n12494 , n12490 , n12493 );
not ( n12495 , n12488 );
buf ( n12496 , n12491 );
nand ( n12497 , n12495 , n12496 );
nand ( n12498 , n12494 , n12497 );
not ( n12499 , n12498 );
xor ( n12500 , n12487 , n12499 );
buf ( n12501 , n5310 );
not ( n12502 , n12501 );
buf ( n12503 , n5311 );
nand ( n12504 , n6622 , n12503 );
buf ( n12505 , n5312 );
buf ( n12506 , n12505 );
and ( n12507 , n12504 , n12506 );
not ( n12508 , n12504 );
not ( n12509 , n12505 );
and ( n12510 , n12508 , n12509 );
nor ( n12511 , n12507 , n12510 );
not ( n12512 , n12511 );
or ( n12513 , n12502 , n12512 );
or ( n12514 , n12511 , n12501 );
nand ( n12515 , n12513 , n12514 );
xnor ( n12516 , n12500 , n12515 );
not ( n12517 , n12516 );
buf ( n12518 , n5313 );
buf ( n12519 , n12518 );
not ( n12520 , n12519 );
and ( n12521 , n12517 , n12520 );
buf ( n12522 , n12486 );
xor ( n12523 , n12522 , n12498 );
xnor ( n12524 , n12523 , n12515 );
buf ( n12525 , n12524 );
and ( n12526 , n12525 , n12519 );
nor ( n12527 , n12521 , n12526 );
not ( n12528 , n8678 );
not ( n12529 , n8702 );
or ( n12530 , n12528 , n12529 );
nand ( n12531 , n12530 , n8706 );
not ( n12532 , n12531 );
and ( n12533 , n12527 , n12532 );
not ( n12534 , n12527 );
and ( n12535 , n12534 , n12531 );
nor ( n12536 , n12533 , n12535 );
not ( n12537 , n12536 );
and ( n12538 , n12485 , n12537 );
and ( n12539 , n12484 , n12536 );
nor ( n12540 , n12538 , n12539 );
and ( n12541 , n12381 , n12540 );
not ( n12542 , n12381 );
not ( n12543 , n12540 );
and ( n12544 , n12542 , n12543 );
nor ( n12545 , n12541 , n12544 );
buf ( n12546 , n12545 );
not ( n12547 , n12546 );
buf ( n12548 , n11318 );
xor ( n12549 , n8056 , n12548 );
buf ( n12550 , n5314 );
not ( n12551 , n12550 );
buf ( n12552 , n5315 );
not ( n12553 , n12552 );
buf ( n12554 , n5316 );
buf ( n12555 , n12554 );
and ( n12556 , n12553 , n12555 );
not ( n12557 , n12553 );
not ( n12558 , n12554 );
and ( n12559 , n12557 , n12558 );
nor ( n12560 , n12556 , n12559 );
xor ( n12561 , n12551 , n12560 );
buf ( n12562 , n5317 );
nand ( n12563 , n7981 , n12562 );
buf ( n12564 , n5318 );
buf ( n12565 , n12564 );
and ( n12566 , n12563 , n12565 );
not ( n12567 , n12563 );
not ( n12568 , n12564 );
and ( n12569 , n12567 , n12568 );
nor ( n12570 , n12566 , n12569 );
not ( n12571 , n12570 );
buf ( n12572 , n5319 );
nand ( n12573 , n8344 , n12572 );
buf ( n12574 , n5320 );
not ( n12575 , n12574 );
and ( n12576 , n12573 , n12575 );
not ( n12577 , n12573 );
buf ( n12578 , n12574 );
and ( n12579 , n12577 , n12578 );
nor ( n12580 , n12576 , n12579 );
not ( n12581 , n12580 );
or ( n12582 , n12571 , n12581 );
not ( n12583 , n12580 );
not ( n12584 , n12570 );
nand ( n12585 , n12583 , n12584 );
nand ( n12586 , n12582 , n12585 );
xnor ( n12587 , n12561 , n12586 );
xnor ( n12588 , n12549 , n12587 );
buf ( n12589 , n5321 );
not ( n12590 , n12589 );
not ( n12591 , n8665 );
not ( n12592 , n12591 );
not ( n12593 , n12592 );
or ( n12594 , n12590 , n12593 );
not ( n12595 , n12589 );
nand ( n12596 , n12595 , n12591 );
nand ( n12597 , n12594 , n12596 );
buf ( n12598 , n5322 );
buf ( n12599 , n12598 );
not ( n12600 , n12599 );
buf ( n12601 , n5323 );
not ( n12602 , n12601 );
not ( n12603 , n12602 );
or ( n12604 , n12600 , n12603 );
not ( n12605 , n12598 );
buf ( n12606 , n12601 );
nand ( n12607 , n12605 , n12606 );
nand ( n12608 , n12604 , n12607 );
buf ( n12609 , n5324 );
not ( n12610 , n12609 );
and ( n12611 , n12608 , n12610 );
not ( n12612 , n12608 );
buf ( n12613 , n12609 );
and ( n12614 , n12612 , n12613 );
nor ( n12615 , n12611 , n12614 );
buf ( n12616 , n5325 );
nand ( n12617 , n7909 , n12616 );
buf ( n12618 , n5326 );
buf ( n12619 , n12618 );
and ( n12620 , n12617 , n12619 );
not ( n12621 , n12617 );
not ( n12622 , n12618 );
and ( n12623 , n12621 , n12622 );
nor ( n12624 , n12620 , n12623 );
xor ( n12625 , n12615 , n12624 );
buf ( n12626 , n5327 );
nand ( n12627 , n7442 , n12626 );
buf ( n12628 , n5328 );
buf ( n12629 , n12628 );
and ( n12630 , n12627 , n12629 );
not ( n12631 , n12627 );
not ( n12632 , n12628 );
and ( n12633 , n12631 , n12632 );
nor ( n12634 , n12630 , n12633 );
xnor ( n12635 , n12625 , n12634 );
not ( n12636 , n12635 );
not ( n12637 , n12636 );
and ( n12638 , n12597 , n12637 );
not ( n12639 , n12597 );
buf ( n12640 , n12635 );
not ( n12641 , n12640 );
and ( n12642 , n12639 , n12641 );
nor ( n12643 , n12638 , n12642 );
nand ( n12644 , n12588 , n12643 );
not ( n12645 , n12644 );
buf ( n12646 , n5329 );
buf ( n12647 , n12646 );
not ( n12648 , n12647 );
buf ( n12649 , n5330 );
not ( n12650 , n12649 );
not ( n12651 , n12650 );
or ( n12652 , n12648 , n12651 );
not ( n12653 , n12646 );
buf ( n12654 , n12649 );
nand ( n12655 , n12653 , n12654 );
nand ( n12656 , n12652 , n12655 );
buf ( n12657 , n5331 );
not ( n12658 , n12657 );
and ( n12659 , n12656 , n12658 );
not ( n12660 , n12656 );
buf ( n12661 , n12657 );
and ( n12662 , n12660 , n12661 );
nor ( n12663 , n12659 , n12662 );
buf ( n12664 , n5332 );
nand ( n12665 , n8387 , n12664 );
buf ( n12666 , n5333 );
buf ( n12667 , n12666 );
and ( n12668 , n12665 , n12667 );
not ( n12669 , n12665 );
not ( n12670 , n12666 );
and ( n12671 , n12669 , n12670 );
nor ( n12672 , n12668 , n12671 );
xor ( n12673 , n12663 , n12672 );
buf ( n12674 , n5334 );
nand ( n12675 , n8971 , n12674 );
buf ( n12676 , n5335 );
buf ( n12677 , n12676 );
and ( n12678 , n12675 , n12677 );
not ( n12679 , n12675 );
not ( n12680 , n12676 );
and ( n12681 , n12679 , n12680 );
nor ( n12682 , n12678 , n12681 );
xnor ( n12683 , n12673 , n12682 );
not ( n12684 , n12683 );
not ( n12685 , n12684 );
not ( n12686 , n12685 );
not ( n12687 , n12686 );
buf ( n12688 , n5336 );
not ( n12689 , n12688 );
not ( n12690 , n12689 );
buf ( n12691 , n5337 );
buf ( n12692 , n12691 );
not ( n12693 , n12692 );
buf ( n12694 , n5338 );
not ( n12695 , n12694 );
not ( n12696 , n12695 );
or ( n12697 , n12693 , n12696 );
not ( n12698 , n12691 );
buf ( n12699 , n12694 );
nand ( n12700 , n12698 , n12699 );
nand ( n12701 , n12697 , n12700 );
buf ( n12702 , n5339 );
not ( n12703 , n12702 );
and ( n12704 , n12701 , n12703 );
not ( n12705 , n12701 );
buf ( n12706 , n12702 );
and ( n12707 , n12705 , n12706 );
nor ( n12708 , n12704 , n12707 );
buf ( n12709 , n5340 );
nand ( n12710 , n7865 , n12709 );
buf ( n12711 , n5341 );
buf ( n12712 , n12711 );
and ( n12713 , n12710 , n12712 );
not ( n12714 , n12710 );
not ( n12715 , n12711 );
and ( n12716 , n12714 , n12715 );
nor ( n12717 , n12713 , n12716 );
not ( n12718 , n12717 );
xor ( n12719 , n12708 , n12718 );
buf ( n12720 , n5342 );
nand ( n12721 , n6851 , n12720 );
buf ( n12722 , n5343 );
not ( n12723 , n12722 );
and ( n12724 , n12721 , n12723 );
not ( n12725 , n12721 );
buf ( n12726 , n12722 );
and ( n12727 , n12725 , n12726 );
nor ( n12728 , n12724 , n12727 );
buf ( n12729 , n12728 );
xnor ( n12730 , n12719 , n12729 );
not ( n12731 , n12730 );
or ( n12732 , n12690 , n12731 );
not ( n12733 , n12689 );
not ( n12734 , n12717 );
not ( n12735 , n12728 );
or ( n12736 , n12734 , n12735 );
or ( n12737 , n12717 , n12728 );
nand ( n12738 , n12736 , n12737 );
and ( n12739 , n12738 , n12708 );
not ( n12740 , n12738 );
not ( n12741 , n12708 );
and ( n12742 , n12740 , n12741 );
nor ( n12743 , n12739 , n12742 );
nand ( n12744 , n12733 , n12743 );
nand ( n12745 , n12732 , n12744 );
not ( n12746 , n12745 );
or ( n12747 , n12687 , n12746 );
not ( n12748 , n12683 );
buf ( n12749 , n12748 );
or ( n12750 , n12745 , n12749 );
nand ( n12751 , n12747 , n12750 );
buf ( n12752 , n12751 );
not ( n12753 , n12752 );
and ( n12754 , n12645 , n12753 );
not ( n12755 , n12643 );
not ( n12756 , n12755 );
nand ( n12757 , n12756 , n12588 );
and ( n12758 , n12757 , n12752 );
nor ( n12759 , n12754 , n12758 );
not ( n12760 , n12759 );
not ( n12761 , n12760 );
nand ( n12762 , n11925 , n11779 );
buf ( n12763 , n5344 );
buf ( n12764 , n12763 );
not ( n12765 , n12764 );
buf ( n12766 , n5345 );
buf ( n12767 , n12766 );
not ( n12768 , n12767 );
buf ( n12769 , n5346 );
not ( n12770 , n12769 );
not ( n12771 , n12770 );
or ( n12772 , n12768 , n12771 );
not ( n12773 , n12766 );
buf ( n12774 , n12769 );
nand ( n12775 , n12773 , n12774 );
nand ( n12776 , n12772 , n12775 );
buf ( n12777 , n5347 );
not ( n12778 , n12777 );
and ( n12779 , n12776 , n12778 );
not ( n12780 , n12776 );
buf ( n12781 , n12777 );
and ( n12782 , n12780 , n12781 );
nor ( n12783 , n12779 , n12782 );
buf ( n12784 , n5348 );
nand ( n12785 , n7412 , n12784 );
buf ( n12786 , n5349 );
not ( n12787 , n12786 );
and ( n12788 , n12785 , n12787 );
not ( n12789 , n12785 );
buf ( n12790 , n12786 );
and ( n12791 , n12789 , n12790 );
nor ( n12792 , n12788 , n12791 );
xor ( n12793 , n12783 , n12792 );
buf ( n12794 , n5350 );
nand ( n12795 , n7356 , n12794 );
buf ( n12796 , n5351 );
not ( n12797 , n12796 );
and ( n12798 , n12795 , n12797 );
not ( n12799 , n12795 );
buf ( n12800 , n12796 );
and ( n12801 , n12799 , n12800 );
nor ( n12802 , n12798 , n12801 );
xnor ( n12803 , n12793 , n12802 );
not ( n12804 , n12803 );
not ( n12805 , n12804 );
or ( n12806 , n12765 , n12805 );
not ( n12807 , n12804 );
not ( n12808 , n12763 );
nand ( n12809 , n12807 , n12808 );
nand ( n12810 , n12806 , n12809 );
and ( n12811 , n12810 , n7755 );
not ( n12812 , n12810 );
and ( n12813 , n12812 , n7756 );
nor ( n12814 , n12811 , n12813 );
not ( n12815 , n12814 );
and ( n12816 , n12762 , n12815 );
not ( n12817 , n12762 );
and ( n12818 , n12817 , n12814 );
nor ( n12819 , n12816 , n12818 );
not ( n12820 , n12819 );
not ( n12821 , n12820 );
or ( n12822 , n12761 , n12821 );
nand ( n12823 , n12819 , n12759 );
nand ( n12824 , n12822 , n12823 );
not ( n12825 , n12824 );
or ( n12826 , n12547 , n12825 );
or ( n12827 , n12824 , n12546 );
nand ( n12828 , n12826 , n12827 );
not ( n12829 , n12828 );
or ( n12830 , n11932 , n12829 );
not ( n12831 , n11931 );
xor ( n12832 , n12824 , n12545 );
nand ( n12833 , n12831 , n12832 );
nand ( n12834 , n12830 , n12833 );
buf ( n12835 , n5352 );
not ( n12836 , n12835 );
buf ( n12837 , n5353 );
buf ( n12838 , n12837 );
and ( n12839 , n12836 , n12838 );
not ( n12840 , n12836 );
not ( n12841 , n12837 );
and ( n12842 , n12840 , n12841 );
nor ( n12843 , n12839 , n12842 );
not ( n12844 , n12843 );
buf ( n12845 , n5354 );
buf ( n12846 , n12845 );
not ( n12847 , n12846 );
and ( n12848 , n12844 , n12847 );
and ( n12849 , n12843 , n12846 );
nor ( n12850 , n12848 , n12849 );
not ( n12851 , n12850 );
buf ( n12852 , n5355 );
xor ( n12853 , n12852 , n12119 );
buf ( n12854 , n5356 );
nand ( n12855 , n10577 , n12854 );
buf ( n12856 , n5357 );
not ( n12857 , n12856 );
and ( n12858 , n12855 , n12857 );
not ( n12859 , n12855 );
buf ( n12860 , n12856 );
and ( n12861 , n12859 , n12860 );
nor ( n12862 , n12858 , n12861 );
xnor ( n12863 , n12853 , n12862 );
not ( n12864 , n12863 );
or ( n12865 , n12851 , n12864 );
or ( n12866 , n12863 , n12850 );
nand ( n12867 , n12865 , n12866 );
and ( n12868 , n12867 , n10589 );
not ( n12869 , n12867 );
buf ( n12870 , n10588 );
and ( n12871 , n12869 , n12870 );
nor ( n12872 , n12868 , n12871 );
buf ( n12873 , n5358 );
not ( n12874 , n12873 );
buf ( n12875 , n5359 );
not ( n12876 , n12875 );
buf ( n12877 , n5360 );
buf ( n12878 , n12877 );
nand ( n12879 , n12876 , n12878 );
not ( n12880 , n12877 );
buf ( n12881 , n12875 );
nand ( n12882 , n12880 , n12881 );
and ( n12883 , n12879 , n12882 );
xor ( n12884 , n12874 , n12883 );
buf ( n12885 , n5361 );
nand ( n12886 , n6816 , n12885 );
buf ( n12887 , n5362 );
buf ( n12888 , n12887 );
and ( n12889 , n12886 , n12888 );
not ( n12890 , n12886 );
not ( n12891 , n12887 );
and ( n12892 , n12890 , n12891 );
nor ( n12893 , n12889 , n12892 );
not ( n12894 , n12893 );
buf ( n12895 , n5363 );
not ( n12896 , n12895 );
and ( n12897 , n12894 , n12896 );
and ( n12898 , n12893 , n12895 );
nor ( n12899 , n12897 , n12898 );
xnor ( n12900 , n12884 , n12899 );
not ( n12901 , n12900 );
not ( n12902 , n12901 );
buf ( n12903 , n5364 );
buf ( n12904 , n12903 );
not ( n12905 , n12904 );
buf ( n12906 , n5365 );
nand ( n12907 , n7865 , n12906 );
buf ( n12908 , n5366 );
buf ( n12909 , n12908 );
and ( n12910 , n12907 , n12909 );
not ( n12911 , n12907 );
not ( n12912 , n12908 );
and ( n12913 , n12911 , n12912 );
nor ( n12914 , n12910 , n12913 );
not ( n12915 , n12914 );
buf ( n12916 , n5367 );
nand ( n12917 , n7412 , n12916 );
buf ( n12918 , n5368 );
not ( n12919 , n12918 );
and ( n12920 , n12917 , n12919 );
not ( n12921 , n12917 );
buf ( n12922 , n12918 );
and ( n12923 , n12921 , n12922 );
nor ( n12924 , n12920 , n12923 );
not ( n12925 , n12924 );
or ( n12926 , n12915 , n12925 );
or ( n12927 , n12914 , n12924 );
nand ( n12928 , n12926 , n12927 );
buf ( n12929 , n5369 );
buf ( n12930 , n12929 );
not ( n12931 , n12930 );
buf ( n12932 , n5370 );
not ( n12933 , n12932 );
not ( n12934 , n12933 );
or ( n12935 , n12931 , n12934 );
not ( n12936 , n12929 );
buf ( n12937 , n12932 );
nand ( n12938 , n12936 , n12937 );
nand ( n12939 , n12935 , n12938 );
buf ( n12940 , n5371 );
not ( n12941 , n12940 );
and ( n12942 , n12939 , n12941 );
not ( n12943 , n12939 );
buf ( n12944 , n12940 );
and ( n12945 , n12943 , n12944 );
nor ( n12946 , n12942 , n12945 );
and ( n12947 , n12928 , n12946 );
not ( n12948 , n12928 );
not ( n12949 , n12946 );
and ( n12950 , n12948 , n12949 );
nor ( n12951 , n12947 , n12950 );
not ( n12952 , n12951 );
or ( n12953 , n12905 , n12952 );
or ( n12954 , n12951 , n12904 );
nand ( n12955 , n12953 , n12954 );
not ( n12956 , n12955 );
or ( n12957 , n12902 , n12956 );
buf ( n12958 , n12873 );
xor ( n12959 , n12958 , n12883 );
xor ( n12960 , n12959 , n12899 );
not ( n12961 , n12960 );
or ( n12962 , n12955 , n12961 );
nand ( n12963 , n12957 , n12962 );
nand ( n12964 , n12872 , n12963 );
not ( n12965 , n12964 );
not ( n12966 , n11057 );
buf ( n12967 , n5372 );
buf ( n12968 , n12967 );
not ( n12969 , n12968 );
buf ( n12970 , n5373 );
not ( n12971 , n12970 );
not ( n12972 , n12971 );
or ( n12973 , n12969 , n12972 );
not ( n12974 , n12967 );
buf ( n12975 , n12970 );
nand ( n12976 , n12974 , n12975 );
nand ( n12977 , n12973 , n12976 );
buf ( n12978 , n5374 );
buf ( n12979 , n12978 );
and ( n12980 , n12977 , n12979 );
not ( n12981 , n12977 );
not ( n12982 , n12978 );
and ( n12983 , n12981 , n12982 );
nor ( n12984 , n12980 , n12983 );
buf ( n12985 , n5375 );
nand ( n12986 , n6985 , n12985 );
buf ( n12987 , n5376 );
buf ( n12988 , n12987 );
and ( n12989 , n12986 , n12988 );
not ( n12990 , n12986 );
not ( n12991 , n12987 );
and ( n12992 , n12990 , n12991 );
nor ( n12993 , n12989 , n12992 );
not ( n12994 , n12993 );
xor ( n12995 , n12984 , n12994 );
buf ( n12996 , n5377 );
nand ( n12997 , n9619 , n12996 );
buf ( n12998 , n5378 );
not ( n12999 , n12998 );
and ( n13000 , n12997 , n12999 );
not ( n13001 , n12997 );
buf ( n13002 , n12998 );
and ( n13003 , n13001 , n13002 );
nor ( n13004 , n13000 , n13003 );
xnor ( n13005 , n12995 , n13004 );
not ( n13006 , n13005 );
or ( n13007 , n12966 , n13006 );
not ( n13008 , n11057 );
xor ( n13009 , n12984 , n12993 );
xnor ( n13010 , n13009 , n13004 );
nand ( n13011 , n13008 , n13010 );
nand ( n13012 , n13007 , n13011 );
and ( n13013 , n13012 , n7933 );
not ( n13014 , n13012 );
not ( n13015 , n7931 );
not ( n13016 , n13015 );
and ( n13017 , n13014 , n13016 );
nor ( n13018 , n13013 , n13017 );
not ( n13019 , n13018 );
not ( n13020 , n13019 );
and ( n13021 , n12965 , n13020 );
and ( n13022 , n12964 , n13019 );
nor ( n13023 , n13021 , n13022 );
not ( n13024 , n13023 );
buf ( n13025 , n5379 );
buf ( n13026 , n13025 );
not ( n13027 , n10613 );
xor ( n13028 , n10635 , n13027 );
buf ( n13029 , n10603 );
xnor ( n13030 , n13028 , n13029 );
xor ( n13031 , n13026 , n13030 );
not ( n13032 , n11542 );
xnor ( n13033 , n13031 , n13032 );
not ( n13034 , n13033 );
buf ( n13035 , n5380 );
buf ( n13036 , n13035 );
not ( n13037 , n13036 );
buf ( n13038 , n5381 );
not ( n13039 , n13038 );
buf ( n13040 , n5382 );
buf ( n13041 , n13040 );
and ( n13042 , n13039 , n13041 );
not ( n13043 , n13039 );
not ( n13044 , n13040 );
and ( n13045 , n13043 , n13044 );
nor ( n13046 , n13042 , n13045 );
not ( n13047 , n13046 );
or ( n13048 , n13037 , n13047 );
or ( n13049 , n13046 , n13036 );
nand ( n13050 , n13048 , n13049 );
not ( n13051 , n13050 );
buf ( n13052 , n5383 );
buf ( n13053 , n5384 );
not ( n13054 , n13053 );
xor ( n13055 , n13052 , n13054 );
buf ( n13056 , n5385 );
nand ( n13057 , n6905 , n13056 );
buf ( n13058 , n5386 );
not ( n13059 , n13058 );
and ( n13060 , n13057 , n13059 );
not ( n13061 , n13057 );
buf ( n13062 , n13058 );
and ( n13063 , n13061 , n13062 );
nor ( n13064 , n13060 , n13063 );
xnor ( n13065 , n13055 , n13064 );
not ( n13066 , n13065 );
not ( n13067 , n13066 );
or ( n13068 , n13051 , n13067 );
or ( n13069 , n13066 , n13050 );
nand ( n13070 , n13068 , n13069 );
not ( n13071 , n13070 );
buf ( n13072 , n11671 );
not ( n13073 , n13072 );
and ( n13074 , n13071 , n13073 );
and ( n13075 , n13070 , n11673 );
nor ( n13076 , n13074 , n13075 );
nand ( n13077 , n13034 , n13076 );
buf ( n13078 , n5387 );
buf ( n13079 , n13078 );
not ( n13080 , n13079 );
not ( n13081 , n8190 );
or ( n13082 , n13080 , n13081 );
not ( n13083 , n13078 );
nand ( n13084 , n8164 , n13083 );
nand ( n13085 , n13082 , n13084 );
not ( n13086 , n13085 );
buf ( n13087 , n8186 );
not ( n13088 , n13087 );
or ( n13089 , n13086 , n13088 );
or ( n13090 , n13087 , n13085 );
nand ( n13091 , n13089 , n13090 );
buf ( n13092 , n5388 );
buf ( n13093 , n13092 );
not ( n13094 , n13093 );
buf ( n13095 , n5389 );
not ( n13096 , n13095 );
not ( n13097 , n13096 );
or ( n13098 , n13094 , n13097 );
not ( n13099 , n13092 );
buf ( n13100 , n13095 );
nand ( n13101 , n13099 , n13100 );
nand ( n13102 , n13098 , n13101 );
buf ( n13103 , n5390 );
not ( n13104 , n13103 );
and ( n13105 , n13102 , n13104 );
not ( n13106 , n13102 );
buf ( n13107 , n13103 );
and ( n13108 , n13106 , n13107 );
nor ( n13109 , n13105 , n13108 );
xor ( n13110 , n13109 , n8353 );
buf ( n13111 , n5391 );
nand ( n13112 , n7617 , n13111 );
buf ( n13113 , n5392 );
not ( n13114 , n13113 );
and ( n13115 , n13112 , n13114 );
not ( n13116 , n13112 );
buf ( n13117 , n13113 );
and ( n13118 , n13116 , n13117 );
nor ( n13119 , n13115 , n13118 );
xnor ( n13120 , n13110 , n13119 );
buf ( n13121 , n13120 );
and ( n13122 , n13091 , n13121 );
not ( n13123 , n13091 );
xor ( n13124 , n13109 , n8353 );
xor ( n13125 , n13124 , n13119 );
and ( n13126 , n13123 , n13125 );
nor ( n13127 , n13122 , n13126 );
and ( n13128 , n13077 , n13127 );
not ( n13129 , n13077 );
not ( n13130 , n13127 );
and ( n13131 , n13129 , n13130 );
nor ( n13132 , n13128 , n13131 );
not ( n13133 , n13132 );
or ( n13134 , n13024 , n13133 );
or ( n13135 , n13132 , n13023 );
nand ( n13136 , n13134 , n13135 );
not ( n13137 , n7114 );
buf ( n13138 , n5393 );
not ( n13139 , n13138 );
buf ( n13140 , n5394 );
not ( n13141 , n13140 );
buf ( n13142 , n5395 );
buf ( n13143 , n13142 );
nand ( n13144 , n13141 , n13143 );
not ( n13145 , n13142 );
buf ( n13146 , n13140 );
nand ( n13147 , n13145 , n13146 );
and ( n13148 , n13144 , n13147 );
xor ( n13149 , n13139 , n13148 );
buf ( n13150 , n5396 );
buf ( n13151 , n5397 );
not ( n13152 , n13151 );
xor ( n13153 , n13150 , n13152 );
buf ( n13154 , n5398 );
nand ( n13155 , n10577 , n13154 );
xnor ( n13156 , n13153 , n13155 );
xnor ( n13157 , n13149 , n13156 );
buf ( n13158 , n13157 );
not ( n13159 , n13158 );
or ( n13160 , n13137 , n13159 );
not ( n13161 , n7114 );
buf ( n13162 , n13138 );
xor ( n13163 , n13162 , n13148 );
xnor ( n13164 , n13163 , n13156 );
buf ( n13165 , n13164 );
nand ( n13166 , n13161 , n13165 );
nand ( n13167 , n13160 , n13166 );
buf ( n13168 , n5399 );
buf ( n13169 , n13168 );
not ( n13170 , n13169 );
buf ( n13171 , n5400 );
not ( n13172 , n13171 );
not ( n13173 , n13172 );
or ( n13174 , n13170 , n13173 );
not ( n13175 , n13168 );
buf ( n13176 , n13171 );
nand ( n13177 , n13175 , n13176 );
nand ( n13178 , n13174 , n13177 );
not ( n13179 , n13178 );
buf ( n13180 , n5401 );
nand ( n13181 , n6863 , n13180 );
buf ( n13182 , n5402 );
buf ( n13183 , n13182 );
and ( n13184 , n13181 , n13183 );
not ( n13185 , n13181 );
not ( n13186 , n13182 );
and ( n13187 , n13185 , n13186 );
nor ( n13188 , n13184 , n13187 );
not ( n13189 , n13188 );
buf ( n13190 , n5403 );
nand ( n13191 , n6760 , n13190 );
buf ( n13192 , n5404 );
buf ( n13193 , n13192 );
and ( n13194 , n13191 , n13193 );
not ( n13195 , n13191 );
not ( n13196 , n13192 );
and ( n13197 , n13195 , n13196 );
nor ( n13198 , n13194 , n13197 );
not ( n13199 , n13198 );
not ( n13200 , n13199 );
or ( n13201 , n13189 , n13200 );
not ( n13202 , n13188 );
nand ( n13203 , n13198 , n13202 );
nand ( n13204 , n13201 , n13203 );
buf ( n13205 , n5405 );
buf ( n13206 , n13205 );
and ( n13207 , n13204 , n13206 );
not ( n13208 , n13204 );
not ( n13209 , n13205 );
and ( n13210 , n13208 , n13209 );
nor ( n13211 , n13207 , n13210 );
not ( n13212 , n13211 );
not ( n13213 , n13212 );
or ( n13214 , n13179 , n13213 );
not ( n13215 , n13178 );
nand ( n13216 , n13211 , n13215 );
nand ( n13217 , n13214 , n13216 );
buf ( n13218 , n13217 );
and ( n13219 , n13167 , n13218 );
not ( n13220 , n13167 );
xor ( n13221 , n13206 , n13178 );
xnor ( n13222 , n13221 , n13204 );
buf ( n13223 , n13222 );
and ( n13224 , n13220 , n13223 );
nor ( n13225 , n13219 , n13224 );
not ( n13226 , n9233 );
xor ( n13227 , n11614 , n11618 );
xnor ( n13228 , n13227 , n11628 );
buf ( n13229 , n13228 );
not ( n13230 , n13229 );
or ( n13231 , n13226 , n13230 );
buf ( n13232 , n11629 );
nand ( n13233 , n13232 , n9229 );
nand ( n13234 , n13231 , n13233 );
not ( n13235 , n13234 );
not ( n13236 , n11592 );
buf ( n13237 , n13236 );
not ( n13238 , n13237 );
and ( n13239 , n13235 , n13238 );
and ( n13240 , n13234 , n13237 );
nor ( n13241 , n13239 , n13240 );
nand ( n13242 , n13225 , n13241 );
not ( n13243 , n13242 );
not ( n13244 , n7756 );
buf ( n13245 , n5406 );
nand ( n13246 , n6660 , n13245 );
buf ( n13247 , n5407 );
not ( n13248 , n13247 );
and ( n13249 , n13246 , n13248 );
not ( n13250 , n13246 );
buf ( n13251 , n13247 );
and ( n13252 , n13250 , n13251 );
nor ( n13253 , n13249 , n13252 );
buf ( n13254 , n13253 );
not ( n13255 , n13254 );
buf ( n13256 , n12803 );
not ( n13257 , n13256 );
not ( n13258 , n13257 );
or ( n13259 , n13255 , n13258 );
not ( n13260 , n13254 );
nand ( n13261 , n13260 , n12807 );
nand ( n13262 , n13259 , n13261 );
not ( n13263 , n13262 );
or ( n13264 , n13244 , n13263 );
or ( n13265 , n7756 , n13262 );
nand ( n13266 , n13264 , n13265 );
not ( n13267 , n13266 );
and ( n13268 , n13243 , n13267 );
and ( n13269 , n13242 , n13266 );
nor ( n13270 , n13268 , n13269 );
and ( n13271 , n13136 , n13270 );
not ( n13272 , n13136 );
not ( n13273 , n13270 );
and ( n13274 , n13272 , n13273 );
nor ( n13275 , n13271 , n13274 );
not ( n13276 , n13275 );
not ( n13277 , n13276 );
buf ( n13278 , n5408 );
buf ( n13279 , n13278 );
not ( n13280 , n13279 );
buf ( n13281 , n5409 );
buf ( n13282 , n13281 );
not ( n13283 , n13282 );
buf ( n13284 , n5410 );
not ( n13285 , n13284 );
not ( n13286 , n13285 );
or ( n13287 , n13283 , n13286 );
not ( n13288 , n13281 );
buf ( n13289 , n13284 );
nand ( n13290 , n13288 , n13289 );
nand ( n13291 , n13287 , n13290 );
buf ( n13292 , n5411 );
buf ( n13293 , n13292 );
and ( n13294 , n13291 , n13293 );
not ( n13295 , n13291 );
not ( n13296 , n13292 );
and ( n13297 , n13295 , n13296 );
nor ( n13298 , n13294 , n13297 );
buf ( n13299 , n5412 );
nand ( n13300 , n6706 , n13299 );
buf ( n13301 , n5413 );
buf ( n13302 , n13301 );
and ( n13303 , n13300 , n13302 );
not ( n13304 , n13300 );
not ( n13305 , n13301 );
and ( n13306 , n13304 , n13305 );
nor ( n13307 , n13303 , n13306 );
xor ( n13308 , n13298 , n13307 );
buf ( n13309 , n5414 );
nand ( n13310 , n6622 , n13309 );
buf ( n13311 , n5415 );
buf ( n13312 , n13311 );
and ( n13313 , n13310 , n13312 );
not ( n13314 , n13310 );
not ( n13315 , n13311 );
and ( n13316 , n13314 , n13315 );
nor ( n13317 , n13313 , n13316 );
not ( n13318 , n13317 );
xnor ( n13319 , n13308 , n13318 );
not ( n13320 , n13319 );
not ( n13321 , n13320 );
or ( n13322 , n13280 , n13321 );
not ( n13323 , n13279 );
not ( n13324 , n13320 );
nand ( n13325 , n13323 , n13324 );
nand ( n13326 , n13322 , n13325 );
not ( n13327 , n13326 );
buf ( n13328 , n5416 );
buf ( n13329 , n5417 );
not ( n13330 , n13329 );
buf ( n13331 , n5418 );
buf ( n13332 , n13331 );
and ( n13333 , n13330 , n13332 );
not ( n13334 , n13330 );
not ( n13335 , n13331 );
and ( n13336 , n13334 , n13335 );
nor ( n13337 , n13333 , n13336 );
xor ( n13338 , n13328 , n13337 );
buf ( n13339 , n5419 );
xor ( n13340 , n13339 , n11881 );
xnor ( n13341 , n13340 , n11876 );
xnor ( n13342 , n13338 , n13341 );
not ( n13343 , n13342 );
not ( n13344 , n13343 );
and ( n13345 , n13327 , n13344 );
and ( n13346 , n13326 , n13343 );
nor ( n13347 , n13345 , n13346 );
buf ( n13348 , n5420 );
buf ( n13349 , n13348 );
not ( n13350 , n13349 );
buf ( n13351 , n5421 );
buf ( n13352 , n13351 );
not ( n13353 , n13352 );
buf ( n13354 , n5422 );
not ( n13355 , n13354 );
not ( n13356 , n13355 );
or ( n13357 , n13353 , n13356 );
not ( n13358 , n13351 );
buf ( n13359 , n13354 );
nand ( n13360 , n13358 , n13359 );
nand ( n13361 , n13357 , n13360 );
buf ( n13362 , n5423 );
not ( n13363 , n13362 );
and ( n13364 , n13361 , n13363 );
not ( n13365 , n13361 );
buf ( n13366 , n13362 );
and ( n13367 , n13365 , n13366 );
nor ( n13368 , n13364 , n13367 );
buf ( n13369 , n5424 );
nand ( n13370 , n6934 , n13369 );
buf ( n13371 , n5425 );
buf ( n13372 , n13371 );
and ( n13373 , n13370 , n13372 );
not ( n13374 , n13370 );
not ( n13375 , n13371 );
and ( n13376 , n13374 , n13375 );
nor ( n13377 , n13373 , n13376 );
xor ( n13378 , n13368 , n13377 );
buf ( n13379 , n6660 );
buf ( n13380 , n5426 );
nand ( n13381 , n13379 , n13380 );
buf ( n13382 , n5427 );
not ( n13383 , n13382 );
and ( n13384 , n13381 , n13383 );
not ( n13385 , n13381 );
buf ( n13386 , n13382 );
and ( n13387 , n13385 , n13386 );
nor ( n13388 , n13384 , n13387 );
xnor ( n13389 , n13378 , n13388 );
buf ( n13390 , n13389 );
buf ( n13391 , n13390 );
not ( n13392 , n13391 );
or ( n13393 , n13350 , n13392 );
not ( n13394 , n13349 );
not ( n13395 , n13389 );
buf ( n13396 , n13395 );
nand ( n13397 , n13394 , n13396 );
nand ( n13398 , n13393 , n13397 );
buf ( n13399 , n11823 );
not ( n13400 , n13399 );
and ( n13401 , n13398 , n13400 );
not ( n13402 , n13398 );
buf ( n13403 , n11822 );
not ( n13404 , n13403 );
and ( n13405 , n13402 , n13404 );
nor ( n13406 , n13401 , n13405 );
nand ( n13407 , n13347 , n13406 );
not ( n13408 , n13407 );
buf ( n13409 , n5428 );
nand ( n13410 , n7442 , n13409 );
buf ( n13411 , n5429 );
not ( n13412 , n13411 );
and ( n13413 , n13410 , n13412 );
not ( n13414 , n13410 );
buf ( n13415 , n13411 );
and ( n13416 , n13414 , n13415 );
nor ( n13417 , n13413 , n13416 );
buf ( n13418 , n5430 );
buf ( n13419 , n13418 );
not ( n13420 , n13419 );
buf ( n13421 , n5431 );
not ( n13422 , n13421 );
not ( n13423 , n13422 );
or ( n13424 , n13420 , n13423 );
not ( n13425 , n13418 );
buf ( n13426 , n13421 );
nand ( n13427 , n13425 , n13426 );
nand ( n13428 , n13424 , n13427 );
buf ( n13429 , n5432 );
buf ( n13430 , n13429 );
and ( n13431 , n13428 , n13430 );
not ( n13432 , n13428 );
not ( n13433 , n13429 );
and ( n13434 , n13432 , n13433 );
nor ( n13435 , n13431 , n13434 );
buf ( n13436 , n5433 );
nand ( n13437 , n7299 , n13436 );
buf ( n13438 , n5434 );
buf ( n13439 , n13438 );
and ( n13440 , n13437 , n13439 );
not ( n13441 , n13437 );
not ( n13442 , n13438 );
and ( n13443 , n13441 , n13442 );
nor ( n13444 , n13440 , n13443 );
xor ( n13445 , n13435 , n13444 );
buf ( n13446 , n5435 );
nand ( n13447 , n6622 , n13446 );
buf ( n13448 , n5436 );
buf ( n13449 , n13448 );
and ( n13450 , n13447 , n13449 );
not ( n13451 , n13447 );
not ( n13452 , n13448 );
and ( n13453 , n13451 , n13452 );
nor ( n13454 , n13450 , n13453 );
not ( n13455 , n13454 );
xnor ( n13456 , n13445 , n13455 );
not ( n13457 , n13456 );
not ( n13458 , n13457 );
not ( n13459 , n13458 );
xor ( n13460 , n13417 , n13459 );
not ( n13461 , n11385 );
buf ( n13462 , n5437 );
not ( n13463 , n13462 );
not ( n13464 , n13463 );
or ( n13465 , n13461 , n13464 );
not ( n13466 , n11384 );
buf ( n13467 , n13462 );
nand ( n13468 , n13466 , n13467 );
nand ( n13469 , n13465 , n13468 );
not ( n13470 , n13469 );
buf ( n13471 , n5438 );
not ( n13472 , n13471 );
buf ( n13473 , n5439 );
nand ( n13474 , n6760 , n13473 );
not ( n13475 , n13474 );
buf ( n13476 , n5440 );
not ( n13477 , n13476 );
and ( n13478 , n13475 , n13477 );
nand ( n13479 , n6863 , n13473 );
and ( n13480 , n13479 , n13476 );
nor ( n13481 , n13478 , n13480 );
xor ( n13482 , n13472 , n13481 );
buf ( n13483 , n5441 );
nand ( n13484 , n6934 , n13483 );
not ( n13485 , n13484 );
buf ( n13486 , n5442 );
not ( n13487 , n13486 );
and ( n13488 , n13485 , n13487 );
nand ( n13489 , n7921 , n13483 );
and ( n13490 , n13489 , n13486 );
nor ( n13491 , n13488 , n13490 );
xnor ( n13492 , n13482 , n13491 );
not ( n13493 , n13492 );
not ( n13494 , n13493 );
or ( n13495 , n13470 , n13494 );
not ( n13496 , n13469 );
nand ( n13497 , n13496 , n13492 );
nand ( n13498 , n13495 , n13497 );
buf ( n13499 , n13498 );
not ( n13500 , n13499 );
xnor ( n13501 , n13460 , n13500 );
not ( n13502 , n13501 );
not ( n13503 , n13502 );
or ( n13504 , n13408 , n13503 );
or ( n13505 , n13502 , n13407 );
nand ( n13506 , n13504 , n13505 );
not ( n13507 , n13506 );
not ( n13508 , n13507 );
buf ( n13509 , n5443 );
buf ( n13510 , n13509 );
not ( n13511 , n13510 );
buf ( n13512 , n5444 );
not ( n13513 , n13512 );
not ( n13514 , n13513 );
or ( n13515 , n13511 , n13514 );
not ( n13516 , n13509 );
buf ( n13517 , n13512 );
nand ( n13518 , n13516 , n13517 );
nand ( n13519 , n13515 , n13518 );
buf ( n13520 , n5445 );
not ( n13521 , n13520 );
and ( n13522 , n13519 , n13521 );
not ( n13523 , n13519 );
buf ( n13524 , n13520 );
and ( n13525 , n13523 , n13524 );
nor ( n13526 , n13522 , n13525 );
buf ( n13527 , n5446 );
nand ( n13528 , n6863 , n13527 );
buf ( n13529 , n5447 );
buf ( n13530 , n13529 );
and ( n13531 , n13528 , n13530 );
not ( n13532 , n13528 );
not ( n13533 , n13529 );
and ( n13534 , n13532 , n13533 );
nor ( n13535 , n13531 , n13534 );
xor ( n13536 , n13526 , n13535 );
buf ( n13537 , n5448 );
nand ( n13538 , n6804 , n13537 );
buf ( n13539 , n5449 );
not ( n13540 , n13539 );
and ( n13541 , n13538 , n13540 );
not ( n13542 , n13538 );
buf ( n13543 , n13539 );
and ( n13544 , n13542 , n13543 );
nor ( n13545 , n13541 , n13544 );
xnor ( n13546 , n13536 , n13545 );
not ( n13547 , n13546 );
not ( n13548 , n13547 );
xor ( n13549 , n8529 , n13548 );
buf ( n13550 , n5450 );
buf ( n13551 , n5451 );
buf ( n13552 , n13551 );
not ( n13553 , n13552 );
buf ( n13554 , n5452 );
not ( n13555 , n13554 );
not ( n13556 , n13555 );
or ( n13557 , n13553 , n13556 );
not ( n13558 , n13551 );
buf ( n13559 , n13554 );
nand ( n13560 , n13558 , n13559 );
nand ( n13561 , n13557 , n13560 );
xor ( n13562 , n13550 , n13561 );
buf ( n13563 , n5453 );
buf ( n13564 , n5454 );
buf ( n13565 , n13564 );
xor ( n13566 , n13563 , n13565 );
buf ( n13567 , n5455 );
nand ( n13568 , n7617 , n13567 );
xnor ( n13569 , n13566 , n13568 );
not ( n13570 , n13569 );
xnor ( n13571 , n13562 , n13570 );
buf ( n13572 , n13571 );
xnor ( n13573 , n13549 , n13572 );
not ( n13574 , n13573 );
not ( n13575 , n13574 );
buf ( n13576 , n7489 );
not ( n13577 , n13576 );
buf ( n13578 , n5456 );
buf ( n13579 , n13578 );
buf ( n13580 , n5457 );
buf ( n13581 , n13580 );
not ( n13582 , n13581 );
buf ( n13583 , n5458 );
not ( n13584 , n13583 );
not ( n13585 , n13584 );
or ( n13586 , n13582 , n13585 );
not ( n13587 , n13580 );
buf ( n13588 , n13583 );
nand ( n13589 , n13587 , n13588 );
nand ( n13590 , n13586 , n13589 );
buf ( n13591 , n5459 );
buf ( n13592 , n13591 );
and ( n13593 , n13590 , n13592 );
not ( n13594 , n13590 );
not ( n13595 , n13591 );
and ( n13596 , n13594 , n13595 );
nor ( n13597 , n13593 , n13596 );
buf ( n13598 , n5460 );
nand ( n13599 , n6660 , n13598 );
buf ( n13600 , n5461 );
not ( n13601 , n13600 );
and ( n13602 , n13599 , n13601 );
not ( n13603 , n13599 );
buf ( n13604 , n13600 );
and ( n13605 , n13603 , n13604 );
nor ( n13606 , n13602 , n13605 );
xor ( n13607 , n13597 , n13606 );
buf ( n13608 , n5462 );
nand ( n13609 , n7082 , n13608 );
buf ( n13610 , n5463 );
not ( n13611 , n13610 );
and ( n13612 , n13609 , n13611 );
not ( n13613 , n13609 );
buf ( n13614 , n13610 );
and ( n13615 , n13613 , n13614 );
nor ( n13616 , n13612 , n13615 );
xor ( n13617 , n13607 , n13616 );
buf ( n13618 , n13617 );
xor ( n13619 , n13579 , n13618 );
not ( n13620 , n13619 );
or ( n13621 , n13577 , n13620 );
or ( n13622 , n13619 , n13576 );
nand ( n13623 , n13621 , n13622 );
not ( n13624 , n9568 );
buf ( n13625 , n5464 );
buf ( n13626 , n13625 );
not ( n13627 , n13626 );
buf ( n13628 , n5465 );
not ( n13629 , n13628 );
not ( n13630 , n13629 );
or ( n13631 , n13627 , n13630 );
not ( n13632 , n13625 );
buf ( n13633 , n13628 );
nand ( n13634 , n13632 , n13633 );
nand ( n13635 , n13631 , n13634 );
buf ( n13636 , n5466 );
not ( n13637 , n13636 );
and ( n13638 , n13635 , n13637 );
not ( n13639 , n13635 );
buf ( n13640 , n13636 );
and ( n13641 , n13639 , n13640 );
nor ( n13642 , n13638 , n13641 );
buf ( n13643 , n5467 );
nand ( n13644 , n8740 , n13643 );
buf ( n13645 , n5468 );
buf ( n13646 , n13645 );
and ( n13647 , n13644 , n13646 );
not ( n13648 , n13644 );
not ( n13649 , n13645 );
and ( n13650 , n13648 , n13649 );
nor ( n13651 , n13647 , n13650 );
xor ( n13652 , n13642 , n13651 );
buf ( n13653 , n5469 );
nand ( n13654 , n10107 , n13653 );
buf ( n13655 , n5470 );
buf ( n13656 , n13655 );
and ( n13657 , n13654 , n13656 );
not ( n13658 , n13654 );
not ( n13659 , n13655 );
and ( n13660 , n13658 , n13659 );
nor ( n13661 , n13657 , n13660 );
not ( n13662 , n13661 );
xnor ( n13663 , n13652 , n13662 );
not ( n13664 , n13663 );
or ( n13665 , n13624 , n13664 );
not ( n13666 , n13663 );
nand ( n13667 , n13666 , n9564 );
nand ( n13668 , n13665 , n13667 );
not ( n13669 , n13668 );
buf ( n13670 , n5471 );
buf ( n13671 , n13670 );
not ( n13672 , n13671 );
buf ( n13673 , n5472 );
not ( n13674 , n13673 );
not ( n13675 , n13674 );
or ( n13676 , n13672 , n13675 );
not ( n13677 , n13670 );
buf ( n13678 , n13673 );
nand ( n13679 , n13677 , n13678 );
nand ( n13680 , n13676 , n13679 );
buf ( n13681 , n5473 );
not ( n13682 , n13681 );
and ( n13683 , n13680 , n13682 );
not ( n13684 , n13680 );
buf ( n13685 , n13681 );
and ( n13686 , n13684 , n13685 );
nor ( n13687 , n13683 , n13686 );
buf ( n13688 , n5474 );
nand ( n13689 , n7750 , n13688 );
buf ( n13690 , n5475 );
buf ( n13691 , n13690 );
and ( n13692 , n13689 , n13691 );
not ( n13693 , n13689 );
not ( n13694 , n13690 );
and ( n13695 , n13693 , n13694 );
nor ( n13696 , n13692 , n13695 );
xor ( n13697 , n13687 , n13696 );
buf ( n13698 , n5476 );
nand ( n13699 , n8971 , n13698 );
buf ( n13700 , n5477 );
not ( n13701 , n13700 );
and ( n13702 , n13699 , n13701 );
not ( n13703 , n13699 );
buf ( n13704 , n13700 );
and ( n13705 , n13703 , n13704 );
nor ( n13706 , n13702 , n13705 );
xnor ( n13707 , n13697 , n13706 );
buf ( n13708 , n13707 );
buf ( n13709 , n13708 );
not ( n13710 , n13709 );
and ( n13711 , n13669 , n13710 );
and ( n13712 , n13668 , n13709 );
nor ( n13713 , n13711 , n13712 );
nor ( n13714 , n13623 , n13713 );
not ( n13715 , n13714 );
and ( n13716 , n13575 , n13715 );
and ( n13717 , n13574 , n13714 );
nor ( n13718 , n13716 , n13717 );
not ( n13719 , n13718 );
not ( n13720 , n13719 );
or ( n13721 , n13508 , n13720 );
nand ( n13722 , n13718 , n13506 );
nand ( n13723 , n13721 , n13722 );
not ( n13724 , n13723 );
not ( n13725 , n13724 );
or ( n13726 , n13277 , n13725 );
nand ( n13727 , n13275 , n13723 );
nand ( n13728 , n13726 , n13727 );
not ( n13729 , n13728 );
not ( n13730 , n13729 );
and ( n13731 , n12834 , n13730 );
not ( n13732 , n12834 );
buf ( n13733 , n13728 );
not ( n13734 , n13733 );
and ( n13735 , n13732 , n13734 );
nor ( n13736 , n13731 , n13735 );
buf ( n13737 , n9619 );
buf ( n13738 , n6601 );
nor ( n13739 , n13737 , n13738 );
buf ( n13740 , n5478 );
not ( n13741 , n13740 );
not ( n13742 , n13741 );
or ( n13743 , n13739 , n13742 );
buf ( n13744 , n13743 );
not ( n13745 , n13744 );
buf ( n13746 , n13745 );
not ( n13747 , n13746 );
nor ( n13748 , n13736 , n13747 );
not ( n13749 , n13748 );
or ( n13750 , n11754 , n13749 );
not ( n13751 , n13736 );
buf ( n13752 , n13743 );
buf ( n13753 , n13752 );
nor ( n13754 , n13751 , n13753 );
nand ( n13755 , n13754 , n11754 );
and ( n13756 , n13739 , n13741 );
buf ( n13757 , n13756 );
buf ( n13758 , n13757 );
buf ( n13759 , n5479 );
buf ( n13760 , n13759 );
nand ( n13761 , n13758 , n13760 );
nand ( n13762 , n13750 , n13755 , n13761 );
buf ( n13763 , n13762 );
buf ( n13764 , n13763 );
not ( n13765 , n12958 );
buf ( n13766 , n13756 );
buf ( n13767 , n13766 );
not ( n13768 , n13767 );
or ( n13769 , n13765 , n13768 );
buf ( n13770 , n5480 );
buf ( n13771 , n13770 );
not ( n13772 , n13771 );
buf ( n13773 , n5481 );
not ( n13774 , n13773 );
not ( n13775 , n13774 );
or ( n13776 , n13772 , n13775 );
not ( n13777 , n13770 );
buf ( n13778 , n13773 );
nand ( n13779 , n13777 , n13778 );
nand ( n13780 , n13776 , n13779 );
buf ( n13781 , n5482 );
buf ( n13782 , n13781 );
and ( n13783 , n13780 , n13782 );
not ( n13784 , n13780 );
not ( n13785 , n13781 );
and ( n13786 , n13784 , n13785 );
nor ( n13787 , n13783 , n13786 );
buf ( n13788 , n5483 );
nand ( n13789 , n6816 , n13788 );
buf ( n13790 , n5484 );
buf ( n13791 , n13790 );
and ( n13792 , n13789 , n13791 );
not ( n13793 , n13789 );
not ( n13794 , n13790 );
and ( n13795 , n13793 , n13794 );
nor ( n13796 , n13792 , n13795 );
xor ( n13797 , n13787 , n13796 );
xnor ( n13798 , n13797 , n7451 );
not ( n13799 , n13798 );
not ( n13800 , n13799 );
not ( n13801 , n11842 );
buf ( n13802 , n5485 );
buf ( n13803 , n13802 );
not ( n13804 , n13803 );
not ( n13805 , n13578 );
not ( n13806 , n13805 );
or ( n13807 , n13804 , n13806 );
not ( n13808 , n13802 );
nand ( n13809 , n13808 , n13579 );
nand ( n13810 , n13807 , n13809 );
buf ( n13811 , n5486 );
buf ( n13812 , n13811 );
and ( n13813 , n13810 , n13812 );
not ( n13814 , n13810 );
not ( n13815 , n13811 );
and ( n13816 , n13814 , n13815 );
nor ( n13817 , n13813 , n13816 );
buf ( n13818 , n5487 );
nand ( n13819 , n7183 , n13818 );
buf ( n13820 , n5488 );
buf ( n13821 , n13820 );
and ( n13822 , n13819 , n13821 );
not ( n13823 , n13819 );
not ( n13824 , n13820 );
and ( n13825 , n13823 , n13824 );
nor ( n13826 , n13822 , n13825 );
xor ( n13827 , n13817 , n13826 );
buf ( n13828 , n5489 );
nand ( n13829 , n7442 , n13828 );
buf ( n13830 , n5490 );
not ( n13831 , n13830 );
and ( n13832 , n13829 , n13831 );
not ( n13833 , n13829 );
buf ( n13834 , n13830 );
and ( n13835 , n13833 , n13834 );
nor ( n13836 , n13832 , n13835 );
xnor ( n13837 , n13827 , n13836 );
not ( n13838 , n13837 );
not ( n13839 , n13838 );
or ( n13840 , n13801 , n13839 );
xor ( n13841 , n13817 , n13826 );
xnor ( n13842 , n13841 , n13836 );
nand ( n13843 , n13842 , n11845 );
nand ( n13844 , n13840 , n13843 );
not ( n13845 , n13844 );
or ( n13846 , n13800 , n13845 );
or ( n13847 , n13844 , n13799 );
nand ( n13848 , n13846 , n13847 );
not ( n13849 , n13848 );
not ( n13850 , n10893 );
not ( n13851 , n6633 );
or ( n13852 , n13850 , n13851 );
or ( n13853 , n6638 , n10893 );
nand ( n13854 , n13852 , n13853 );
and ( n13855 , n13854 , n6678 );
not ( n13856 , n13854 );
buf ( n13857 , n6676 );
and ( n13858 , n13856 , n13857 );
or ( n13859 , n13855 , n13858 );
nand ( n13860 , n13849 , n13859 );
not ( n13861 , n13860 );
buf ( n13862 , n5491 );
buf ( n13863 , n13862 );
not ( n13864 , n13863 );
buf ( n13865 , n5492 );
buf ( n13866 , n13865 );
not ( n13867 , n13866 );
buf ( n13868 , n5493 );
not ( n13869 , n13868 );
not ( n13870 , n13869 );
or ( n13871 , n13867 , n13870 );
not ( n13872 , n13865 );
buf ( n13873 , n13868 );
nand ( n13874 , n13872 , n13873 );
nand ( n13875 , n13871 , n13874 );
buf ( n13876 , n5494 );
not ( n13877 , n13876 );
and ( n13878 , n13875 , n13877 );
not ( n13879 , n13875 );
buf ( n13880 , n13876 );
and ( n13881 , n13879 , n13880 );
nor ( n13882 , n13878 , n13881 );
buf ( n13883 , n5495 );
nand ( n13884 , n7043 , n13883 );
buf ( n13885 , n5496 );
buf ( n13886 , n13885 );
and ( n13887 , n13884 , n13886 );
not ( n13888 , n13884 );
not ( n13889 , n13885 );
and ( n13890 , n13888 , n13889 );
nor ( n13891 , n13887 , n13890 );
xor ( n13892 , n13882 , n13891 );
buf ( n13893 , n5497 );
nand ( n13894 , n6945 , n13893 );
buf ( n13895 , n5498 );
not ( n13896 , n13895 );
and ( n13897 , n13894 , n13896 );
not ( n13898 , n13894 );
buf ( n13899 , n13895 );
and ( n13900 , n13898 , n13899 );
nor ( n13901 , n13897 , n13900 );
xnor ( n13902 , n13892 , n13901 );
not ( n13903 , n13902 );
or ( n13904 , n13864 , n13903 );
or ( n13905 , n13902 , n13863 );
nand ( n13906 , n13904 , n13905 );
buf ( n13907 , n5499 );
buf ( n13908 , n13907 );
not ( n13909 , n13908 );
buf ( n13910 , n5500 );
not ( n13911 , n13910 );
not ( n13912 , n13911 );
or ( n13913 , n13909 , n13912 );
not ( n13914 , n13907 );
buf ( n13915 , n13910 );
nand ( n13916 , n13914 , n13915 );
nand ( n13917 , n13913 , n13916 );
buf ( n13918 , n5501 );
buf ( n13919 , n13918 );
and ( n13920 , n13917 , n13919 );
not ( n13921 , n13917 );
not ( n13922 , n13918 );
and ( n13923 , n13921 , n13922 );
nor ( n13924 , n13920 , n13923 );
buf ( n13925 , n5502 );
nand ( n13926 , n7616 , n13925 );
buf ( n13927 , n5503 );
buf ( n13928 , n13927 );
and ( n13929 , n13926 , n13928 );
not ( n13930 , n13926 );
not ( n13931 , n13927 );
and ( n13932 , n13930 , n13931 );
nor ( n13933 , n13929 , n13932 );
xor ( n13934 , n13924 , n13933 );
buf ( n13935 , n5504 );
nand ( n13936 , n7288 , n13935 );
buf ( n13937 , n5505 );
not ( n13938 , n13937 );
and ( n13939 , n13936 , n13938 );
not ( n13940 , n13936 );
buf ( n13941 , n13937 );
and ( n13942 , n13940 , n13941 );
nor ( n13943 , n13939 , n13942 );
xnor ( n13944 , n13934 , n13943 );
buf ( n13945 , n13944 );
not ( n13946 , n13945 );
and ( n13947 , n13906 , n13946 );
not ( n13948 , n13906 );
and ( n13949 , n13948 , n13945 );
nor ( n13950 , n13947 , n13949 );
not ( n13951 , n13950 );
not ( n13952 , n13951 );
and ( n13953 , n13861 , n13952 );
and ( n13954 , n13860 , n13951 );
nor ( n13955 , n13953 , n13954 );
not ( n13956 , n13955 );
not ( n13957 , n13956 );
nand ( n13958 , n13848 , n13950 );
not ( n13959 , n13958 );
buf ( n13960 , n5506 );
not ( n13961 , n13960 );
not ( n13962 , n13961 );
not ( n13963 , n9623 );
or ( n13964 , n13962 , n13963 );
not ( n13965 , n13961 );
nand ( n13966 , n13965 , n9629 );
nand ( n13967 , n13964 , n13966 );
buf ( n13968 , n5507 );
buf ( n13969 , n13968 );
not ( n13970 , n13969 );
buf ( n13971 , n5508 );
not ( n13972 , n13971 );
not ( n13973 , n13972 );
or ( n13974 , n13970 , n13973 );
not ( n13975 , n13968 );
buf ( n13976 , n13971 );
nand ( n13977 , n13975 , n13976 );
nand ( n13978 , n13974 , n13977 );
buf ( n13979 , n5509 );
not ( n13980 , n13979 );
and ( n13981 , n13978 , n13980 );
not ( n13982 , n13978 );
buf ( n13983 , n13979 );
and ( n13984 , n13982 , n13983 );
nor ( n13985 , n13981 , n13984 );
buf ( n13986 , n5510 );
nand ( n13987 , n7981 , n13986 );
buf ( n13988 , n5511 );
not ( n13989 , n13988 );
and ( n13990 , n13987 , n13989 );
not ( n13991 , n13987 );
buf ( n13992 , n13988 );
and ( n13993 , n13991 , n13992 );
nor ( n13994 , n13990 , n13993 );
xor ( n13995 , n13985 , n13994 );
buf ( n13996 , n5512 );
nand ( n13997 , n7515 , n13996 );
buf ( n13998 , n5513 );
not ( n13999 , n13998 );
and ( n14000 , n13997 , n13999 );
not ( n14001 , n13997 );
buf ( n14002 , n13998 );
and ( n14003 , n14001 , n14002 );
nor ( n14004 , n14000 , n14003 );
xnor ( n14005 , n13995 , n14004 );
not ( n14006 , n14005 );
not ( n14007 , n14006 );
not ( n14008 , n14007 );
and ( n14009 , n13967 , n14008 );
not ( n14010 , n13967 );
and ( n14011 , n14010 , n14007 );
nor ( n14012 , n14009 , n14011 );
not ( n14013 , n14012 );
not ( n14014 , n14013 );
and ( n14015 , n13959 , n14014 );
and ( n14016 , n13958 , n14013 );
nor ( n14017 , n14015 , n14016 );
xor ( n14018 , n10474 , n8072 );
not ( n14019 , n11298 );
buf ( n14020 , n5514 );
not ( n14021 , n14020 );
not ( n14022 , n14021 );
or ( n14023 , n14019 , n14022 );
not ( n14024 , n11297 );
buf ( n14025 , n14020 );
nand ( n14026 , n14024 , n14025 );
nand ( n14027 , n14023 , n14026 );
buf ( n14028 , n5515 );
not ( n14029 , n14028 );
and ( n14030 , n14027 , n14029 );
not ( n14031 , n14027 );
buf ( n14032 , n14028 );
and ( n14033 , n14031 , n14032 );
nor ( n14034 , n14030 , n14033 );
buf ( n14035 , n5516 );
nand ( n14036 , n7288 , n14035 );
buf ( n14037 , n5517 );
buf ( n14038 , n14037 );
and ( n14039 , n14036 , n14038 );
not ( n14040 , n14036 );
not ( n14041 , n14037 );
and ( n14042 , n14040 , n14041 );
nor ( n14043 , n14039 , n14042 );
xor ( n14044 , n14034 , n14043 );
buf ( n14045 , n5518 );
nand ( n14046 , n8520 , n14045 );
buf ( n14047 , n5519 );
not ( n14048 , n14047 );
and ( n14049 , n14046 , n14048 );
not ( n14050 , n14046 );
buf ( n14051 , n14047 );
and ( n14052 , n14050 , n14051 );
nor ( n14053 , n14049 , n14052 );
xnor ( n14054 , n14044 , n14053 );
not ( n14055 , n14054 );
buf ( n14056 , n14055 );
xnor ( n14057 , n14018 , n14056 );
not ( n14058 , n14057 );
xor ( n14059 , n8444 , n11768 );
xnor ( n14060 , n14059 , n11776 );
buf ( n14061 , n14060 );
not ( n14062 , n14061 );
not ( n14063 , n6696 );
buf ( n14064 , n5520 );
buf ( n14065 , n14064 );
not ( n14066 , n14065 );
buf ( n14067 , n5521 );
not ( n14068 , n14067 );
not ( n14069 , n14068 );
or ( n14070 , n14066 , n14069 );
not ( n14071 , n14064 );
buf ( n14072 , n14067 );
nand ( n14073 , n14071 , n14072 );
nand ( n14074 , n14070 , n14073 );
buf ( n14075 , n5522 );
not ( n14076 , n14075 );
and ( n14077 , n14074 , n14076 );
not ( n14078 , n14074 );
buf ( n14079 , n14075 );
and ( n14080 , n14078 , n14079 );
nor ( n14081 , n14077 , n14080 );
buf ( n14082 , n5523 );
nand ( n14083 , n7981 , n14082 );
buf ( n14084 , n5524 );
buf ( n14085 , n14084 );
and ( n14086 , n14083 , n14085 );
not ( n14087 , n14083 );
not ( n14088 , n14084 );
and ( n14089 , n14087 , n14088 );
nor ( n14090 , n14086 , n14089 );
xor ( n14091 , n14081 , n14090 );
buf ( n14092 , n5525 );
nand ( n14093 , n6706 , n14092 );
buf ( n14094 , n5526 );
not ( n14095 , n14094 );
and ( n14096 , n14093 , n14095 );
not ( n14097 , n14093 );
buf ( n14098 , n14094 );
and ( n14099 , n14097 , n14098 );
nor ( n14100 , n14096 , n14099 );
xnor ( n14101 , n14091 , n14100 );
not ( n14102 , n14101 );
or ( n14103 , n14063 , n14102 );
not ( n14104 , n14090 );
not ( n14105 , n14100 );
or ( n14106 , n14104 , n14105 );
or ( n14107 , n14090 , n14100 );
nand ( n14108 , n14106 , n14107 );
not ( n14109 , n14081 );
and ( n14110 , n14108 , n14109 );
not ( n14111 , n14108 );
and ( n14112 , n14111 , n14081 );
nor ( n14113 , n14110 , n14112 );
nand ( n14114 , n14113 , n6692 );
nand ( n14115 , n14103 , n14114 );
not ( n14116 , n14115 );
or ( n14117 , n14062 , n14116 );
not ( n14118 , n14115 );
nand ( n14119 , n14118 , n11778 );
nand ( n14120 , n14117 , n14119 );
not ( n14121 , n14120 );
nand ( n14122 , n14058 , n14121 );
buf ( n14123 , n5527 );
buf ( n14124 , n14123 );
not ( n14125 , n14124 );
buf ( n14126 , n5528 );
not ( n14127 , n14126 );
not ( n14128 , n14127 );
or ( n14129 , n14125 , n14128 );
not ( n14130 , n14123 );
buf ( n14131 , n14126 );
nand ( n14132 , n14130 , n14131 );
nand ( n14133 , n14129 , n14132 );
buf ( n14134 , n5529 );
not ( n14135 , n14134 );
and ( n14136 , n14133 , n14135 );
not ( n14137 , n14133 );
buf ( n14138 , n14134 );
and ( n14139 , n14137 , n14138 );
nor ( n14140 , n14136 , n14139 );
buf ( n14141 , n5530 );
nand ( n14142 , n6803 , n14141 );
buf ( n14143 , n5531 );
buf ( n14144 , n14143 );
and ( n14145 , n14142 , n14144 );
not ( n14146 , n14142 );
not ( n14147 , n14143 );
and ( n14148 , n14146 , n14147 );
nor ( n14149 , n14145 , n14148 );
xor ( n14150 , n14140 , n14149 );
buf ( n14151 , n5532 );
nand ( n14152 , n6816 , n14151 );
buf ( n14153 , n5533 );
not ( n14154 , n14153 );
and ( n14155 , n14152 , n14154 );
not ( n14156 , n14152 );
buf ( n14157 , n14153 );
and ( n14158 , n14156 , n14157 );
nor ( n14159 , n14155 , n14158 );
xnor ( n14160 , n14150 , n14159 );
not ( n14161 , n14160 );
buf ( n14162 , n5534 );
buf ( n14163 , n14162 );
not ( n14164 , n14163 );
and ( n14165 , n14161 , n14164 );
and ( n14166 , n14160 , n14163 );
nor ( n14167 , n14165 , n14166 );
buf ( n14168 , n5535 );
buf ( n14169 , n14168 );
not ( n14170 , n14169 );
buf ( n14171 , n5536 );
not ( n14172 , n14171 );
not ( n14173 , n14172 );
or ( n14174 , n14170 , n14173 );
not ( n14175 , n14168 );
buf ( n14176 , n14171 );
nand ( n14177 , n14175 , n14176 );
nand ( n14178 , n14174 , n14177 );
buf ( n14179 , n5537 );
buf ( n14180 , n14179 );
and ( n14181 , n14178 , n14180 );
not ( n14182 , n14178 );
not ( n14183 , n14179 );
and ( n14184 , n14182 , n14183 );
nor ( n14185 , n14181 , n14184 );
not ( n14186 , n14185 );
buf ( n14187 , n5538 );
nand ( n14188 , n7195 , n14187 );
buf ( n14189 , n5539 );
buf ( n14190 , n14189 );
and ( n14191 , n14188 , n14190 );
not ( n14192 , n14188 );
not ( n14193 , n14189 );
and ( n14194 , n14192 , n14193 );
nor ( n14195 , n14191 , n14194 );
xor ( n14196 , n14186 , n14195 );
buf ( n14197 , n5540 );
nand ( n14198 , n8971 , n14197 );
buf ( n14199 , n5541 );
not ( n14200 , n14199 );
and ( n14201 , n14198 , n14200 );
not ( n14202 , n14198 );
buf ( n14203 , n14199 );
and ( n14204 , n14202 , n14203 );
nor ( n14205 , n14201 , n14204 );
xnor ( n14206 , n14196 , n14205 );
not ( n14207 , n14206 );
not ( n14208 , n14207 );
and ( n14209 , n14167 , n14208 );
not ( n14210 , n14167 );
xor ( n14211 , n14185 , n14195 );
xnor ( n14212 , n14211 , n14205 );
buf ( n14213 , n14212 );
and ( n14214 , n14210 , n14213 );
nor ( n14215 , n14209 , n14214 );
not ( n14216 , n14215 );
and ( n14217 , n14122 , n14216 );
not ( n14218 , n14122 );
and ( n14219 , n14218 , n14215 );
nor ( n14220 , n14217 , n14219 );
xor ( n14221 , n14017 , n14220 );
buf ( n14222 , n5542 );
buf ( n14223 , n14222 );
not ( n14224 , n14223 );
buf ( n14225 , n5543 );
buf ( n14226 , n5544 );
not ( n14227 , n14226 );
buf ( n14228 , n5545 );
buf ( n14229 , n14228 );
nand ( n14230 , n14227 , n14229 );
not ( n14231 , n14228 );
buf ( n14232 , n14226 );
nand ( n14233 , n14231 , n14232 );
and ( n14234 , n14230 , n14233 );
xor ( n14235 , n14225 , n14234 );
buf ( n14236 , n5546 );
buf ( n14237 , n5547 );
xor ( n14238 , n14236 , n14237 );
buf ( n14239 , n5548 );
nand ( n14240 , n7184 , n14239 );
xnor ( n14241 , n14238 , n14240 );
xnor ( n14242 , n14235 , n14241 );
not ( n14243 , n14242 );
not ( n14244 , n14243 );
or ( n14245 , n14224 , n14244 );
not ( n14246 , n14242 );
or ( n14247 , n14246 , n14223 );
nand ( n14248 , n14245 , n14247 );
buf ( n14249 , n5549 );
not ( n14250 , n14249 );
buf ( n14251 , n5550 );
buf ( n14252 , n14251 );
not ( n14253 , n14252 );
buf ( n14254 , n5551 );
not ( n14255 , n14254 );
not ( n14256 , n14255 );
or ( n14257 , n14253 , n14256 );
not ( n14258 , n14251 );
buf ( n14259 , n14254 );
nand ( n14260 , n14258 , n14259 );
nand ( n14261 , n14257 , n14260 );
not ( n14262 , n14261 );
xor ( n14263 , n14250 , n14262 );
buf ( n14264 , n5552 );
nand ( n14265 , n7094 , n14264 );
buf ( n14266 , n5553 );
buf ( n14267 , n14266 );
and ( n14268 , n14265 , n14267 );
not ( n14269 , n14265 );
not ( n14270 , n14266 );
and ( n14271 , n14269 , n14270 );
nor ( n14272 , n14268 , n14271 );
not ( n14273 , n14272 );
buf ( n14274 , n5554 );
nand ( n14275 , n6608 , n14274 );
buf ( n14276 , n5555 );
buf ( n14277 , n14276 );
and ( n14278 , n14275 , n14277 );
not ( n14279 , n14275 );
not ( n14280 , n14276 );
and ( n14281 , n14279 , n14280 );
nor ( n14282 , n14278 , n14281 );
not ( n14283 , n14282 );
not ( n14284 , n14283 );
or ( n14285 , n14273 , n14284 );
not ( n14286 , n14272 );
nand ( n14287 , n14282 , n14286 );
nand ( n14288 , n14285 , n14287 );
xnor ( n14289 , n14263 , n14288 );
not ( n14290 , n14289 );
and ( n14291 , n14248 , n14290 );
not ( n14292 , n14248 );
buf ( n14293 , n14289 );
and ( n14294 , n14292 , n14293 );
nor ( n14295 , n14291 , n14294 );
not ( n14296 , n14295 );
not ( n14297 , n13640 );
buf ( n14298 , n5556 );
buf ( n14299 , n14298 );
not ( n14300 , n14299 );
buf ( n14301 , n5557 );
not ( n14302 , n14301 );
not ( n14303 , n14302 );
or ( n14304 , n14300 , n14303 );
not ( n14305 , n14298 );
buf ( n14306 , n14301 );
nand ( n14307 , n14305 , n14306 );
nand ( n14308 , n14304 , n14307 );
buf ( n14309 , n5558 );
buf ( n14310 , n14309 );
and ( n14311 , n14308 , n14310 );
not ( n14312 , n14308 );
not ( n14313 , n14309 );
and ( n14314 , n14312 , n14313 );
nor ( n14315 , n14311 , n14314 );
buf ( n14316 , n5559 );
nand ( n14317 , n6851 , n14316 );
buf ( n14318 , n5560 );
buf ( n14319 , n14318 );
and ( n14320 , n14317 , n14319 );
not ( n14321 , n14317 );
not ( n14322 , n14318 );
and ( n14323 , n14321 , n14322 );
nor ( n14324 , n14320 , n14323 );
not ( n14325 , n14324 );
xor ( n14326 , n14315 , n14325 );
buf ( n14327 , n5561 );
nand ( n14328 , n9159 , n14327 );
buf ( n14329 , n5562 );
not ( n14330 , n14329 );
and ( n14331 , n14328 , n14330 );
not ( n14332 , n14328 );
buf ( n14333 , n14329 );
and ( n14334 , n14332 , n14333 );
nor ( n14335 , n14331 , n14334 );
xnor ( n14336 , n14326 , n14335 );
buf ( n14337 , n14336 );
not ( n14338 , n14337 );
or ( n14339 , n14297 , n14338 );
xor ( n14340 , n14315 , n14324 );
xnor ( n14341 , n14340 , n14335 );
buf ( n14342 , n14341 );
buf ( n14343 , n14342 );
nand ( n14344 , n14343 , n13637 );
nand ( n14345 , n14339 , n14344 );
buf ( n14346 , n5563 );
buf ( n14347 , n14346 );
not ( n14348 , n14347 );
buf ( n14349 , n5564 );
not ( n14350 , n14349 );
not ( n14351 , n14350 );
or ( n14352 , n14348 , n14351 );
not ( n14353 , n14346 );
buf ( n14354 , n14349 );
nand ( n14355 , n14353 , n14354 );
nand ( n14356 , n14352 , n14355 );
buf ( n14357 , n5565 );
buf ( n14358 , n14357 );
and ( n14359 , n14356 , n14358 );
not ( n14360 , n14356 );
not ( n14361 , n14357 );
and ( n14362 , n14360 , n14361 );
nor ( n14363 , n14359 , n14362 );
buf ( n14364 , n5566 );
nand ( n14365 , n7133 , n14364 );
buf ( n14366 , n5567 );
buf ( n14367 , n14366 );
and ( n14368 , n14365 , n14367 );
not ( n14369 , n14365 );
not ( n14370 , n14366 );
and ( n14371 , n14369 , n14370 );
nor ( n14372 , n14368 , n14371 );
xor ( n14373 , n14363 , n14372 );
buf ( n14374 , n5568 );
nand ( n14375 , n8269 , n14374 );
buf ( n14376 , n5569 );
not ( n14377 , n14376 );
and ( n14378 , n14375 , n14377 );
not ( n14379 , n14375 );
buf ( n14380 , n14376 );
and ( n14381 , n14379 , n14380 );
nor ( n14382 , n14378 , n14381 );
xnor ( n14383 , n14373 , n14382 );
not ( n14384 , n14383 );
buf ( n14385 , n14384 );
not ( n14386 , n14385 );
and ( n14387 , n14345 , n14386 );
not ( n14388 , n14345 );
and ( n14389 , n14388 , n14385 );
nor ( n14390 , n14387 , n14389 );
nand ( n14391 , n14296 , n14390 );
buf ( n14392 , n5570 );
buf ( n14393 , n14392 );
not ( n14394 , n14393 );
buf ( n14395 , n5571 );
not ( n14396 , n14395 );
not ( n14397 , n14396 );
or ( n14398 , n14394 , n14397 );
not ( n14399 , n14392 );
buf ( n14400 , n14395 );
nand ( n14401 , n14399 , n14400 );
nand ( n14402 , n14398 , n14401 );
buf ( n14403 , n5572 );
buf ( n14404 , n14403 );
and ( n14405 , n14402 , n14404 );
not ( n14406 , n14402 );
not ( n14407 , n14403 );
and ( n14408 , n14406 , n14407 );
nor ( n14409 , n14405 , n14408 );
buf ( n14410 , n5573 );
nand ( n14411 , n7230 , n14410 );
buf ( n14412 , n5574 );
buf ( n14413 , n14412 );
and ( n14414 , n14411 , n14413 );
not ( n14415 , n14411 );
not ( n14416 , n14412 );
and ( n14417 , n14415 , n14416 );
nor ( n14418 , n14414 , n14417 );
xor ( n14419 , n14409 , n14418 );
buf ( n14420 , n5575 );
nand ( n14421 , n8934 , n14420 );
buf ( n14422 , n5576 );
buf ( n14423 , n14422 );
and ( n14424 , n14421 , n14423 );
not ( n14425 , n14421 );
not ( n14426 , n14422 );
and ( n14427 , n14425 , n14426 );
nor ( n14428 , n14424 , n14427 );
xnor ( n14429 , n14419 , n14428 );
buf ( n14430 , n14429 );
not ( n14431 , n14430 );
buf ( n14432 , n5577 );
not ( n14433 , n14432 );
not ( n14434 , n14433 );
buf ( n14435 , n5578 );
buf ( n14436 , n14435 );
not ( n14437 , n14436 );
buf ( n14438 , n5579 );
not ( n14439 , n14438 );
not ( n14440 , n14439 );
or ( n14441 , n14437 , n14440 );
not ( n14442 , n14435 );
buf ( n14443 , n14438 );
nand ( n14444 , n14442 , n14443 );
nand ( n14445 , n14441 , n14444 );
buf ( n14446 , n5580 );
buf ( n14447 , n14446 );
and ( n14448 , n14445 , n14447 );
not ( n14449 , n14445 );
not ( n14450 , n14446 );
and ( n14451 , n14449 , n14450 );
nor ( n14452 , n14448 , n14451 );
buf ( n14453 , n5581 );
nand ( n14454 , n8134 , n14453 );
buf ( n14455 , n5582 );
buf ( n14456 , n14455 );
and ( n14457 , n14454 , n14456 );
not ( n14458 , n14454 );
not ( n14459 , n14455 );
and ( n14460 , n14458 , n14459 );
nor ( n14461 , n14457 , n14460 );
xor ( n14462 , n14452 , n14461 );
xnor ( n14463 , n14462 , n10657 );
not ( n14464 , n14463 );
not ( n14465 , n14464 );
or ( n14466 , n14434 , n14465 );
or ( n14467 , n14464 , n14433 );
nand ( n14468 , n14466 , n14467 );
not ( n14469 , n14468 );
or ( n14470 , n14431 , n14469 );
not ( n14471 , n14429 );
not ( n14472 , n14471 );
or ( n14473 , n14468 , n14472 );
nand ( n14474 , n14470 , n14473 );
buf ( n14475 , n14474 );
not ( n14476 , n14475 );
and ( n14477 , n14391 , n14476 );
not ( n14478 , n14391 );
and ( n14479 , n14478 , n14475 );
nor ( n14480 , n14477 , n14479 );
xnor ( n14481 , n14221 , n14480 );
not ( n14482 , n14481 );
not ( n14483 , n14482 );
not ( n14484 , n11201 );
not ( n14485 , n10540 );
or ( n14486 , n14484 , n14485 );
nand ( n14487 , n10543 , n11197 );
nand ( n14488 , n14486 , n14487 );
not ( n14489 , n9394 );
xor ( n14490 , n14488 , n14489 );
not ( n14491 , n14490 );
not ( n14492 , n11691 );
buf ( n14493 , n10374 );
not ( n14494 , n14493 );
not ( n14495 , n14494 );
or ( n14496 , n14492 , n14495 );
nand ( n14497 , n14493 , n11694 );
nand ( n14498 , n14496 , n14497 );
not ( n14499 , n14498 );
buf ( n14500 , n5583 );
buf ( n14501 , n5584 );
buf ( n14502 , n14501 );
not ( n14503 , n14502 );
buf ( n14504 , n5585 );
not ( n14505 , n14504 );
not ( n14506 , n14505 );
or ( n14507 , n14503 , n14506 );
not ( n14508 , n14501 );
buf ( n14509 , n14504 );
nand ( n14510 , n14508 , n14509 );
nand ( n14511 , n14507 , n14510 );
xor ( n14512 , n14500 , n14511 );
buf ( n14513 , n5586 );
buf ( n14514 , n5587 );
not ( n14515 , n14514 );
xor ( n14516 , n14513 , n14515 );
buf ( n14517 , n5588 );
nand ( n14518 , n9159 , n14517 );
xnor ( n14519 , n14516 , n14518 );
xnor ( n14520 , n14512 , n14519 );
buf ( n14521 , n14520 );
not ( n14522 , n14521 );
not ( n14523 , n14522 );
and ( n14524 , n14499 , n14523 );
and ( n14525 , n14522 , n14498 );
nor ( n14526 , n14524 , n14525 );
not ( n14527 , n14526 );
nand ( n14528 , n14491 , n14527 );
not ( n14529 , n14528 );
buf ( n14530 , n5589 );
buf ( n14531 , n14530 );
not ( n14532 , n14531 );
buf ( n14533 , n8279 );
not ( n14534 , n14533 );
not ( n14535 , n14534 );
or ( n14536 , n14532 , n14535 );
buf ( n14537 , n8280 );
or ( n14538 , n14537 , n14531 );
nand ( n14539 , n14536 , n14538 );
not ( n14540 , n8238 );
and ( n14541 , n14539 , n14540 );
not ( n14542 , n14539 );
and ( n14543 , n14542 , n8238 );
nor ( n14544 , n14541 , n14543 );
not ( n14545 , n14544 );
and ( n14546 , n14529 , n14545 );
and ( n14547 , n14528 , n14544 );
nor ( n14548 , n14546 , n14547 );
buf ( n14549 , n8357 );
not ( n14550 , n14549 );
buf ( n14551 , n5590 );
nand ( n14552 , n8134 , n14551 );
buf ( n14553 , n5591 );
buf ( n14554 , n14553 );
and ( n14555 , n14552 , n14554 );
not ( n14556 , n14552 );
not ( n14557 , n14553 );
and ( n14558 , n14556 , n14557 );
nor ( n14559 , n14555 , n14558 );
not ( n14560 , n14559 );
buf ( n14561 , n5592 );
nand ( n14562 , n12401 , n14561 );
buf ( n14563 , n5593 );
not ( n14564 , n14563 );
and ( n14565 , n14562 , n14564 );
not ( n14566 , n14562 );
buf ( n14567 , n14563 );
and ( n14568 , n14566 , n14567 );
nor ( n14569 , n14565 , n14568 );
not ( n14570 , n14569 );
or ( n14571 , n14560 , n14570 );
or ( n14572 , n14559 , n14569 );
nand ( n14573 , n14571 , n14572 );
not ( n14574 , n12904 );
buf ( n14575 , n5594 );
not ( n14576 , n14575 );
not ( n14577 , n14576 );
or ( n14578 , n14574 , n14577 );
not ( n14579 , n12903 );
buf ( n14580 , n14575 );
nand ( n14581 , n14579 , n14580 );
nand ( n14582 , n14578 , n14581 );
buf ( n14583 , n5595 );
buf ( n14584 , n14583 );
and ( n14585 , n14582 , n14584 );
not ( n14586 , n14582 );
not ( n14587 , n14583 );
and ( n14588 , n14586 , n14587 );
nor ( n14589 , n14585 , n14588 );
not ( n14590 , n14589 );
xor ( n14591 , n14573 , n14590 );
buf ( n14592 , n14591 );
not ( n14593 , n14592 );
or ( n14594 , n14550 , n14593 );
xor ( n14595 , n14589 , n14559 );
xnor ( n14596 , n14595 , n14569 );
buf ( n14597 , n14596 );
nand ( n14598 , n14597 , n8358 );
nand ( n14599 , n14594 , n14598 );
buf ( n14600 , n9302 );
and ( n14601 , n14599 , n14600 );
not ( n14602 , n14599 );
buf ( n14603 , n9294 );
and ( n14604 , n14602 , n14603 );
nor ( n14605 , n14601 , n14604 );
not ( n14606 , n14605 );
buf ( n14607 , n5596 );
buf ( n14608 , n14607 );
buf ( n14609 , n5597 );
buf ( n14610 , n14609 );
not ( n14611 , n14610 );
buf ( n14612 , n5598 );
not ( n14613 , n14612 );
not ( n14614 , n14613 );
or ( n14615 , n14611 , n14614 );
not ( n14616 , n14609 );
buf ( n14617 , n14612 );
nand ( n14618 , n14616 , n14617 );
nand ( n14619 , n14615 , n14618 );
buf ( n14620 , n5599 );
not ( n14621 , n14620 );
and ( n14622 , n14619 , n14621 );
not ( n14623 , n14619 );
buf ( n14624 , n14620 );
and ( n14625 , n14623 , n14624 );
nor ( n14626 , n14622 , n14625 );
buf ( n14627 , n5600 );
nand ( n14628 , n7133 , n14627 );
buf ( n14629 , n5601 );
xor ( n14630 , n14628 , n14629 );
xor ( n14631 , n14626 , n14630 );
buf ( n14632 , n5602 );
nand ( n14633 , n6945 , n14632 );
buf ( n14634 , n5603 );
not ( n14635 , n14634 );
and ( n14636 , n14633 , n14635 );
not ( n14637 , n14633 );
buf ( n14638 , n14634 );
and ( n14639 , n14637 , n14638 );
nor ( n14640 , n14636 , n14639 );
xnor ( n14641 , n14631 , n14640 );
not ( n14642 , n14641 );
xor ( n14643 , n14608 , n14642 );
buf ( n14644 , n5604 );
buf ( n14645 , n5605 );
buf ( n14646 , n14645 );
not ( n14647 , n14646 );
buf ( n14648 , n5606 );
not ( n14649 , n14648 );
not ( n14650 , n14649 );
or ( n14651 , n14647 , n14650 );
not ( n14652 , n14645 );
buf ( n14653 , n14648 );
nand ( n14654 , n14652 , n14653 );
nand ( n14655 , n14651 , n14654 );
xor ( n14656 , n14644 , n14655 );
buf ( n14657 , n5607 );
buf ( n14658 , n5608 );
xor ( n14659 , n14657 , n14658 );
buf ( n14660 , n5609 );
nand ( n14661 , n9159 , n14660 );
xnor ( n14662 , n14659 , n14661 );
xnor ( n14663 , n14656 , n14662 );
buf ( n14664 , n14663 );
xnor ( n14665 , n14643 , n14664 );
nand ( n14666 , n14606 , n14665 );
not ( n14667 , n14666 );
not ( n14668 , n9244 );
buf ( n14669 , n5610 );
not ( n14670 , n14669 );
not ( n14671 , n14670 );
buf ( n14672 , n5611 );
buf ( n14673 , n14672 );
not ( n14674 , n14673 );
buf ( n14675 , n5612 );
not ( n14676 , n14675 );
not ( n14677 , n14676 );
or ( n14678 , n14674 , n14677 );
not ( n14679 , n14672 );
buf ( n14680 , n14675 );
nand ( n14681 , n14679 , n14680 );
nand ( n14682 , n14678 , n14681 );
buf ( n14683 , n5613 );
not ( n14684 , n14683 );
and ( n14685 , n14682 , n14684 );
not ( n14686 , n14682 );
buf ( n14687 , n14683 );
and ( n14688 , n14686 , n14687 );
nor ( n14689 , n14685 , n14688 );
buf ( n14690 , n5614 );
nand ( n14691 , n7616 , n14690 );
buf ( n14692 , n5615 );
not ( n14693 , n14692 );
and ( n14694 , n14691 , n14693 );
not ( n14695 , n14691 );
buf ( n14696 , n14692 );
and ( n14697 , n14695 , n14696 );
nor ( n14698 , n14694 , n14697 );
not ( n14699 , n14698 );
xor ( n14700 , n14689 , n14699 );
buf ( n14701 , n5616 );
nand ( n14702 , n7299 , n14701 );
buf ( n14703 , n5617 );
buf ( n14704 , n14703 );
and ( n14705 , n14702 , n14704 );
not ( n14706 , n14702 );
not ( n14707 , n14703 );
and ( n14708 , n14706 , n14707 );
nor ( n14709 , n14705 , n14708 );
buf ( n14710 , n14709 );
xnor ( n14711 , n14700 , n14710 );
not ( n14712 , n14711 );
or ( n14713 , n14671 , n14712 );
not ( n14714 , n14709 );
not ( n14715 , n14698 );
or ( n14716 , n14714 , n14715 );
or ( n14717 , n14709 , n14698 );
nand ( n14718 , n14716 , n14717 );
and ( n14719 , n14718 , n14689 );
not ( n14720 , n14718 );
not ( n14721 , n14689 );
and ( n14722 , n14720 , n14721 );
nor ( n14723 , n14719 , n14722 );
buf ( n14724 , n14669 );
nand ( n14725 , n14723 , n14724 );
nand ( n14726 , n14713 , n14725 );
not ( n14727 , n14726 );
or ( n14728 , n14668 , n14727 );
or ( n14729 , n14726 , n9244 );
nand ( n14730 , n14728 , n14729 );
not ( n14731 , n14730 );
and ( n14732 , n14667 , n14731 );
and ( n14733 , n14666 , n14730 );
nor ( n14734 , n14732 , n14733 );
not ( n14735 , n14734 );
and ( n14736 , n14548 , n14735 );
not ( n14737 , n14548 );
and ( n14738 , n14737 , n14734 );
nor ( n14739 , n14736 , n14738 );
not ( n14740 , n14739 );
not ( n14741 , n14740 );
and ( n14742 , n14483 , n14741 );
and ( n14743 , n14482 , n14740 );
nor ( n14744 , n14742 , n14743 );
not ( n14745 , n14744 );
or ( n14746 , n13957 , n14745 );
not ( n14747 , n13956 );
not ( n14748 , n14739 );
not ( n14749 , n14481 );
or ( n14750 , n14748 , n14749 );
not ( n14751 , n14481 );
nand ( n14752 , n14751 , n14740 );
nand ( n14753 , n14750 , n14752 );
nand ( n14754 , n14747 , n14753 );
nand ( n14755 , n14746 , n14754 );
not ( n14756 , n10808 );
buf ( n14757 , n14756 );
not ( n14758 , n14757 );
buf ( n14759 , n5618 );
buf ( n14760 , n14759 );
not ( n14761 , n14760 );
buf ( n14762 , n5619 );
buf ( n14763 , n14762 );
not ( n14764 , n14763 );
not ( n14765 , n13961 );
or ( n14766 , n14764 , n14765 );
not ( n14767 , n14762 );
buf ( n14768 , n13960 );
nand ( n14769 , n14767 , n14768 );
nand ( n14770 , n14766 , n14769 );
buf ( n14771 , n5620 );
not ( n14772 , n14771 );
and ( n14773 , n14770 , n14772 );
not ( n14774 , n14770 );
buf ( n14775 , n14771 );
and ( n14776 , n14774 , n14775 );
nor ( n14777 , n14773 , n14776 );
buf ( n14778 , n5621 );
nand ( n14779 , n6851 , n14778 );
buf ( n14780 , n5622 );
buf ( n14781 , n14780 );
and ( n14782 , n14779 , n14781 );
not ( n14783 , n14779 );
not ( n14784 , n14780 );
and ( n14785 , n14783 , n14784 );
nor ( n14786 , n14782 , n14785 );
xor ( n14787 , n14777 , n14786 );
buf ( n14788 , n5623 );
nand ( n14789 , n8785 , n14788 );
buf ( n14790 , n5624 );
not ( n14791 , n14790 );
and ( n14792 , n14789 , n14791 );
not ( n14793 , n14789 );
buf ( n14794 , n14790 );
and ( n14795 , n14793 , n14794 );
nor ( n14796 , n14792 , n14795 );
xnor ( n14797 , n14787 , n14796 );
not ( n14798 , n14797 );
or ( n14799 , n14761 , n14798 );
not ( n14800 , n14797 );
not ( n14801 , n14800 );
or ( n14802 , n14801 , n14760 );
nand ( n14803 , n14799 , n14802 );
not ( n14804 , n14803 );
or ( n14805 , n14758 , n14804 );
not ( n14806 , n10809 );
or ( n14807 , n14803 , n14806 );
nand ( n14808 , n14805 , n14807 );
not ( n14809 , n14808 );
buf ( n14810 , n12318 );
not ( n14811 , n14810 );
buf ( n14812 , n5625 );
nand ( n14813 , n6815 , n14812 );
buf ( n14814 , n5626 );
buf ( n14815 , n14814 );
and ( n14816 , n14813 , n14815 );
not ( n14817 , n14813 );
not ( n14818 , n14814 );
and ( n14819 , n14817 , n14818 );
nor ( n14820 , n14816 , n14819 );
buf ( n14821 , n14820 );
not ( n14822 , n14821 );
not ( n14823 , n14822 );
buf ( n14824 , n5627 );
buf ( n14825 , n14824 );
not ( n14826 , n14825 );
buf ( n14827 , n5628 );
not ( n14828 , n14827 );
not ( n14829 , n14828 );
or ( n14830 , n14826 , n14829 );
not ( n14831 , n14824 );
buf ( n14832 , n14827 );
nand ( n14833 , n14831 , n14832 );
nand ( n14834 , n14830 , n14833 );
buf ( n14835 , n5629 );
not ( n14836 , n14835 );
and ( n14837 , n14834 , n14836 );
not ( n14838 , n14834 );
buf ( n14839 , n14835 );
and ( n14840 , n14838 , n14839 );
nor ( n14841 , n14837 , n14840 );
buf ( n14842 , n5630 );
nand ( n14843 , n7299 , n14842 );
buf ( n14844 , n5631 );
buf ( n14845 , n14844 );
and ( n14846 , n14843 , n14845 );
not ( n14847 , n14843 );
not ( n14848 , n14844 );
and ( n14849 , n14847 , n14848 );
nor ( n14850 , n14846 , n14849 );
xor ( n14851 , n14841 , n14850 );
buf ( n14852 , n5632 );
nand ( n14853 , n8519 , n14852 );
buf ( n14854 , n5633 );
buf ( n14855 , n14854 );
and ( n14856 , n14853 , n14855 );
not ( n14857 , n14853 );
not ( n14858 , n14854 );
and ( n14859 , n14857 , n14858 );
nor ( n14860 , n14856 , n14859 );
not ( n14861 , n14860 );
xnor ( n14862 , n14851 , n14861 );
not ( n14863 , n14862 );
or ( n14864 , n14823 , n14863 );
xor ( n14865 , n14841 , n14860 );
buf ( n14866 , n14850 );
xnor ( n14867 , n14865 , n14866 );
nand ( n14868 , n14867 , n14821 );
nand ( n14869 , n14864 , n14868 );
not ( n14870 , n14869 );
or ( n14871 , n14811 , n14870 );
or ( n14872 , n14869 , n14810 );
nand ( n14873 , n14871 , n14872 );
not ( n14874 , n14873 );
not ( n14875 , n14521 );
buf ( n14876 , n11705 );
not ( n14877 , n14876 );
not ( n14878 , n10374 );
or ( n14879 , n14877 , n14878 );
or ( n14880 , n10374 , n14876 );
nand ( n14881 , n14879 , n14880 );
not ( n14882 , n14881 );
not ( n14883 , n14882 );
or ( n14884 , n14875 , n14883 );
nand ( n14885 , n14522 , n14881 );
nand ( n14886 , n14884 , n14885 );
nand ( n14887 , n14874 , n14886 );
not ( n14888 , n14887 );
or ( n14889 , n14809 , n14888 );
not ( n14890 , n14873 );
nand ( n14891 , n14890 , n14886 );
or ( n14892 , n14891 , n14808 );
nand ( n14893 , n14889 , n14892 );
not ( n14894 , n14893 );
not ( n14895 , n8612 );
buf ( n14896 , n5634 );
nand ( n14897 , n6945 , n14896 );
buf ( n14898 , n5635 );
not ( n14899 , n14898 );
and ( n14900 , n14897 , n14899 );
not ( n14901 , n14897 );
buf ( n14902 , n14898 );
and ( n14903 , n14901 , n14902 );
nor ( n14904 , n14900 , n14903 );
buf ( n14905 , n14904 );
and ( n14906 , n14905 , n8581 );
not ( n14907 , n14905 );
and ( n14908 , n14907 , n8580 );
nor ( n14909 , n14906 , n14908 );
not ( n14910 , n14909 );
and ( n14911 , n14895 , n14910 );
and ( n14912 , n8612 , n14909 );
nor ( n14913 , n14911 , n14912 );
not ( n14914 , n6772 );
buf ( n14915 , n5636 );
not ( n14916 , n14915 );
not ( n14917 , n6727 );
or ( n14918 , n14916 , n14917 );
xor ( n14919 , n6705 , n6725 );
not ( n14920 , n6715 );
xnor ( n14921 , n14919 , n14920 );
or ( n14922 , n14921 , n14915 );
nand ( n14923 , n14918 , n14922 );
not ( n14924 , n14923 );
or ( n14925 , n14914 , n14924 );
or ( n14926 , n14923 , n6773 );
nand ( n14927 , n14925 , n14926 );
nand ( n14928 , n14913 , n14927 );
not ( n14929 , n14928 );
buf ( n14930 , n5637 );
buf ( n14931 , n14930 );
not ( n14932 , n14931 );
buf ( n14933 , n5638 );
not ( n14934 , n14933 );
not ( n14935 , n14934 );
or ( n14936 , n14932 , n14935 );
not ( n14937 , n14930 );
buf ( n14938 , n14933 );
nand ( n14939 , n14937 , n14938 );
nand ( n14940 , n14936 , n14939 );
not ( n14941 , n14940 );
buf ( n14942 , n5639 );
not ( n14943 , n14942 );
buf ( n14944 , n5640 );
nand ( n14945 , n6660 , n14944 );
buf ( n14946 , n5641 );
buf ( n14947 , n14946 );
and ( n14948 , n14945 , n14947 );
not ( n14949 , n14945 );
not ( n14950 , n14946 );
and ( n14951 , n14949 , n14950 );
nor ( n14952 , n14948 , n14951 );
xor ( n14953 , n14943 , n14952 );
buf ( n14954 , n5642 );
nand ( n14955 , n8785 , n14954 );
buf ( n14956 , n5643 );
not ( n14957 , n14956 );
and ( n14958 , n14955 , n14957 );
not ( n14959 , n14955 );
buf ( n14960 , n14956 );
and ( n14961 , n14959 , n14960 );
nor ( n14962 , n14958 , n14961 );
xnor ( n14963 , n14953 , n14962 );
not ( n14964 , n14963 );
or ( n14965 , n14941 , n14964 );
not ( n14966 , n14963 );
not ( n14967 , n14940 );
nand ( n14968 , n14966 , n14967 );
nand ( n14969 , n14965 , n14968 );
not ( n14970 , n14969 );
not ( n14971 , n14970 );
not ( n14972 , n7465 );
buf ( n14973 , n5644 );
buf ( n14974 , n14973 );
not ( n14975 , n14974 );
buf ( n14976 , n5645 );
not ( n14977 , n14976 );
not ( n14978 , n14977 );
or ( n14979 , n14975 , n14978 );
not ( n14980 , n14973 );
buf ( n14981 , n14976 );
nand ( n14982 , n14980 , n14981 );
nand ( n14983 , n14979 , n14982 );
buf ( n14984 , n5646 );
not ( n14985 , n14984 );
and ( n14986 , n14983 , n14985 );
not ( n14987 , n14983 );
buf ( n14988 , n14984 );
and ( n14989 , n14987 , n14988 );
nor ( n14990 , n14986 , n14989 );
buf ( n14991 , n5647 );
nand ( n14992 , n6706 , n14991 );
buf ( n14993 , n5648 );
buf ( n14994 , n14993 );
and ( n14995 , n14992 , n14994 );
not ( n14996 , n14992 );
not ( n14997 , n14993 );
and ( n14998 , n14996 , n14997 );
nor ( n14999 , n14995 , n14998 );
xor ( n15000 , n14990 , n14999 );
buf ( n15001 , n5649 );
nand ( n15002 , n8785 , n15001 );
buf ( n15003 , n5650 );
buf ( n15004 , n15003 );
and ( n15005 , n15002 , n15004 );
not ( n15006 , n15002 );
not ( n15007 , n15003 );
and ( n15008 , n15006 , n15007 );
nor ( n15009 , n15005 , n15008 );
xnor ( n15010 , n15000 , n15009 );
not ( n15011 , n15010 );
not ( n15012 , n15011 );
or ( n15013 , n14972 , n15012 );
or ( n15014 , n15011 , n7465 );
nand ( n15015 , n15013 , n15014 );
not ( n15016 , n15015 );
and ( n15017 , n14971 , n15016 );
and ( n15018 , n14970 , n15015 );
nor ( n15019 , n15017 , n15018 );
not ( n15020 , n15019 );
not ( n15021 , n15020 );
and ( n15022 , n14929 , n15021 );
and ( n15023 , n14928 , n15020 );
nor ( n15024 , n15022 , n15023 );
not ( n15025 , n15024 );
or ( n15026 , n14894 , n15025 );
or ( n15027 , n15024 , n14893 );
nand ( n15028 , n15026 , n15027 );
not ( n15029 , n12353 );
not ( n15030 , n8976 );
or ( n15031 , n15029 , n15030 );
or ( n15032 , n8976 , n12353 );
nand ( n15033 , n15031 , n15032 );
and ( n15034 , n15033 , n13666 );
not ( n15035 , n15033 );
buf ( n15036 , n13663 );
and ( n15037 , n15035 , n15036 );
nor ( n15038 , n15034 , n15037 );
not ( n15039 , n15038 );
buf ( n15040 , n5651 );
nand ( n15041 , n7515 , n15040 );
buf ( n15042 , n5652 );
buf ( n15043 , n15042 );
and ( n15044 , n15041 , n15043 );
not ( n15045 , n15041 );
not ( n15046 , n15042 );
and ( n15047 , n15045 , n15046 );
nor ( n15048 , n15044 , n15047 );
buf ( n15049 , n15048 );
not ( n15050 , n15049 );
not ( n15051 , n13891 );
xor ( n15052 , n13882 , n15051 );
xnor ( n15053 , n15052 , n13901 );
not ( n15054 , n15053 );
or ( n15055 , n15050 , n15054 );
or ( n15056 , n15053 , n15049 );
nand ( n15057 , n15055 , n15056 );
and ( n15058 , n15057 , n13946 );
not ( n15059 , n15057 );
not ( n15060 , n13944 );
not ( n15061 , n15060 );
and ( n15062 , n15059 , n15061 );
nor ( n15063 , n15058 , n15062 );
not ( n15064 , n15063 );
nand ( n15065 , n15039 , n15064 );
buf ( n15066 , n11300 );
xor ( n15067 , n15066 , n7885 );
xor ( n15068 , n15067 , n7844 );
xor ( n15069 , n15065 , n15068 );
xor ( n15070 , n15028 , n15069 );
buf ( n15071 , n5653 );
nand ( n15072 , n7093 , n15071 );
buf ( n15073 , n5654 );
buf ( n15074 , n15073 );
and ( n15075 , n15072 , n15074 );
not ( n15076 , n15072 );
not ( n15077 , n15073 );
and ( n15078 , n15076 , n15077 );
nor ( n15079 , n15075 , n15078 );
not ( n15080 , n15079 );
buf ( n15081 , n5655 );
buf ( n15082 , n15081 );
not ( n15083 , n15082 );
buf ( n15084 , n5656 );
not ( n15085 , n15084 );
not ( n15086 , n15085 );
or ( n15087 , n15083 , n15086 );
not ( n15088 , n15081 );
buf ( n15089 , n15084 );
nand ( n15090 , n15088 , n15089 );
nand ( n15091 , n15087 , n15090 );
buf ( n15092 , n5657 );
buf ( n15093 , n15092 );
and ( n15094 , n15091 , n15093 );
not ( n15095 , n15091 );
not ( n15096 , n15092 );
and ( n15097 , n15095 , n15096 );
nor ( n15098 , n15094 , n15097 );
buf ( n15099 , n5658 );
nand ( n15100 , n6608 , n15099 );
buf ( n15101 , n5659 );
buf ( n15102 , n15101 );
and ( n15103 , n15100 , n15102 );
not ( n15104 , n15100 );
not ( n15105 , n15101 );
and ( n15106 , n15104 , n15105 );
nor ( n15107 , n15103 , n15106 );
xor ( n15108 , n15098 , n15107 );
buf ( n15109 , n5660 );
nand ( n15110 , n6804 , n15109 );
buf ( n15111 , n5661 );
buf ( n15112 , n15111 );
and ( n15113 , n15110 , n15112 );
not ( n15114 , n15110 );
not ( n15115 , n15111 );
and ( n15116 , n15114 , n15115 );
nor ( n15117 , n15113 , n15116 );
not ( n15118 , n15117 );
xnor ( n15119 , n15108 , n15118 );
buf ( n15120 , n15119 );
not ( n15121 , n15120 );
or ( n15122 , n15080 , n15121 );
or ( n15123 , n15120 , n15079 );
nand ( n15124 , n15122 , n15123 );
and ( n15125 , n15124 , n14597 );
not ( n15126 , n15124 );
buf ( n15127 , n14592 );
and ( n15128 , n15126 , n15127 );
nor ( n15129 , n15125 , n15128 );
not ( n15130 , n15129 );
not ( n15131 , n13651 );
not ( n15132 , n15131 );
not ( n15133 , n14337 );
or ( n15134 , n15132 , n15133 );
not ( n15135 , n15131 );
nand ( n15136 , n15135 , n14342 );
nand ( n15137 , n15134 , n15136 );
and ( n15138 , n15137 , n14386 );
not ( n15139 , n15137 );
and ( n15140 , n15139 , n14385 );
nor ( n15141 , n15138 , n15140 );
nor ( n15142 , n15130 , n15141 );
buf ( n15143 , n5662 );
buf ( n15144 , n15143 );
buf ( n15145 , n5663 );
buf ( n15146 , n15145 );
not ( n15147 , n15146 );
buf ( n15148 , n5664 );
not ( n15149 , n15148 );
not ( n15150 , n15149 );
or ( n15151 , n15147 , n15150 );
not ( n15152 , n15145 );
buf ( n15153 , n15148 );
nand ( n15154 , n15152 , n15153 );
nand ( n15155 , n15151 , n15154 );
buf ( n15156 , n5665 );
not ( n15157 , n15156 );
and ( n15158 , n15155 , n15157 );
not ( n15159 , n15155 );
buf ( n15160 , n15156 );
and ( n15161 , n15159 , n15160 );
nor ( n15162 , n15158 , n15161 );
buf ( n15163 , n5666 );
nand ( n15164 , n7094 , n15163 );
buf ( n15165 , n5667 );
buf ( n15166 , n15165 );
and ( n15167 , n15164 , n15166 );
not ( n15168 , n15164 );
not ( n15169 , n15165 );
and ( n15170 , n15168 , n15169 );
nor ( n15171 , n15167 , n15170 );
xor ( n15172 , n15162 , n15171 );
buf ( n15173 , n5668 );
nand ( n15174 , n6608 , n15173 );
buf ( n15175 , n5669 );
buf ( n15176 , n15175 );
and ( n15177 , n15174 , n15176 );
not ( n15178 , n15174 );
not ( n15179 , n15175 );
and ( n15180 , n15178 , n15179 );
nor ( n15181 , n15177 , n15180 );
not ( n15182 , n15181 );
xnor ( n15183 , n15172 , n15182 );
not ( n15184 , n15183 );
xor ( n15185 , n15144 , n15184 );
buf ( n15186 , n5670 );
not ( n15187 , n15186 );
buf ( n15188 , n5671 );
not ( n15189 , n15188 );
buf ( n15190 , n5672 );
buf ( n15191 , n15190 );
and ( n15192 , n15189 , n15191 );
not ( n15193 , n15189 );
not ( n15194 , n15190 );
and ( n15195 , n15193 , n15194 );
nor ( n15196 , n15192 , n15195 );
xor ( n15197 , n15187 , n15196 );
buf ( n15198 , n5673 );
buf ( n15199 , n5674 );
xor ( n15200 , n15198 , n15199 );
buf ( n15201 , n5675 );
nand ( n15202 , n7184 , n15201 );
xnor ( n15203 , n15200 , n15202 );
xnor ( n15204 , n15197 , n15203 );
not ( n15205 , n15204 );
not ( n15206 , n15205 );
xor ( n15207 , n15185 , n15206 );
and ( n15208 , n15142 , n15207 );
not ( n15209 , n15142 );
not ( n15210 , n15207 );
and ( n15211 , n15209 , n15210 );
nor ( n15212 , n15208 , n15211 );
not ( n15213 , n15212 );
not ( n15214 , n15213 );
buf ( n15215 , n5676 );
not ( n15216 , n15215 );
buf ( n15217 , n5677 );
nand ( n15218 , n6933 , n15217 );
buf ( n15219 , n5678 );
buf ( n15220 , n15219 );
and ( n15221 , n15218 , n15220 );
not ( n15222 , n15218 );
not ( n15223 , n15219 );
and ( n15224 , n15222 , n15223 );
nor ( n15225 , n15221 , n15224 );
xor ( n15226 , n15216 , n15225 );
buf ( n15227 , n5679 );
nand ( n15228 , n7288 , n15227 );
buf ( n15229 , n5680 );
buf ( n15230 , n15229 );
and ( n15231 , n15228 , n15230 );
not ( n15232 , n15228 );
not ( n15233 , n15229 );
and ( n15234 , n15232 , n15233 );
nor ( n15235 , n15231 , n15234 );
xnor ( n15236 , n15226 , n15235 );
not ( n15237 , n15236 );
buf ( n15238 , n5681 );
buf ( n15239 , n15238 );
not ( n15240 , n15239 );
buf ( n15241 , n5682 );
not ( n15242 , n15241 );
not ( n15243 , n15242 );
or ( n15244 , n15240 , n15243 );
not ( n15245 , n15238 );
buf ( n15246 , n15241 );
nand ( n15247 , n15245 , n15246 );
nand ( n15248 , n15244 , n15247 );
not ( n15249 , n15248 );
not ( n15250 , n15249 );
and ( n15251 , n15237 , n15250 );
and ( n15252 , n15236 , n15249 );
nor ( n15253 , n15251 , n15252 );
buf ( n15254 , n15253 );
not ( n15255 , n15254 );
not ( n15256 , n8790 );
buf ( n15257 , n5683 );
nand ( n15258 , n7230 , n15257 );
buf ( n15259 , n5684 );
buf ( n15260 , n15259 );
and ( n15261 , n15258 , n15260 );
not ( n15262 , n15258 );
not ( n15263 , n15259 );
and ( n15264 , n15262 , n15263 );
nor ( n15265 , n15261 , n15264 );
buf ( n15266 , n15265 );
nor ( n15267 , n15256 , n15266 );
not ( n15268 , n15267 );
nand ( n15269 , n15266 , n8791 );
nand ( n15270 , n15268 , n15269 );
not ( n15271 , n15270 );
or ( n15272 , n15255 , n15271 );
buf ( n15273 , n15253 );
or ( n15274 , n15270 , n15273 );
nand ( n15275 , n15272 , n15274 );
buf ( n15276 , n13151 );
and ( n15277 , n13155 , n15276 );
not ( n15278 , n13155 );
and ( n15279 , n15278 , n13152 );
nor ( n15280 , n15277 , n15279 );
not ( n15281 , n15280 );
not ( n15282 , n10895 );
not ( n15283 , n15282 );
or ( n15284 , n15281 , n15283 );
not ( n15285 , n10894 );
buf ( n15286 , n15285 );
not ( n15287 , n15286 );
or ( n15288 , n15287 , n15280 );
nand ( n15289 , n15284 , n15288 );
buf ( n15290 , n5685 );
buf ( n15291 , n15290 );
not ( n15292 , n15291 );
buf ( n15293 , n5686 );
not ( n15294 , n15293 );
not ( n15295 , n15294 );
or ( n15296 , n15292 , n15295 );
not ( n15297 , n15290 );
buf ( n15298 , n15293 );
nand ( n15299 , n15297 , n15298 );
nand ( n15300 , n15296 , n15299 );
buf ( n15301 , n5687 );
not ( n15302 , n15301 );
and ( n15303 , n15300 , n15302 );
not ( n15304 , n15300 );
buf ( n15305 , n15301 );
and ( n15306 , n15304 , n15305 );
nor ( n15307 , n15303 , n15306 );
buf ( n15308 , n5688 );
nand ( n15309 , n7288 , n15308 );
buf ( n15310 , n5689 );
not ( n15311 , n15310 );
and ( n15312 , n15309 , n15311 );
not ( n15313 , n15309 );
buf ( n15314 , n15310 );
and ( n15315 , n15313 , n15314 );
nor ( n15316 , n15312 , n15315 );
xor ( n15317 , n15307 , n15316 );
buf ( n15318 , n5690 );
nand ( n15319 , n7750 , n15318 );
buf ( n15320 , n5691 );
not ( n15321 , n15320 );
and ( n15322 , n15319 , n15321 );
not ( n15323 , n15319 );
buf ( n15324 , n15320 );
and ( n15325 , n15323 , n15324 );
nor ( n15326 , n15322 , n15325 );
xnor ( n15327 , n15317 , n15326 );
not ( n15328 , n15327 );
not ( n15329 , n15328 );
and ( n15330 , n15289 , n15329 );
not ( n15331 , n15289 );
buf ( n15332 , n15327 );
not ( n15333 , n15332 );
not ( n15334 , n15333 );
not ( n15335 , n15334 );
and ( n15336 , n15331 , n15335 );
nor ( n15337 , n15330 , n15336 );
not ( n15338 , n15337 );
nand ( n15339 , n15275 , n15338 );
not ( n15340 , n12442 );
buf ( n15341 , n5692 );
buf ( n15342 , n15341 );
not ( n15343 , n15342 );
buf ( n15344 , n5693 );
not ( n15345 , n15344 );
not ( n15346 , n15345 );
or ( n15347 , n15343 , n15346 );
not ( n15348 , n15341 );
buf ( n15349 , n15344 );
nand ( n15350 , n15348 , n15349 );
nand ( n15351 , n15347 , n15350 );
buf ( n15352 , n5694 );
not ( n15353 , n15352 );
and ( n15354 , n15351 , n15353 );
not ( n15355 , n15351 );
buf ( n15356 , n15352 );
and ( n15357 , n15355 , n15356 );
nor ( n15358 , n15354 , n15357 );
buf ( n15359 , n5695 );
nand ( n15360 , n7909 , n15359 );
buf ( n15361 , n5696 );
not ( n15362 , n15361 );
and ( n15363 , n15360 , n15362 );
not ( n15364 , n15360 );
buf ( n15365 , n15361 );
and ( n15366 , n15364 , n15365 );
nor ( n15367 , n15363 , n15366 );
xor ( n15368 , n15358 , n15367 );
xnor ( n15369 , n15368 , n13417 );
buf ( n15370 , n15369 );
not ( n15371 , n15370 );
not ( n15372 , n15371 );
or ( n15373 , n15340 , n15372 );
nand ( n15374 , n15370 , n12439 );
nand ( n15375 , n15373 , n15374 );
not ( n15376 , n15375 );
buf ( n15377 , n5697 );
buf ( n15378 , n5698 );
not ( n15379 , n15378 );
buf ( n15380 , n5699 );
buf ( n15381 , n15380 );
nand ( n15382 , n15379 , n15381 );
not ( n15383 , n15380 );
buf ( n15384 , n15378 );
nand ( n15385 , n15383 , n15384 );
and ( n15386 , n15382 , n15385 );
xor ( n15387 , n15377 , n15386 );
buf ( n15388 , n5700 );
buf ( n15389 , n5701 );
xor ( n15390 , n15388 , n15389 );
buf ( n15391 , n5702 );
nand ( n15392 , n6945 , n15391 );
xnor ( n15393 , n15390 , n15392 );
xnor ( n15394 , n15387 , n15393 );
buf ( n15395 , n15394 );
not ( n15396 , n15395 );
not ( n15397 , n15396 );
and ( n15398 , n15376 , n15397 );
and ( n15399 , n15375 , n15396 );
nor ( n15400 , n15398 , n15399 );
and ( n15401 , n15339 , n15400 );
not ( n15402 , n15339 );
not ( n15403 , n15400 );
and ( n15404 , n15402 , n15403 );
nor ( n15405 , n15401 , n15404 );
not ( n15406 , n15405 );
not ( n15407 , n15406 );
or ( n15408 , n15214 , n15407 );
nand ( n15409 , n15405 , n15212 );
nand ( n15410 , n15408 , n15409 );
not ( n15411 , n15410 );
and ( n15412 , n15070 , n15411 );
not ( n15413 , n15070 );
and ( n15414 , n15413 , n15410 );
nor ( n15415 , n15412 , n15414 );
buf ( n15416 , n15415 );
and ( n15417 , n14755 , n15416 );
not ( n15418 , n14755 );
and ( n15419 , n15070 , n15410 );
not ( n15420 , n15070 );
and ( n15421 , n15420 , n15411 );
nor ( n15422 , n15419 , n15421 );
buf ( n15423 , n15422 );
and ( n15424 , n15418 , n15423 );
nor ( n15425 , n15417 , n15424 );
not ( n15426 , n15425 );
not ( n15427 , n9430 );
nand ( n15428 , n15426 , n15427 );
not ( n15429 , n11753 );
and ( n15430 , n15428 , n15429 );
not ( n15431 , n15428 );
and ( n15432 , n15431 , n11753 );
nor ( n15433 , n15430 , n15432 );
not ( n15434 , n13746 );
buf ( n15435 , n15434 );
or ( n15436 , n15433 , n15435 );
nand ( n15437 , n13769 , n15436 );
buf ( n15438 , n15437 );
buf ( n15439 , n15438 );
not ( n15440 , n9243 );
buf ( n15441 , n5703 );
buf ( n15442 , n15441 );
not ( n15443 , n15442 );
not ( n15444 , n14723 );
or ( n15445 , n15443 , n15444 );
not ( n15446 , n15442 );
nand ( n15447 , n15446 , n14711 );
nand ( n15448 , n15445 , n15447 );
xor ( n15449 , n15440 , n15448 );
buf ( n15450 , n5704 );
buf ( n15451 , n15450 );
not ( n15452 , n15451 );
not ( n15453 , n12743 );
or ( n15454 , n15452 , n15453 );
or ( n15455 , n12743 , n15451 );
nand ( n15456 , n15454 , n15455 );
not ( n15457 , n15456 );
not ( n15458 , n12748 );
not ( n15459 , n15458 );
not ( n15460 , n15459 );
and ( n15461 , n15457 , n15460 );
and ( n15462 , n15456 , n12749 );
nor ( n15463 , n15461 , n15462 );
nand ( n15464 , n15449 , n15463 );
not ( n15465 , n9947 );
not ( n15466 , n7269 );
buf ( n15467 , n5705 );
not ( n15468 , n15467 );
not ( n15469 , n15468 );
or ( n15470 , n15466 , n15469 );
not ( n15471 , n7268 );
buf ( n15472 , n15467 );
nand ( n15473 , n15471 , n15472 );
nand ( n15474 , n15470 , n15473 );
buf ( n15475 , n5706 );
buf ( n15476 , n15475 );
and ( n15477 , n15474 , n15476 );
not ( n15478 , n15474 );
not ( n15479 , n15475 );
and ( n15480 , n15478 , n15479 );
nor ( n15481 , n15477 , n15480 );
buf ( n15482 , n5707 );
nand ( n15483 , n6816 , n15482 );
buf ( n15484 , n5708 );
buf ( n15485 , n15484 );
and ( n15486 , n15483 , n15485 );
not ( n15487 , n15483 );
not ( n15488 , n15484 );
and ( n15489 , n15487 , n15488 );
nor ( n15490 , n15486 , n15489 );
xor ( n15491 , n15481 , n15490 );
buf ( n15492 , n5709 );
nand ( n15493 , n8971 , n15492 );
buf ( n15494 , n5710 );
not ( n15495 , n15494 );
and ( n15496 , n15493 , n15495 );
not ( n15497 , n15493 );
buf ( n15498 , n15494 );
and ( n15499 , n15497 , n15498 );
nor ( n15500 , n15496 , n15499 );
xnor ( n15501 , n15491 , n15500 );
buf ( n15502 , n15501 );
not ( n15503 , n15502 );
not ( n15504 , n15503 );
or ( n15505 , n15465 , n15504 );
not ( n15506 , n9947 );
not ( n15507 , n15501 );
not ( n15508 , n15507 );
nand ( n15509 , n15506 , n15508 );
nand ( n15510 , n15505 , n15509 );
buf ( n15511 , n5711 );
buf ( n15512 , n15511 );
not ( n15513 , n15512 );
buf ( n15514 , n5712 );
not ( n15515 , n15514 );
not ( n15516 , n15515 );
or ( n15517 , n15513 , n15516 );
not ( n15518 , n15511 );
buf ( n15519 , n15514 );
nand ( n15520 , n15518 , n15519 );
nand ( n15521 , n15517 , n15520 );
buf ( n15522 , n5713 );
buf ( n15523 , n15522 );
and ( n15524 , n15521 , n15523 );
not ( n15525 , n15521 );
not ( n15526 , n15522 );
and ( n15527 , n15525 , n15526 );
nor ( n15528 , n15524 , n15527 );
buf ( n15529 , n5714 );
nand ( n15530 , n6803 , n15529 );
buf ( n15531 , n5715 );
buf ( n15532 , n15531 );
and ( n15533 , n15530 , n15532 );
not ( n15534 , n15530 );
not ( n15535 , n15531 );
and ( n15536 , n15534 , n15535 );
nor ( n15537 , n15533 , n15536 );
xor ( n15538 , n15528 , n15537 );
buf ( n15539 , n5716 );
nand ( n15540 , n7921 , n15539 );
buf ( n15541 , n5717 );
not ( n15542 , n15541 );
and ( n15543 , n15540 , n15542 );
not ( n15544 , n15540 );
buf ( n15545 , n15541 );
and ( n15546 , n15544 , n15545 );
nor ( n15547 , n15543 , n15546 );
xnor ( n15548 , n15538 , n15547 );
buf ( n15549 , n15548 );
not ( n15550 , n15549 );
and ( n15551 , n15510 , n15550 );
not ( n15552 , n15510 );
and ( n15553 , n15552 , n15549 );
nor ( n15554 , n15551 , n15553 );
xor ( n15555 , n15464 , n15554 );
not ( n15556 , n15555 );
buf ( n15557 , n9596 );
not ( n15558 , n15557 );
xor ( n15559 , n13642 , n13661 );
xnor ( n15560 , n15559 , n15131 );
not ( n15561 , n15560 );
not ( n15562 , n15561 );
or ( n15563 , n15558 , n15562 );
or ( n15564 , n13666 , n15557 );
nand ( n15565 , n15563 , n15564 );
and ( n15566 , n15565 , n13709 );
not ( n15567 , n15565 );
not ( n15568 , n13708 );
and ( n15569 , n15567 , n15568 );
nor ( n15570 , n15566 , n15569 );
not ( n15571 , n15570 );
not ( n15572 , n15571 );
buf ( n15573 , n5718 );
buf ( n15574 , n15573 );
not ( n15575 , n15574 );
buf ( n15576 , n5719 );
not ( n15577 , n15576 );
not ( n15578 , n15577 );
or ( n15579 , n15575 , n15578 );
not ( n15580 , n15573 );
buf ( n15581 , n15576 );
nand ( n15582 , n15580 , n15581 );
nand ( n15583 , n15579 , n15582 );
not ( n15584 , n15583 );
not ( n15585 , n15584 );
buf ( n15586 , n5720 );
buf ( n15587 , n5721 );
not ( n15588 , n15587 );
xor ( n15589 , n15586 , n15588 );
buf ( n15590 , n5722 );
not ( n15591 , n15590 );
buf ( n15592 , n5723 );
nand ( n15593 , n6851 , n15592 );
not ( n15594 , n15593 );
or ( n15595 , n15591 , n15594 );
nand ( n15596 , n7230 , n15592 );
or ( n15597 , n15596 , n15590 );
nand ( n15598 , n15595 , n15597 );
xnor ( n15599 , n15589 , n15598 );
not ( n15600 , n15599 );
or ( n15601 , n15585 , n15600 );
or ( n15602 , n15599 , n15584 );
nand ( n15603 , n15601 , n15602 );
buf ( n15604 , n15603 );
not ( n15605 , n15604 );
buf ( n15606 , n5724 );
nand ( n15607 , n7412 , n15606 );
buf ( n15608 , n5725 );
buf ( n15609 , n15608 );
and ( n15610 , n15607 , n15609 );
not ( n15611 , n15607 );
not ( n15612 , n15608 );
and ( n15613 , n15611 , n15612 );
nor ( n15614 , n15610 , n15613 );
not ( n15615 , n15614 );
buf ( n15616 , n5726 );
nand ( n15617 , n10107 , n15616 );
buf ( n15618 , n5727 );
not ( n15619 , n15618 );
and ( n15620 , n15617 , n15619 );
not ( n15621 , n15617 );
buf ( n15622 , n15618 );
and ( n15623 , n15621 , n15622 );
nor ( n15624 , n15620 , n15623 );
not ( n15625 , n15624 );
or ( n15626 , n15615 , n15625 );
or ( n15627 , n15614 , n15624 );
nand ( n15628 , n15626 , n15627 );
buf ( n15629 , n5728 );
buf ( n15630 , n15629 );
not ( n15631 , n15630 );
buf ( n15632 , n5729 );
not ( n15633 , n15632 );
not ( n15634 , n15633 );
or ( n15635 , n15631 , n15634 );
not ( n15636 , n15629 );
buf ( n15637 , n15632 );
nand ( n15638 , n15636 , n15637 );
nand ( n15639 , n15635 , n15638 );
buf ( n15640 , n5730 );
not ( n15641 , n15640 );
and ( n15642 , n15639 , n15641 );
not ( n15643 , n15639 );
buf ( n15644 , n15640 );
and ( n15645 , n15643 , n15644 );
nor ( n15646 , n15642 , n15645 );
xnor ( n15647 , n15628 , n15646 );
not ( n15648 , n15647 );
buf ( n15649 , n13377 );
not ( n15650 , n15649 );
and ( n15651 , n15648 , n15650 );
and ( n15652 , n15647 , n15649 );
nor ( n15653 , n15651 , n15652 );
not ( n15654 , n15653 );
and ( n15655 , n15605 , n15654 );
and ( n15656 , n15604 , n15653 );
nor ( n15657 , n15655 , n15656 );
buf ( n15658 , n5731 );
buf ( n15659 , n15658 );
not ( n15660 , n15659 );
buf ( n15661 , n5732 );
not ( n15662 , n15661 );
not ( n15663 , n15662 );
or ( n15664 , n15660 , n15663 );
not ( n15665 , n15658 );
buf ( n15666 , n15661 );
nand ( n15667 , n15665 , n15666 );
nand ( n15668 , n15664 , n15667 );
buf ( n15669 , n5733 );
buf ( n15670 , n15669 );
and ( n15671 , n15668 , n15670 );
not ( n15672 , n15668 );
not ( n15673 , n15669 );
and ( n15674 , n15672 , n15673 );
nor ( n15675 , n15671 , n15674 );
buf ( n15676 , n5734 );
nand ( n15677 , n10204 , n15676 );
buf ( n15678 , n5735 );
not ( n15679 , n15678 );
and ( n15680 , n15677 , n15679 );
not ( n15681 , n15677 );
buf ( n15682 , n15678 );
and ( n15683 , n15681 , n15682 );
nor ( n15684 , n15680 , n15683 );
xor ( n15685 , n15675 , n15684 );
buf ( n15686 , n5736 );
nand ( n15687 , n6906 , n15686 );
buf ( n15688 , n5737 );
not ( n15689 , n15688 );
and ( n15690 , n15687 , n15689 );
not ( n15691 , n15687 );
buf ( n15692 , n15688 );
and ( n15693 , n15691 , n15692 );
nor ( n15694 , n15690 , n15693 );
xnor ( n15695 , n15685 , n15694 );
not ( n15696 , n15695 );
not ( n15697 , n15696 );
not ( n15698 , n15697 );
not ( n15699 , n15698 );
buf ( n15700 , n5738 );
buf ( n15701 , n15700 );
not ( n15702 , n15701 );
buf ( n15703 , n5739 );
not ( n15704 , n15703 );
not ( n15705 , n15704 );
or ( n15706 , n15702 , n15705 );
not ( n15707 , n15700 );
buf ( n15708 , n15703 );
nand ( n15709 , n15707 , n15708 );
nand ( n15710 , n15706 , n15709 );
buf ( n15711 , n5740 );
buf ( n15712 , n15711 );
and ( n15713 , n15710 , n15712 );
not ( n15714 , n15710 );
not ( n15715 , n15711 );
and ( n15716 , n15714 , n15715 );
nor ( n15717 , n15713 , n15716 );
buf ( n15718 , n5741 );
nand ( n15719 , n7865 , n15718 );
buf ( n15720 , n5742 );
not ( n15721 , n15720 );
and ( n15722 , n15719 , n15721 );
not ( n15723 , n15719 );
buf ( n15724 , n15720 );
and ( n15725 , n15723 , n15724 );
nor ( n15726 , n15722 , n15725 );
xor ( n15727 , n15717 , n15726 );
buf ( n15728 , n5743 );
nand ( n15729 , n9159 , n15728 );
buf ( n15730 , n5744 );
not ( n15731 , n15730 );
and ( n15732 , n15729 , n15731 );
not ( n15733 , n15729 );
buf ( n15734 , n15730 );
and ( n15735 , n15733 , n15734 );
nor ( n15736 , n15732 , n15735 );
xnor ( n15737 , n15727 , n15736 );
not ( n15738 , n15737 );
not ( n15739 , n15738 );
not ( n15740 , n15739 );
not ( n15741 , n7742 );
and ( n15742 , n15740 , n15741 );
buf ( n15743 , n15737 );
and ( n15744 , n15743 , n7742 );
nor ( n15745 , n15742 , n15744 );
not ( n15746 , n15745 );
or ( n15747 , n15699 , n15746 );
buf ( n15748 , n15695 );
buf ( n15749 , n15748 );
not ( n15750 , n15749 );
or ( n15751 , n15745 , n15750 );
nand ( n15752 , n15747 , n15751 );
nand ( n15753 , n15657 , n15752 );
not ( n15754 , n15753 );
or ( n15755 , n15572 , n15754 );
or ( n15756 , n15753 , n15571 );
nand ( n15757 , n15755 , n15756 );
not ( n15758 , n15757 );
buf ( n15759 , n5745 );
buf ( n15760 , n15759 );
not ( n15761 , n15760 );
buf ( n15762 , n5746 );
not ( n15763 , n15762 );
not ( n15764 , n15763 );
or ( n15765 , n15761 , n15764 );
not ( n15766 , n15759 );
buf ( n15767 , n15762 );
nand ( n15768 , n15766 , n15767 );
nand ( n15769 , n15765 , n15768 );
not ( n15770 , n15769 );
buf ( n15771 , n5747 );
not ( n15772 , n15771 );
buf ( n15773 , n5748 );
nand ( n15774 , n7865 , n15773 );
buf ( n15775 , n5749 );
buf ( n15776 , n15775 );
and ( n15777 , n15774 , n15776 );
not ( n15778 , n15774 );
not ( n15779 , n15775 );
and ( n15780 , n15778 , n15779 );
nor ( n15781 , n15777 , n15780 );
xor ( n15782 , n15772 , n15781 );
buf ( n15783 , n5750 );
nand ( n15784 , n6863 , n15783 );
buf ( n15785 , n5751 );
buf ( n15786 , n15785 );
and ( n15787 , n15784 , n15786 );
not ( n15788 , n15784 );
not ( n15789 , n15785 );
and ( n15790 , n15788 , n15789 );
nor ( n15791 , n15787 , n15790 );
xnor ( n15792 , n15782 , n15791 );
xor ( n15793 , n15770 , n15792 );
not ( n15794 , n15793 );
buf ( n15795 , n9331 );
not ( n15796 , n15795 );
not ( n15797 , n14531 );
buf ( n15798 , n5752 );
not ( n15799 , n15798 );
not ( n15800 , n15799 );
or ( n15801 , n15797 , n15800 );
not ( n15802 , n14530 );
buf ( n15803 , n15798 );
nand ( n15804 , n15802 , n15803 );
nand ( n15805 , n15801 , n15804 );
not ( n15806 , n8240 );
and ( n15807 , n15805 , n15806 );
not ( n15808 , n15805 );
and ( n15809 , n15808 , n8241 );
nor ( n15810 , n15807 , n15809 );
buf ( n15811 , n5753 );
nand ( n15812 , n6660 , n15811 );
buf ( n15813 , n5754 );
buf ( n15814 , n15813 );
and ( n15815 , n15812 , n15814 );
not ( n15816 , n15812 );
not ( n15817 , n15813 );
and ( n15818 , n15816 , n15817 );
nor ( n15819 , n15815 , n15818 );
xor ( n15820 , n15810 , n15819 );
buf ( n15821 , n5755 );
nand ( n15822 , n7477 , n15821 );
buf ( n15823 , n5756 );
buf ( n15824 , n15823 );
and ( n15825 , n15822 , n15824 );
not ( n15826 , n15822 );
not ( n15827 , n15823 );
and ( n15828 , n15826 , n15827 );
nor ( n15829 , n15825 , n15828 );
xnor ( n15830 , n15820 , n15829 );
not ( n15831 , n15830 );
or ( n15832 , n15796 , n15831 );
or ( n15833 , n15830 , n15795 );
nand ( n15834 , n15832 , n15833 );
not ( n15835 , n15834 );
and ( n15836 , n15794 , n15835 );
not ( n15837 , n15769 );
not ( n15838 , n15792 );
not ( n15839 , n15838 );
or ( n15840 , n15837 , n15839 );
nand ( n15841 , n15792 , n15770 );
nand ( n15842 , n15840 , n15841 );
not ( n15843 , n15842 );
and ( n15844 , n15843 , n15834 );
nor ( n15845 , n15836 , n15844 );
buf ( n15846 , n5757 );
buf ( n15847 , n15846 );
nand ( n15848 , n8581 , n15847 );
not ( n15849 , n15848 );
not ( n15850 , n8580 );
nor ( n15851 , n15850 , n15847 );
nor ( n15852 , n15849 , n15851 );
not ( n15853 , n15852 );
not ( n15854 , n8612 );
or ( n15855 , n15853 , n15854 );
or ( n15856 , n8612 , n15852 );
nand ( n15857 , n15855 , n15856 );
nand ( n15858 , n15845 , n15857 );
not ( n15859 , n15858 );
buf ( n15860 , n5758 );
buf ( n15861 , n15860 );
not ( n15862 , n15861 );
buf ( n15863 , n5759 );
not ( n15864 , n15863 );
not ( n15865 , n15864 );
or ( n15866 , n15862 , n15865 );
not ( n15867 , n15860 );
buf ( n15868 , n15863 );
nand ( n15869 , n15867 , n15868 );
nand ( n15870 , n15866 , n15869 );
buf ( n15871 , n5760 );
buf ( n15872 , n15871 );
and ( n15873 , n15870 , n15872 );
not ( n15874 , n15870 );
not ( n15875 , n15871 );
and ( n15876 , n15874 , n15875 );
nor ( n15877 , n15873 , n15876 );
buf ( n15878 , n5761 );
nand ( n15879 , n7477 , n15878 );
buf ( n15880 , n5762 );
buf ( n15881 , n15880 );
and ( n15882 , n15879 , n15881 );
not ( n15883 , n15879 );
not ( n15884 , n15880 );
and ( n15885 , n15883 , n15884 );
nor ( n15886 , n15882 , n15885 );
xor ( n15887 , n15877 , n15886 );
buf ( n15888 , n5763 );
nand ( n15889 , n10204 , n15888 );
buf ( n15890 , n5764 );
not ( n15891 , n15890 );
and ( n15892 , n15889 , n15891 );
not ( n15893 , n15889 );
buf ( n15894 , n15890 );
and ( n15895 , n15893 , n15894 );
nor ( n15896 , n15892 , n15895 );
buf ( n15897 , n15896 );
xnor ( n15898 , n15887 , n15897 );
not ( n15899 , n15898 );
buf ( n15900 , n8690 );
not ( n15901 , n15900 );
and ( n15902 , n15899 , n15901 );
and ( n15903 , n15898 , n15900 );
nor ( n15904 , n15902 , n15903 );
buf ( n15905 , n5765 );
buf ( n15906 , n15905 );
not ( n15907 , n15906 );
buf ( n15908 , n5766 );
not ( n15909 , n15908 );
not ( n15910 , n15909 );
or ( n15911 , n15907 , n15910 );
not ( n15912 , n15905 );
buf ( n15913 , n15908 );
nand ( n15914 , n15912 , n15913 );
nand ( n15915 , n15911 , n15914 );
buf ( n15916 , n5767 );
not ( n15917 , n15916 );
and ( n15918 , n15915 , n15917 );
not ( n15919 , n15915 );
buf ( n15920 , n15916 );
and ( n15921 , n15919 , n15920 );
nor ( n15922 , n15918 , n15921 );
buf ( n15923 , n5768 );
nand ( n15924 , n7401 , n15923 );
buf ( n15925 , n5769 );
buf ( n15926 , n15925 );
and ( n15927 , n15924 , n15926 );
not ( n15928 , n15924 );
not ( n15929 , n15925 );
and ( n15930 , n15928 , n15929 );
nor ( n15931 , n15927 , n15930 );
xor ( n15932 , n15922 , n15931 );
xnor ( n15933 , n15932 , n8104 );
buf ( n15934 , n15933 );
and ( n15935 , n15904 , n15934 );
not ( n15936 , n15904 );
buf ( n15937 , n15934 );
not ( n15938 , n15937 );
and ( n15939 , n15936 , n15938 );
nor ( n15940 , n15935 , n15939 );
not ( n15941 , n15940 );
and ( n15942 , n15859 , n15941 );
and ( n15943 , n15858 , n15940 );
nor ( n15944 , n15942 , n15943 );
not ( n15945 , n15944 );
or ( n15946 , n15758 , n15945 );
or ( n15947 , n15944 , n15757 );
nand ( n15948 , n15946 , n15947 );
buf ( n15949 , n14418 );
buf ( n15950 , n5770 );
buf ( n15951 , n15950 );
not ( n15952 , n15951 );
buf ( n15953 , n5771 );
not ( n15954 , n15953 );
not ( n15955 , n15954 );
or ( n15956 , n15952 , n15955 );
not ( n15957 , n15950 );
buf ( n15958 , n15953 );
nand ( n15959 , n15957 , n15958 );
nand ( n15960 , n15956 , n15959 );
buf ( n15961 , n5772 );
not ( n15962 , n15961 );
and ( n15963 , n15960 , n15962 );
not ( n15964 , n15960 );
buf ( n15965 , n15961 );
and ( n15966 , n15964 , n15965 );
nor ( n15967 , n15963 , n15966 );
buf ( n15968 , n5773 );
nand ( n15969 , n7401 , n15968 );
buf ( n15970 , n5774 );
buf ( n15971 , n15970 );
and ( n15972 , n15969 , n15971 );
not ( n15973 , n15969 );
not ( n15974 , n15970 );
and ( n15975 , n15973 , n15974 );
nor ( n15976 , n15972 , n15975 );
xor ( n15977 , n15967 , n15976 );
buf ( n15978 , n5775 );
nand ( n15979 , n7356 , n15978 );
buf ( n15980 , n5776 );
not ( n15981 , n15980 );
and ( n15982 , n15979 , n15981 );
not ( n15983 , n15979 );
buf ( n15984 , n15980 );
and ( n15985 , n15983 , n15984 );
nor ( n15986 , n15982 , n15985 );
xor ( n15987 , n15977 , n15986 );
buf ( n15988 , n15987 );
buf ( n15989 , n15988 );
xor ( n15990 , n15949 , n15989 );
buf ( n15991 , n10734 );
xnor ( n15992 , n15990 , n15991 );
not ( n15993 , n15992 );
buf ( n15994 , n5777 );
buf ( n15995 , n15994 );
not ( n15996 , n15995 );
not ( n15997 , n11269 );
or ( n15998 , n15996 , n15997 );
or ( n15999 , n11269 , n15995 );
nand ( n16000 , n15998 , n15999 );
and ( n16001 , n16000 , n11229 );
not ( n16002 , n16000 );
not ( n16003 , n11229 );
and ( n16004 , n16002 , n16003 );
nor ( n16005 , n16001 , n16004 );
not ( n16006 , n16005 );
nand ( n16007 , n15993 , n16006 );
not ( n16008 , n10641 );
buf ( n16009 , n5778 );
nand ( n16010 , n6817 , n16009 );
buf ( n16011 , n16010 );
buf ( n16012 , n5779 );
xor ( n16013 , n16011 , n16012 );
not ( n16014 , n16013 );
not ( n16015 , n10588 );
or ( n16016 , n16014 , n16015 );
or ( n16017 , n10588 , n16013 );
nand ( n16018 , n16016 , n16017 );
not ( n16019 , n16018 );
or ( n16020 , n16008 , n16019 );
or ( n16021 , n16018 , n10641 );
nand ( n16022 , n16020 , n16021 );
not ( n16023 , n16022 );
and ( n16024 , n16007 , n16023 );
not ( n16025 , n16007 );
and ( n16026 , n16025 , n16022 );
nor ( n16027 , n16024 , n16026 );
not ( n16028 , n16027 );
and ( n16029 , n15948 , n16028 );
not ( n16030 , n15948 );
and ( n16031 , n16030 , n16027 );
nor ( n16032 , n16029 , n16031 );
not ( n16033 , n16032 );
buf ( n16034 , n5780 );
nand ( n16035 , n7094 , n16034 );
buf ( n16036 , n5781 );
buf ( n16037 , n16036 );
and ( n16038 , n16035 , n16037 );
not ( n16039 , n16035 );
not ( n16040 , n16036 );
and ( n16041 , n16039 , n16040 );
nor ( n16042 , n16038 , n16041 );
buf ( n16043 , n16042 );
not ( n16044 , n16043 );
not ( n16045 , n7931 );
or ( n16046 , n16044 , n16045 );
or ( n16047 , n7931 , n16043 );
nand ( n16048 , n16046 , n16047 );
and ( n16049 , n16048 , n7977 );
not ( n16050 , n16048 );
and ( n16051 , n16050 , n7970 );
nor ( n16052 , n16049 , n16051 );
buf ( n16053 , n16052 );
not ( n16054 , n16053 );
buf ( n16055 , n5782 );
buf ( n16056 , n16055 );
not ( n16057 , n16056 );
buf ( n16058 , n5783 );
not ( n16059 , n16058 );
not ( n16060 , n16059 );
or ( n16061 , n16057 , n16060 );
not ( n16062 , n16055 );
buf ( n16063 , n16058 );
nand ( n16064 , n16062 , n16063 );
nand ( n16065 , n16061 , n16064 );
buf ( n16066 , n5784 );
buf ( n16067 , n16066 );
and ( n16068 , n16065 , n16067 );
not ( n16069 , n16065 );
not ( n16070 , n16066 );
and ( n16071 , n16069 , n16070 );
nor ( n16072 , n16068 , n16071 );
buf ( n16073 , n5785 );
nand ( n16074 , n6804 , n16073 );
buf ( n16075 , n5786 );
not ( n16076 , n16075 );
and ( n16077 , n16074 , n16076 );
not ( n16078 , n16074 );
buf ( n16079 , n16075 );
and ( n16080 , n16078 , n16079 );
nor ( n16081 , n16077 , n16080 );
xor ( n16082 , n16072 , n16081 );
buf ( n16083 , n5787 );
nand ( n16084 , n8971 , n16083 );
buf ( n16085 , n5788 );
not ( n16086 , n16085 );
and ( n16087 , n16084 , n16086 );
not ( n16088 , n16084 );
buf ( n16089 , n16085 );
and ( n16090 , n16088 , n16089 );
nor ( n16091 , n16087 , n16090 );
xnor ( n16092 , n16082 , n16091 );
buf ( n16093 , n16092 );
not ( n16094 , n16093 );
buf ( n16095 , n5789 );
not ( n16096 , n16095 );
xor ( n16097 , n9148 , n9157 );
xnor ( n16098 , n16097 , n9168 );
not ( n16099 , n16098 );
or ( n16100 , n16096 , n16099 );
or ( n16101 , n16098 , n16095 );
nand ( n16102 , n16100 , n16101 );
not ( n16103 , n16102 );
or ( n16104 , n16094 , n16103 );
or ( n16105 , n16102 , n16093 );
nand ( n16106 , n16104 , n16105 );
not ( n16107 , n16106 );
not ( n16108 , n12602 );
buf ( n16109 , n5790 );
buf ( n16110 , n5791 );
buf ( n16111 , n16110 );
not ( n16112 , n16111 );
buf ( n16113 , n5792 );
not ( n16114 , n16113 );
not ( n16115 , n16114 );
or ( n16116 , n16112 , n16115 );
not ( n16117 , n16110 );
buf ( n16118 , n16113 );
nand ( n16119 , n16117 , n16118 );
nand ( n16120 , n16116 , n16119 );
xor ( n16121 , n16109 , n16120 );
not ( n16122 , n13083 );
buf ( n16123 , n5793 );
nand ( n16124 , n7865 , n16123 );
buf ( n16125 , n5794 );
buf ( n16126 , n16125 );
and ( n16127 , n16124 , n16126 );
not ( n16128 , n16124 );
not ( n16129 , n16125 );
and ( n16130 , n16128 , n16129 );
nor ( n16131 , n16127 , n16130 );
not ( n16132 , n16131 );
not ( n16133 , n16132 );
or ( n16134 , n16122 , n16133 );
nand ( n16135 , n16131 , n13079 );
nand ( n16136 , n16134 , n16135 );
xor ( n16137 , n16121 , n16136 );
not ( n16138 , n16137 );
or ( n16139 , n16108 , n16138 );
not ( n16140 , n12602 );
xor ( n16141 , n16109 , n16120 );
xnor ( n16142 , n16141 , n16136 );
nand ( n16143 , n16140 , n16142 );
nand ( n16144 , n16139 , n16143 );
buf ( n16145 , n5795 );
buf ( n16146 , n16145 );
not ( n16147 , n16146 );
buf ( n16148 , n5796 );
not ( n16149 , n16148 );
not ( n16150 , n16149 );
or ( n16151 , n16147 , n16150 );
not ( n16152 , n16145 );
buf ( n16153 , n16148 );
nand ( n16154 , n16152 , n16153 );
nand ( n16155 , n16151 , n16154 );
buf ( n16156 , n5797 );
not ( n16157 , n16156 );
and ( n16158 , n16155 , n16157 );
not ( n16159 , n16155 );
buf ( n16160 , n16156 );
and ( n16161 , n16159 , n16160 );
nor ( n16162 , n16158 , n16161 );
buf ( n16163 , n5798 );
nand ( n16164 , n7412 , n16163 );
buf ( n16165 , n5799 );
buf ( n16166 , n16165 );
and ( n16167 , n16164 , n16166 );
not ( n16168 , n16164 );
not ( n16169 , n16165 );
and ( n16170 , n16168 , n16169 );
nor ( n16171 , n16167 , n16170 );
xor ( n16172 , n16162 , n16171 );
buf ( n16173 , n5800 );
nand ( n16174 , n8821 , n16173 );
buf ( n16175 , n5801 );
buf ( n16176 , n16175 );
and ( n16177 , n16174 , n16176 );
not ( n16178 , n16174 );
not ( n16179 , n16175 );
and ( n16180 , n16178 , n16179 );
nor ( n16181 , n16177 , n16180 );
xnor ( n16182 , n16172 , n16181 );
buf ( n16183 , n16182 );
not ( n16184 , n16183 );
and ( n16185 , n16144 , n16184 );
not ( n16186 , n16144 );
and ( n16187 , n16186 , n16183 );
nor ( n16188 , n16185 , n16187 );
not ( n16189 , n16188 );
nand ( n16190 , n16107 , n16189 );
not ( n16191 , n16190 );
or ( n16192 , n16054 , n16191 );
or ( n16193 , n16190 , n16053 );
nand ( n16194 , n16192 , n16193 );
not ( n16195 , n16194 );
not ( n16196 , n15463 );
nand ( n16197 , n16196 , n15554 );
not ( n16198 , n16197 );
buf ( n16199 , n5802 );
nand ( n16200 , n6985 , n16199 );
buf ( n16201 , n5803 );
not ( n16202 , n16201 );
and ( n16203 , n16200 , n16202 );
not ( n16204 , n16200 );
buf ( n16205 , n16201 );
and ( n16206 , n16204 , n16205 );
nor ( n16207 , n16203 , n16206 );
not ( n16208 , n16207 );
not ( n16209 , n12525 );
or ( n16210 , n16208 , n16209 );
not ( n16211 , n16207 );
not ( n16212 , n12524 );
nand ( n16213 , n16211 , n16212 );
nand ( n16214 , n16210 , n16213 );
and ( n16215 , n16214 , n12531 );
not ( n16216 , n16214 );
and ( n16217 , n16216 , n12532 );
nor ( n16218 , n16215 , n16217 );
buf ( n16219 , n16218 );
not ( n16220 , n16219 );
or ( n16221 , n16198 , n16220 );
or ( n16222 , n16219 , n16197 );
nand ( n16223 , n16221 , n16222 );
not ( n16224 , n16223 );
not ( n16225 , n16224 );
or ( n16226 , n16195 , n16225 );
not ( n16227 , n16194 );
nand ( n16228 , n16227 , n16223 );
nand ( n16229 , n16226 , n16228 );
not ( n16230 , n16229 );
and ( n16231 , n16033 , n16230 );
not ( n16232 , n16033 );
not ( n16233 , n16230 );
and ( n16234 , n16232 , n16233 );
nor ( n16235 , n16231 , n16234 );
not ( n16236 , n16235 );
or ( n16237 , n15556 , n16236 );
not ( n16238 , n15555 );
not ( n16239 , n16229 );
not ( n16240 , n16032 );
or ( n16241 , n16239 , n16240 );
nand ( n16242 , n16033 , n16230 );
nand ( n16243 , n16241 , n16242 );
nand ( n16244 , n16238 , n16243 );
nand ( n16245 , n16237 , n16244 );
buf ( n16246 , n5804 );
buf ( n16247 , n16246 );
not ( n16248 , n16247 );
not ( n16249 , n11868 );
or ( n16250 , n16248 , n16249 );
or ( n16251 , n11868 , n16247 );
nand ( n16252 , n16250 , n16251 );
buf ( n16253 , n5805 );
buf ( n16254 , n16253 );
not ( n16255 , n16254 );
buf ( n16256 , n5806 );
not ( n16257 , n16256 );
not ( n16258 , n16257 );
or ( n16259 , n16255 , n16258 );
not ( n16260 , n16253 );
buf ( n16261 , n16256 );
nand ( n16262 , n16260 , n16261 );
nand ( n16263 , n16259 , n16262 );
not ( n16264 , n16263 );
buf ( n16265 , n5807 );
buf ( n16266 , n5808 );
not ( n16267 , n16266 );
xor ( n16268 , n16265 , n16267 );
buf ( n16269 , n5809 );
not ( n16270 , n16269 );
buf ( n16271 , n5810 );
nand ( n16272 , n6660 , n16271 );
not ( n16273 , n16272 );
or ( n16274 , n16270 , n16273 );
nand ( n16275 , n12401 , n16271 );
or ( n16276 , n16275 , n16269 );
nand ( n16277 , n16274 , n16276 );
xnor ( n16278 , n16268 , n16277 );
not ( n16279 , n16278 );
not ( n16280 , n16279 );
or ( n16281 , n16264 , n16280 );
not ( n16282 , n16263 );
nand ( n16283 , n16278 , n16282 );
nand ( n16284 , n16281 , n16283 );
buf ( n16285 , n16284 );
buf ( n16286 , n16285 );
and ( n16287 , n16252 , n16286 );
not ( n16288 , n16252 );
not ( n16289 , n16285 );
and ( n16290 , n16288 , n16289 );
nor ( n16291 , n16287 , n16290 );
buf ( n16292 , n5811 );
buf ( n16293 , n16292 );
not ( n16294 , n16293 );
buf ( n16295 , n15183 );
not ( n16296 , n16295 );
or ( n16297 , n16294 , n16296 );
or ( n16298 , n16295 , n16293 );
nand ( n16299 , n16297 , n16298 );
buf ( n16300 , n14921 );
and ( n16301 , n16299 , n16300 );
not ( n16302 , n16299 );
not ( n16303 , n16300 );
and ( n16304 , n16302 , n16303 );
nor ( n16305 , n16301 , n16304 );
nand ( n16306 , n16291 , n16305 );
not ( n16307 , n16306 );
not ( n16308 , n10509 );
not ( n16309 , n14055 );
not ( n16310 , n16309 );
or ( n16311 , n16308 , n16310 );
not ( n16312 , n16309 );
nand ( n16313 , n16312 , n10505 );
nand ( n16314 , n16311 , n16313 );
buf ( n16315 , n5812 );
buf ( n16316 , n16315 );
not ( n16317 , n16316 );
buf ( n16318 , n5813 );
not ( n16319 , n16318 );
not ( n16320 , n16319 );
or ( n16321 , n16317 , n16320 );
not ( n16322 , n16315 );
buf ( n16323 , n16318 );
nand ( n16324 , n16322 , n16323 );
nand ( n16325 , n16321 , n16324 );
buf ( n16326 , n5814 );
not ( n16327 , n16326 );
and ( n16328 , n16325 , n16327 );
not ( n16329 , n16325 );
buf ( n16330 , n16326 );
and ( n16331 , n16329 , n16330 );
nor ( n16332 , n16328 , n16331 );
not ( n16333 , n16332 );
buf ( n16334 , n5815 );
nand ( n16335 , n8343 , n16334 );
buf ( n16336 , n5816 );
buf ( n16337 , n16336 );
and ( n16338 , n16335 , n16337 );
not ( n16339 , n16335 );
not ( n16340 , n16336 );
and ( n16341 , n16339 , n16340 );
nor ( n16342 , n16338 , n16341 );
not ( n16343 , n16342 );
buf ( n16344 , n5817 );
nand ( n16345 , n7195 , n16344 );
buf ( n16346 , n5818 );
not ( n16347 , n16346 );
xor ( n16348 , n16345 , n16347 );
not ( n16349 , n16348 );
or ( n16350 , n16343 , n16349 );
or ( n16351 , n16342 , n16348 );
nand ( n16352 , n16350 , n16351 );
not ( n16353 , n16352 );
or ( n16354 , n16333 , n16353 );
or ( n16355 , n16352 , n16332 );
nand ( n16356 , n16354 , n16355 );
buf ( n16357 , n16356 );
and ( n16358 , n16314 , n16357 );
not ( n16359 , n16314 );
xor ( n16360 , n16332 , n16342 );
xnor ( n16361 , n16360 , n16348 );
not ( n16362 , n16361 );
not ( n16363 , n16362 );
and ( n16364 , n16359 , n16363 );
nor ( n16365 , n16358 , n16364 );
not ( n16366 , n16365 );
and ( n16367 , n16307 , n16366 );
and ( n16368 , n16306 , n16365 );
nor ( n16369 , n16367 , n16368 );
not ( n16370 , n16369 );
buf ( n16371 , n13329 );
xor ( n16372 , n16371 , n11269 );
buf ( n16373 , n11923 );
not ( n16374 , n16373 );
xnor ( n16375 , n16372 , n16374 );
xor ( n16376 , n8503 , n13548 );
not ( n16377 , n13572 );
xnor ( n16378 , n16376 , n16377 );
not ( n16379 , n16378 );
nand ( n16380 , n16375 , n16379 );
buf ( n16381 , n5819 );
buf ( n16382 , n16381 );
not ( n16383 , n16382 );
buf ( n16384 , n5820 );
buf ( n16385 , n16384 );
not ( n16386 , n16385 );
not ( n16387 , n12845 );
not ( n16388 , n16387 );
or ( n16389 , n16386 , n16388 );
not ( n16390 , n16384 );
nand ( n16391 , n16390 , n12846 );
nand ( n16392 , n16389 , n16391 );
buf ( n16393 , n5821 );
buf ( n16394 , n16393 );
and ( n16395 , n16392 , n16394 );
not ( n16396 , n16392 );
not ( n16397 , n16393 );
and ( n16398 , n16396 , n16397 );
nor ( n16399 , n16395 , n16398 );
buf ( n16400 , n5822 );
nand ( n16401 , n7093 , n16400 );
buf ( n16402 , n5823 );
not ( n16403 , n16402 );
and ( n16404 , n16401 , n16403 );
not ( n16405 , n16401 );
buf ( n16406 , n16402 );
and ( n16407 , n16405 , n16406 );
nor ( n16408 , n16404 , n16407 );
xor ( n16409 , n16399 , n16408 );
buf ( n16410 , n5824 );
nand ( n16411 , n10204 , n16410 );
buf ( n16412 , n5825 );
not ( n16413 , n16412 );
and ( n16414 , n16411 , n16413 );
not ( n16415 , n16411 );
buf ( n16416 , n16412 );
and ( n16417 , n16415 , n16416 );
nor ( n16418 , n16414 , n16417 );
xnor ( n16419 , n16409 , n16418 );
buf ( n16420 , n16419 );
not ( n16421 , n16420 );
or ( n16422 , n16383 , n16421 );
or ( n16423 , n16420 , n16382 );
nand ( n16424 , n16422 , n16423 );
buf ( n16425 , n5826 );
buf ( n16426 , n16425 );
buf ( n16427 , n5827 );
buf ( n16428 , n16427 );
not ( n16429 , n16428 );
buf ( n16430 , n5828 );
not ( n16431 , n16430 );
not ( n16432 , n16431 );
or ( n16433 , n16429 , n16432 );
not ( n16434 , n16427 );
buf ( n16435 , n16430 );
nand ( n16436 , n16434 , n16435 );
nand ( n16437 , n16433 , n16436 );
xor ( n16438 , n16426 , n16437 );
xor ( n16439 , n10547 , n16012 );
xnor ( n16440 , n16439 , n16010 );
xnor ( n16441 , n16438 , n16440 );
buf ( n16442 , n16441 );
not ( n16443 , n16442 );
and ( n16444 , n16424 , n16443 );
not ( n16445 , n16424 );
buf ( n16446 , n16442 );
and ( n16447 , n16445 , n16446 );
nor ( n16448 , n16444 , n16447 );
not ( n16449 , n16448 );
and ( n16450 , n16380 , n16449 );
not ( n16451 , n16380 );
and ( n16452 , n16451 , n16448 );
nor ( n16453 , n16450 , n16452 );
not ( n16454 , n16453 );
or ( n16455 , n16370 , n16454 );
or ( n16456 , n16453 , n16369 );
nand ( n16457 , n16455 , n16456 );
not ( n16458 , n6786 );
buf ( n16459 , n5829 );
buf ( n16460 , n16459 );
not ( n16461 , n16460 );
buf ( n16462 , n5830 );
not ( n16463 , n16462 );
not ( n16464 , n16463 );
or ( n16465 , n16461 , n16464 );
not ( n16466 , n16459 );
buf ( n16467 , n16462 );
nand ( n16468 , n16466 , n16467 );
nand ( n16469 , n16465 , n16468 );
buf ( n16470 , n5831 );
buf ( n16471 , n16470 );
and ( n16472 , n16469 , n16471 );
not ( n16473 , n16469 );
not ( n16474 , n16470 );
and ( n16475 , n16473 , n16474 );
nor ( n16476 , n16472 , n16475 );
xor ( n16477 , n16476 , n12217 );
buf ( n16478 , n5832 );
nand ( n16479 , n7785 , n16478 );
buf ( n16480 , n5833 );
not ( n16481 , n16480 );
and ( n16482 , n16479 , n16481 );
not ( n16483 , n16479 );
buf ( n16484 , n16480 );
and ( n16485 , n16483 , n16484 );
nor ( n16486 , n16482 , n16485 );
xnor ( n16487 , n16477 , n16486 );
buf ( n16488 , n16487 );
not ( n16489 , n16488 );
or ( n16490 , n16458 , n16489 );
not ( n16491 , n16487 );
not ( n16492 , n16491 );
or ( n16493 , n16492 , n6786 );
nand ( n16494 , n16490 , n16493 );
buf ( n16495 , n5834 );
buf ( n16496 , n16495 );
not ( n16497 , n16496 );
buf ( n16498 , n5835 );
not ( n16499 , n16498 );
not ( n16500 , n16499 );
or ( n16501 , n16497 , n16500 );
not ( n16502 , n16495 );
buf ( n16503 , n16498 );
nand ( n16504 , n16502 , n16503 );
nand ( n16505 , n16501 , n16504 );
buf ( n16506 , n5836 );
not ( n16507 , n16506 );
and ( n16508 , n16505 , n16507 );
not ( n16509 , n16505 );
buf ( n16510 , n16506 );
and ( n16511 , n16509 , n16510 );
nor ( n16512 , n16508 , n16511 );
buf ( n16513 , n5837 );
nand ( n16514 , n7183 , n16513 );
buf ( n16515 , n5838 );
not ( n16516 , n16515 );
and ( n16517 , n16514 , n16516 );
not ( n16518 , n16514 );
buf ( n16519 , n16515 );
and ( n16520 , n16518 , n16519 );
nor ( n16521 , n16517 , n16520 );
xor ( n16522 , n16512 , n16521 );
buf ( n16523 , n5839 );
nand ( n16524 , n7515 , n16523 );
buf ( n16525 , n5840 );
buf ( n16526 , n16525 );
and ( n16527 , n16524 , n16526 );
not ( n16528 , n16524 );
not ( n16529 , n16525 );
and ( n16530 , n16528 , n16529 );
nor ( n16531 , n16527 , n16530 );
xor ( n16532 , n16522 , n16531 );
not ( n16533 , n16532 );
and ( n16534 , n16494 , n16533 );
not ( n16535 , n16494 );
not ( n16536 , n16532 );
not ( n16537 , n16536 );
not ( n16538 , n16537 );
not ( n16539 , n16538 );
and ( n16540 , n16535 , n16539 );
nor ( n16541 , n16534 , n16540 );
not ( n16542 , n9575 );
not ( n16543 , n15560 );
or ( n16544 , n16542 , n16543 );
not ( n16545 , n9575 );
nand ( n16546 , n16545 , n15561 );
nand ( n16547 , n16544 , n16546 );
and ( n16548 , n16547 , n15568 );
not ( n16549 , n16547 );
and ( n16550 , n16549 , n13708 );
nor ( n16551 , n16548 , n16550 );
nand ( n16552 , n16541 , n16551 );
not ( n16553 , n16552 );
xor ( n16554 , n8356 , n8365 );
xnor ( n16555 , n16554 , n8381 );
xor ( n16556 , n13100 , n16555 );
and ( n16557 , n16556 , n8441 );
not ( n16558 , n16556 );
and ( n16559 , n16558 , n8434 );
nor ( n16560 , n16557 , n16559 );
not ( n16561 , n16560 );
not ( n16562 , n16561 );
and ( n16563 , n16553 , n16562 );
and ( n16564 , n16552 , n16561 );
nor ( n16565 , n16563 , n16564 );
not ( n16566 , n16565 );
buf ( n16567 , n5841 );
buf ( n16568 , n5842 );
buf ( n16569 , n16568 );
not ( n16570 , n16569 );
buf ( n16571 , n5843 );
not ( n16572 , n16571 );
not ( n16573 , n16572 );
or ( n16574 , n16570 , n16573 );
not ( n16575 , n16568 );
buf ( n16576 , n16571 );
nand ( n16577 , n16575 , n16576 );
nand ( n16578 , n16574 , n16577 );
xor ( n16579 , n16567 , n16578 );
buf ( n16580 , n5844 );
xor ( n16581 , n7063 , n16580 );
buf ( n16582 , n5845 );
nand ( n16583 , n6906 , n16582 );
xnor ( n16584 , n16581 , n16583 );
xnor ( n16585 , n16579 , n16584 );
not ( n16586 , n16585 );
not ( n16587 , n11598 );
buf ( n16588 , n5846 );
buf ( n16589 , n16588 );
not ( n16590 , n16589 );
buf ( n16591 , n5847 );
not ( n16592 , n16591 );
not ( n16593 , n16592 );
or ( n16594 , n16590 , n16593 );
not ( n16595 , n16588 );
buf ( n16596 , n16591 );
nand ( n16597 , n16595 , n16596 );
nand ( n16598 , n16594 , n16597 );
buf ( n16599 , n5848 );
buf ( n16600 , n16599 );
and ( n16601 , n16598 , n16600 );
not ( n16602 , n16598 );
not ( n16603 , n16599 );
and ( n16604 , n16602 , n16603 );
nor ( n16605 , n16601 , n16604 );
buf ( n16606 , n5849 );
nand ( n16607 , n8223 , n16606 );
buf ( n16608 , n5850 );
buf ( n16609 , n16608 );
and ( n16610 , n16607 , n16609 );
not ( n16611 , n16607 );
not ( n16612 , n16608 );
and ( n16613 , n16611 , n16612 );
nor ( n16614 , n16610 , n16613 );
xor ( n16615 , n16605 , n16614 );
buf ( n16616 , n5851 );
nand ( n16617 , n7082 , n16616 );
buf ( n16618 , n5852 );
not ( n16619 , n16618 );
and ( n16620 , n16617 , n16619 );
not ( n16621 , n16617 );
buf ( n16622 , n16618 );
and ( n16623 , n16621 , n16622 );
nor ( n16624 , n16620 , n16623 );
xnor ( n16625 , n16615 , n16624 );
not ( n16626 , n16625 );
not ( n16627 , n16626 );
or ( n16628 , n16587 , n16627 );
or ( n16629 , n16626 , n11598 );
nand ( n16630 , n16628 , n16629 );
and ( n16631 , n16586 , n16630 );
not ( n16632 , n16586 );
not ( n16633 , n16630 );
and ( n16634 , n16632 , n16633 );
nor ( n16635 , n16631 , n16634 );
not ( n16636 , n16635 );
buf ( n16637 , n5853 );
buf ( n16638 , n16637 );
not ( n16639 , n16638 );
buf ( n16640 , n5854 );
not ( n16641 , n16640 );
not ( n16642 , n16641 );
or ( n16643 , n16639 , n16642 );
not ( n16644 , n16637 );
buf ( n16645 , n16640 );
nand ( n16646 , n16644 , n16645 );
nand ( n16647 , n16643 , n16646 );
buf ( n16648 , n5855 );
not ( n16649 , n16648 );
and ( n16650 , n16647 , n16649 );
not ( n16651 , n16647 );
buf ( n16652 , n16648 );
and ( n16653 , n16651 , n16652 );
nor ( n16654 , n16650 , n16653 );
buf ( n16655 , n5856 );
nand ( n16656 , n7477 , n16655 );
buf ( n16657 , n5857 );
buf ( n16658 , n16657 );
and ( n16659 , n16656 , n16658 );
not ( n16660 , n16656 );
not ( n16661 , n16657 );
and ( n16662 , n16660 , n16661 );
nor ( n16663 , n16659 , n16662 );
xor ( n16664 , n16654 , n16663 );
buf ( n16665 , n5858 );
nand ( n16666 , n6863 , n16665 );
buf ( n16667 , n5859 );
not ( n16668 , n16667 );
and ( n16669 , n16666 , n16668 );
not ( n16670 , n16666 );
buf ( n16671 , n16667 );
and ( n16672 , n16670 , n16671 );
nor ( n16673 , n16669 , n16672 );
xnor ( n16674 , n16664 , n16673 );
not ( n16675 , n16674 );
buf ( n16676 , n15186 );
not ( n16677 , n16676 );
and ( n16678 , n16675 , n16677 );
and ( n16679 , n16674 , n16676 );
nor ( n16680 , n16678 , n16679 );
buf ( n16681 , n5860 );
buf ( n16682 , n16681 );
not ( n16683 , n16682 );
buf ( n16684 , n5861 );
not ( n16685 , n16684 );
not ( n16686 , n16685 );
or ( n16687 , n16683 , n16686 );
not ( n16688 , n16681 );
buf ( n16689 , n16684 );
nand ( n16690 , n16688 , n16689 );
nand ( n16691 , n16687 , n16690 );
buf ( n16692 , n5862 );
not ( n16693 , n16692 );
and ( n16694 , n16691 , n16693 );
not ( n16695 , n16691 );
buf ( n16696 , n16692 );
and ( n16697 , n16695 , n16696 );
nor ( n16698 , n16694 , n16697 );
buf ( n16699 , n5863 );
nand ( n16700 , n7043 , n16699 );
buf ( n16701 , n5864 );
buf ( n16702 , n16701 );
and ( n16703 , n16700 , n16702 );
not ( n16704 , n16700 );
not ( n16705 , n16701 );
and ( n16706 , n16704 , n16705 );
nor ( n16707 , n16703 , n16706 );
xor ( n16708 , n16698 , n16707 );
buf ( n16709 , n5865 );
nand ( n16710 , n8785 , n16709 );
buf ( n16711 , n5866 );
buf ( n16712 , n16711 );
and ( n16713 , n16710 , n16712 );
not ( n16714 , n16710 );
not ( n16715 , n16711 );
and ( n16716 , n16714 , n16715 );
nor ( n16717 , n16713 , n16716 );
xnor ( n16718 , n16708 , n16717 );
buf ( n16719 , n16718 );
not ( n16720 , n16719 );
and ( n16721 , n16680 , n16720 );
not ( n16722 , n16680 );
and ( n16723 , n16722 , n16719 );
nor ( n16724 , n16721 , n16723 );
nand ( n16725 , n16636 , n16724 );
buf ( n16726 , n5867 );
buf ( n16727 , n16726 );
not ( n16728 , n16727 );
not ( n16729 , n11948 );
or ( n16730 , n16728 , n16729 );
not ( n16731 , n16726 );
nand ( n16732 , n9948 , n16731 );
nand ( n16733 , n16730 , n16732 );
not ( n16734 , n16733 );
not ( n16735 , n11997 );
and ( n16736 , n16734 , n16735 );
not ( n16737 , n11996 );
and ( n16738 , n16733 , n16737 );
nor ( n16739 , n16736 , n16738 );
and ( n16740 , n16725 , n16739 );
not ( n16741 , n16725 );
not ( n16742 , n16739 );
and ( n16743 , n16741 , n16742 );
nor ( n16744 , n16740 , n16743 );
not ( n16745 , n16744 );
or ( n16746 , n16566 , n16745 );
or ( n16747 , n16744 , n16565 );
nand ( n16748 , n16746 , n16747 );
buf ( n16749 , n5868 );
buf ( n16750 , n16749 );
not ( n16751 , n12743 );
not ( n16752 , n16751 );
xor ( n16753 , n16750 , n16752 );
buf ( n16754 , n5869 );
buf ( n16755 , n16754 );
not ( n16756 , n16755 );
not ( n16757 , n7430 );
or ( n16758 , n16756 , n16757 );
not ( n16759 , n16754 );
nand ( n16760 , n16759 , n7381 );
nand ( n16761 , n16758 , n16760 );
not ( n16762 , n16761 );
not ( n16763 , n16762 );
buf ( n16764 , n5870 );
buf ( n16765 , n5871 );
not ( n16766 , n16765 );
xor ( n16767 , n16764 , n16766 );
buf ( n16768 , n5872 );
not ( n16769 , n16768 );
buf ( n16770 , n5873 );
nand ( n16771 , n6607 , n16770 );
not ( n16772 , n16771 );
or ( n16773 , n16769 , n16772 );
nand ( n16774 , n7183 , n16770 );
or ( n16775 , n16774 , n16768 );
nand ( n16776 , n16773 , n16775 );
xnor ( n16777 , n16767 , n16776 );
not ( n16778 , n16777 );
or ( n16779 , n16763 , n16778 );
or ( n16780 , n16777 , n16762 );
nand ( n16781 , n16779 , n16780 );
buf ( n16782 , n16781 );
not ( n16783 , n16782 );
xnor ( n16784 , n16753 , n16783 );
nor ( n16785 , n12636 , n15093 );
not ( n16786 , n16785 );
nand ( n16787 , n12641 , n15093 );
nand ( n16788 , n16786 , n16787 );
not ( n16789 , n12924 );
xor ( n16790 , n12946 , n16789 );
buf ( n16791 , n12914 );
xnor ( n16792 , n16790 , n16791 );
buf ( n16793 , n16792 );
and ( n16794 , n16788 , n16793 );
not ( n16795 , n16788 );
buf ( n16796 , n12951 );
and ( n16797 , n16795 , n16796 );
nor ( n16798 , n16794 , n16797 );
nand ( n16799 , n16784 , n16798 );
not ( n16800 , n16799 );
buf ( n16801 , n13902 );
not ( n16802 , n16801 );
buf ( n16803 , n5874 );
not ( n16804 , n16803 );
not ( n16805 , n16804 );
not ( n16806 , n14213 );
or ( n16807 , n16805 , n16806 );
buf ( n16808 , n16803 );
nand ( n16809 , n14206 , n16808 );
nand ( n16810 , n16807 , n16809 );
not ( n16811 , n16810 );
or ( n16812 , n16802 , n16811 );
or ( n16813 , n16810 , n16801 );
nand ( n16814 , n16812 , n16813 );
not ( n16815 , n16814 );
and ( n16816 , n16800 , n16815 );
and ( n16817 , n16799 , n16814 );
nor ( n16818 , n16816 , n16817 );
and ( n16819 , n16748 , n16818 );
not ( n16820 , n16748 );
not ( n16821 , n16818 );
and ( n16822 , n16820 , n16821 );
nor ( n16823 , n16819 , n16822 );
and ( n16824 , n16457 , n16823 );
not ( n16825 , n16457 );
not ( n16826 , n16823 );
and ( n16827 , n16825 , n16826 );
nor ( n16828 , n16824 , n16827 );
not ( n16829 , n16828 );
not ( n16830 , n16829 );
and ( n16831 , n16245 , n16830 );
not ( n16832 , n16245 );
buf ( n16833 , n16828 );
not ( n16834 , n16833 );
and ( n16835 , n16832 , n16834 );
nor ( n16836 , n16831 , n16835 );
not ( n16837 , n13752 );
buf ( n16838 , n16837 );
not ( n16839 , n16838 );
nor ( n16840 , n16836 , n16839 );
nand ( n16841 , n9975 , n10174 );
not ( n16842 , n16841 );
not ( n16843 , n13685 );
buf ( n16844 , n14383 );
not ( n16845 , n16844 );
not ( n16846 , n16845 );
or ( n16847 , n16843 , n16846 );
nand ( n16848 , n16844 , n13682 );
nand ( n16849 , n16847 , n16848 );
buf ( n16850 , n12525 );
xnor ( n16851 , n16849 , n16850 );
not ( n16852 , n16851 );
and ( n16853 , n16842 , n16852 );
not ( n16854 , n10174 );
not ( n16855 , n16854 );
nand ( n16856 , n16855 , n9975 );
and ( n16857 , n16856 , n16851 );
nor ( n16858 , n16853 , n16857 );
not ( n16859 , n16858 );
not ( n16860 , n16859 );
not ( n16861 , n16183 );
and ( n16862 , n12944 , n16861 );
not ( n16863 , n12944 );
and ( n16864 , n16863 , n16183 );
or ( n16865 , n16862 , n16864 );
buf ( n16866 , n5875 );
buf ( n16867 , n16866 );
not ( n16868 , n16867 );
buf ( n16869 , n5876 );
not ( n16870 , n16869 );
not ( n16871 , n16870 );
or ( n16872 , n16868 , n16871 );
not ( n16873 , n16866 );
buf ( n16874 , n16869 );
nand ( n16875 , n16873 , n16874 );
nand ( n16876 , n16872 , n16875 );
not ( n16877 , n13759 );
and ( n16878 , n16876 , n16877 );
not ( n16879 , n16876 );
and ( n16880 , n16879 , n13760 );
nor ( n16881 , n16878 , n16880 );
buf ( n16882 , n5877 );
nand ( n16883 , n7981 , n16882 );
buf ( n16884 , n5878 );
buf ( n16885 , n16884 );
and ( n16886 , n16883 , n16885 );
not ( n16887 , n16883 );
not ( n16888 , n16884 );
and ( n16889 , n16887 , n16888 );
nor ( n16890 , n16886 , n16889 );
xor ( n16891 , n16881 , n16890 );
buf ( n16892 , n5879 );
nand ( n16893 , n6622 , n16892 );
buf ( n16894 , n5880 );
buf ( n16895 , n16894 );
and ( n16896 , n16893 , n16895 );
not ( n16897 , n16893 );
not ( n16898 , n16894 );
and ( n16899 , n16897 , n16898 );
nor ( n16900 , n16896 , n16899 );
xor ( n16901 , n16891 , n16900 );
buf ( n16902 , n16901 );
and ( n16903 , n16865 , n16902 );
not ( n16904 , n16865 );
not ( n16905 , n16902 );
and ( n16906 , n16904 , n16905 );
nor ( n16907 , n16903 , n16906 );
nand ( n16908 , n16907 , n10741 );
not ( n16909 , n16908 );
not ( n16910 , n12408 );
buf ( n16911 , n5881 );
buf ( n16912 , n16911 );
not ( n16913 , n16912 );
buf ( n16914 , n5882 );
not ( n16915 , n16914 );
not ( n16916 , n16915 );
or ( n16917 , n16913 , n16916 );
not ( n16918 , n16911 );
buf ( n16919 , n16914 );
nand ( n16920 , n16918 , n16919 );
nand ( n16921 , n16917 , n16920 );
buf ( n16922 , n5883 );
not ( n16923 , n16922 );
and ( n16924 , n16921 , n16923 );
not ( n16925 , n16921 );
buf ( n16926 , n16922 );
and ( n16927 , n16925 , n16926 );
nor ( n16928 , n16924 , n16927 );
buf ( n16929 , n5884 );
nand ( n16930 , n8387 , n16929 );
buf ( n16931 , n5885 );
buf ( n16932 , n16931 );
and ( n16933 , n16930 , n16932 );
not ( n16934 , n16930 );
not ( n16935 , n16931 );
and ( n16936 , n16934 , n16935 );
nor ( n16937 , n16933 , n16936 );
xor ( n16938 , n16928 , n16937 );
buf ( n16939 , n5886 );
nand ( n16940 , n7184 , n16939 );
buf ( n16941 , n5887 );
buf ( n16942 , n16941 );
and ( n16943 , n16940 , n16942 );
not ( n16944 , n16940 );
not ( n16945 , n16941 );
and ( n16946 , n16944 , n16945 );
nor ( n16947 , n16943 , n16946 );
xor ( n16948 , n16938 , n16947 );
not ( n16949 , n16948 );
or ( n16950 , n16910 , n16949 );
or ( n16951 , n16948 , n12408 );
nand ( n16952 , n16950 , n16951 );
and ( n16953 , n16952 , n15370 );
not ( n16954 , n16952 );
not ( n16955 , n15370 );
and ( n16956 , n16954 , n16955 );
nor ( n16957 , n16953 , n16956 );
not ( n16958 , n16957 );
and ( n16959 , n16909 , n16958 );
nand ( n16960 , n16907 , n10742 );
and ( n16961 , n16960 , n16957 );
nor ( n16962 , n16959 , n16961 );
not ( n16963 , n16962 );
not ( n16964 , n15442 );
not ( n16965 , n14670 );
or ( n16966 , n16964 , n16965 );
not ( n16967 , n15441 );
nand ( n16968 , n16967 , n14724 );
nand ( n16969 , n16966 , n16968 );
buf ( n16970 , n5888 );
buf ( n16971 , n16970 );
and ( n16972 , n16969 , n16971 );
not ( n16973 , n16969 );
not ( n16974 , n16970 );
and ( n16975 , n16973 , n16974 );
nor ( n16976 , n16972 , n16975 );
buf ( n16977 , n5889 );
nand ( n16978 , n7126 , n16977 );
buf ( n16979 , n5890 );
buf ( n16980 , n16979 );
and ( n16981 , n16978 , n16980 );
not ( n16982 , n16978 );
not ( n16983 , n16979 );
and ( n16984 , n16982 , n16983 );
nor ( n16985 , n16981 , n16984 );
xor ( n16986 , n16976 , n16985 );
buf ( n16987 , n5891 );
nand ( n16988 , n9159 , n16987 );
buf ( n16989 , n5892 );
not ( n16990 , n16989 );
and ( n16991 , n16988 , n16990 );
not ( n16992 , n16988 );
buf ( n16993 , n16989 );
and ( n16994 , n16992 , n16993 );
nor ( n16995 , n16991 , n16994 );
xnor ( n16996 , n16986 , n16995 );
not ( n16997 , n16996 );
not ( n16998 , n16997 );
buf ( n16999 , n5893 );
not ( n17000 , n16999 );
and ( n17001 , n16998 , n17000 );
buf ( n17002 , n16996 );
not ( n17003 , n17002 );
and ( n17004 , n17003 , n16999 );
nor ( n17005 , n17001 , n17004 );
buf ( n17006 , n5894 );
buf ( n17007 , n17006 );
not ( n17008 , n17007 );
buf ( n17009 , n5895 );
not ( n17010 , n17009 );
not ( n17011 , n17010 );
or ( n17012 , n17008 , n17011 );
not ( n17013 , n17006 );
buf ( n17014 , n17009 );
nand ( n17015 , n17013 , n17014 );
nand ( n17016 , n17012 , n17015 );
not ( n17017 , n9180 );
and ( n17018 , n17016 , n17017 );
not ( n17019 , n17016 );
and ( n17020 , n17019 , n9181 );
nor ( n17021 , n17018 , n17020 );
not ( n17022 , n17021 );
buf ( n17023 , n5896 );
nand ( n17024 , n7183 , n17023 );
buf ( n17025 , n5897 );
xor ( n17026 , n17024 , n17025 );
xor ( n17027 , n17022 , n17026 );
buf ( n17028 , n5898 );
nand ( n17029 , n7134 , n17028 );
buf ( n17030 , n5899 );
buf ( n17031 , n17030 );
and ( n17032 , n17029 , n17031 );
not ( n17033 , n17029 );
not ( n17034 , n17030 );
and ( n17035 , n17033 , n17034 );
nor ( n17036 , n17032 , n17035 );
xnor ( n17037 , n17027 , n17036 );
not ( n17038 , n17037 );
not ( n17039 , n17038 );
and ( n17040 , n17005 , n17039 );
not ( n17041 , n17005 );
xor ( n17042 , n17021 , n17026 );
xnor ( n17043 , n17042 , n17036 );
buf ( n17044 , n17043 );
and ( n17045 , n17041 , n17044 );
nor ( n17046 , n17040 , n17045 );
not ( n17047 , n17046 );
nand ( n17048 , n17047 , n10281 );
buf ( n17049 , n5900 );
buf ( n17050 , n17049 );
not ( n17051 , n17050 );
not ( n17052 , n13015 );
or ( n17053 , n17051 , n17052 );
not ( n17054 , n17050 );
nand ( n17055 , n17054 , n7931 );
nand ( n17056 , n17053 , n17055 );
not ( n17057 , n17056 );
not ( n17058 , n7970 );
and ( n17059 , n17057 , n17058 );
and ( n17060 , n7970 , n17056 );
nor ( n17061 , n17059 , n17060 );
and ( n17062 , n17048 , n17061 );
not ( n17063 , n17048 );
not ( n17064 , n17061 );
and ( n17065 , n17063 , n17064 );
nor ( n17066 , n17062 , n17065 );
not ( n17067 , n17066 );
or ( n17068 , n16963 , n17067 );
or ( n17069 , n17066 , n16962 );
nand ( n17070 , n17068 , n17069 );
not ( n17071 , n8008 );
buf ( n17072 , n5901 );
buf ( n17073 , n17072 );
not ( n17074 , n17073 );
buf ( n17075 , n5902 );
not ( n17076 , n17075 );
not ( n17077 , n17076 );
or ( n17078 , n17074 , n17077 );
not ( n17079 , n17072 );
buf ( n17080 , n17075 );
nand ( n17081 , n17079 , n17080 );
nand ( n17082 , n17078 , n17081 );
buf ( n17083 , n5903 );
not ( n17084 , n17083 );
and ( n17085 , n17082 , n17084 );
not ( n17086 , n17082 );
buf ( n17087 , n17083 );
and ( n17088 , n17086 , n17087 );
nor ( n17089 , n17085 , n17088 );
buf ( n17090 , n5904 );
nand ( n17091 , n7471 , n17090 );
buf ( n17092 , n5905 );
buf ( n17093 , n17092 );
and ( n17094 , n17091 , n17093 );
not ( n17095 , n17091 );
not ( n17096 , n17092 );
and ( n17097 , n17095 , n17096 );
nor ( n17098 , n17094 , n17097 );
xor ( n17099 , n17089 , n17098 );
buf ( n17100 , n5906 );
nand ( n17101 , n10577 , n17100 );
buf ( n17102 , n5907 );
not ( n17103 , n17102 );
and ( n17104 , n17101 , n17103 );
not ( n17105 , n17101 );
buf ( n17106 , n17102 );
and ( n17107 , n17105 , n17106 );
nor ( n17108 , n17104 , n17107 );
xnor ( n17109 , n17099 , n17108 );
not ( n17110 , n17109 );
or ( n17111 , n17071 , n17110 );
buf ( n17112 , n17109 );
or ( n17113 , n17112 , n8008 );
nand ( n17114 , n17111 , n17113 );
not ( n17115 , n17114 );
not ( n17116 , n17115 );
and ( n17117 , n12586 , n12551 );
not ( n17118 , n12586 );
buf ( n17119 , n12550 );
and ( n17120 , n17118 , n17119 );
nor ( n17121 , n17117 , n17120 );
not ( n17122 , n17121 );
and ( n17123 , n12560 , n17122 );
not ( n17124 , n12560 );
and ( n17125 , n17124 , n17121 );
nor ( n17126 , n17123 , n17125 );
not ( n17127 , n17126 );
not ( n17128 , n17127 );
or ( n17129 , n17116 , n17128 );
nand ( n17130 , n12587 , n17114 );
nand ( n17131 , n17129 , n17130 );
not ( n17132 , n17131 );
nand ( n17133 , n17132 , n9694 );
not ( n17134 , n9490 );
and ( n17135 , n17133 , n17134 );
not ( n17136 , n17133 );
and ( n17137 , n17136 , n9490 );
nor ( n17138 , n17135 , n17137 );
not ( n17139 , n17138 );
and ( n17140 , n17070 , n17139 );
not ( n17141 , n17070 );
and ( n17142 , n17141 , n17138 );
nor ( n17143 , n17140 , n17142 );
not ( n17144 , n17143 );
not ( n17145 , n16589 );
buf ( n17146 , n5908 );
nand ( n17147 , n8519 , n17146 );
buf ( n17148 , n5909 );
buf ( n17149 , n17148 );
and ( n17150 , n17147 , n17149 );
not ( n17151 , n17147 );
not ( n17152 , n17148 );
and ( n17153 , n17151 , n17152 );
nor ( n17154 , n17150 , n17153 );
not ( n17155 , n17154 );
buf ( n17156 , n5910 );
nand ( n17157 , n7955 , n17156 );
buf ( n17158 , n5911 );
not ( n17159 , n17158 );
and ( n17160 , n17157 , n17159 );
not ( n17161 , n17157 );
buf ( n17162 , n17158 );
and ( n17163 , n17161 , n17162 );
nor ( n17164 , n17160 , n17163 );
not ( n17165 , n17164 );
or ( n17166 , n17155 , n17165 );
or ( n17167 , n17154 , n17164 );
nand ( n17168 , n17166 , n17167 );
buf ( n17169 , n5912 );
buf ( n17170 , n17169 );
not ( n17171 , n17170 );
buf ( n17172 , n5913 );
not ( n17173 , n17172 );
not ( n17174 , n17173 );
or ( n17175 , n17171 , n17174 );
not ( n17176 , n17169 );
buf ( n17177 , n17172 );
nand ( n17178 , n17176 , n17177 );
nand ( n17179 , n17175 , n17178 );
buf ( n17180 , n5914 );
buf ( n17181 , n17180 );
and ( n17182 , n17179 , n17181 );
not ( n17183 , n17179 );
not ( n17184 , n17180 );
and ( n17185 , n17183 , n17184 );
nor ( n17186 , n17182 , n17185 );
not ( n17187 , n17186 );
and ( n17188 , n17168 , n17187 );
not ( n17189 , n17168 );
and ( n17190 , n17189 , n17186 );
nor ( n17191 , n17188 , n17190 );
buf ( n17192 , n17191 );
not ( n17193 , n17192 );
or ( n17194 , n17145 , n17193 );
not ( n17195 , n16589 );
buf ( n17196 , n17154 );
xor ( n17197 , n17186 , n17196 );
buf ( n17198 , n17164 );
xnor ( n17199 , n17197 , n17198 );
buf ( n17200 , n17199 );
nand ( n17201 , n17195 , n17200 );
nand ( n17202 , n17194 , n17201 );
buf ( n17203 , n7105 );
and ( n17204 , n17202 , n17203 );
not ( n17205 , n17202 );
xor ( n17206 , n7081 , n7103 );
buf ( n17207 , n7091 );
xnor ( n17208 , n17206 , n17207 );
buf ( n17209 , n17208 );
and ( n17210 , n17205 , n17209 );
nor ( n17211 , n17204 , n17210 );
not ( n17212 , n17211 );
not ( n17213 , n16851 );
nand ( n17214 , n17213 , n16854 );
not ( n17215 , n17214 );
or ( n17216 , n17212 , n17215 );
or ( n17217 , n17211 , n17214 );
nand ( n17218 , n17216 , n17217 );
not ( n17219 , n15302 );
not ( n17220 , n13857 );
or ( n17221 , n17219 , n17220 );
or ( n17222 , n13857 , n15302 );
nand ( n17223 , n17221 , n17222 );
not ( n17224 , n12863 );
not ( n17225 , n12843 );
and ( n17226 , n17224 , n17225 );
and ( n17227 , n12863 , n12843 );
nor ( n17228 , n17226 , n17227 );
buf ( n17229 , n17228 );
and ( n17230 , n17223 , n17229 );
not ( n17231 , n17223 );
not ( n17232 , n17229 );
and ( n17233 , n17231 , n17232 );
nor ( n17234 , n17230 , n17233 );
nand ( n17235 , n17234 , n9787 );
not ( n17236 , n17235 );
buf ( n17237 , n15188 );
not ( n17238 , n17237 );
buf ( n17239 , n16674 );
not ( n17240 , n17239 );
or ( n17241 , n17238 , n17240 );
or ( n17242 , n17239 , n17237 );
nand ( n17243 , n17241 , n17242 );
and ( n17244 , n17243 , n16719 );
not ( n17245 , n17243 );
not ( n17246 , n16718 );
buf ( n17247 , n17246 );
and ( n17248 , n17245 , n17247 );
nor ( n17249 , n17244 , n17248 );
not ( n17250 , n17249 );
and ( n17251 , n17236 , n17250 );
and ( n17252 , n17235 , n17249 );
nor ( n17253 , n17251 , n17252 );
and ( n17254 , n17218 , n17253 );
not ( n17255 , n17218 );
not ( n17256 , n17253 );
and ( n17257 , n17255 , n17256 );
nor ( n17258 , n17254 , n17257 );
not ( n17259 , n17258 );
not ( n17260 , n17259 );
and ( n17261 , n17144 , n17260 );
and ( n17262 , n17259 , n17143 );
nor ( n17263 , n17261 , n17262 );
not ( n17264 , n17263 );
or ( n17265 , n16860 , n17264 );
not ( n17266 , n16859 );
not ( n17267 , n17259 );
not ( n17268 , n17143 );
or ( n17269 , n17267 , n17268 );
not ( n17270 , n17143 );
nand ( n17271 , n17270 , n17258 );
nand ( n17272 , n17269 , n17271 );
nand ( n17273 , n17266 , n17272 );
nand ( n17274 , n17265 , n17273 );
not ( n17275 , n13696 );
not ( n17276 , n16844 );
or ( n17277 , n17275 , n17276 );
or ( n17278 , n16844 , n13696 );
nand ( n17279 , n17277 , n17278 );
not ( n17280 , n17279 );
not ( n17281 , n17280 );
not ( n17282 , n16212 );
or ( n17283 , n17281 , n17282 );
nand ( n17284 , n12525 , n17279 );
nand ( n17285 , n17283 , n17284 );
not ( n17286 , n17285 );
nand ( n17287 , n17286 , n11289 );
not ( n17288 , n17287 );
not ( n17289 , n15793 );
buf ( n17290 , n9341 );
not ( n17291 , n17290 );
not ( n17292 , n15830 );
or ( n17293 , n17291 , n17292 );
or ( n17294 , n15830 , n17290 );
nand ( n17295 , n17293 , n17294 );
not ( n17296 , n17295 );
and ( n17297 , n17289 , n17296 );
and ( n17298 , n15843 , n17295 );
nor ( n17299 , n17297 , n17298 );
not ( n17300 , n17299 );
not ( n17301 , n17300 );
and ( n17302 , n17288 , n17301 );
and ( n17303 , n17287 , n17300 );
nor ( n17304 , n17302 , n17303 );
not ( n17305 , n17304 );
not ( n17306 , n17126 );
buf ( n17307 , n8014 );
not ( n17308 , n17307 );
not ( n17309 , n17109 );
not ( n17310 , n17309 );
or ( n17311 , n17308 , n17310 );
or ( n17312 , n17309 , n17307 );
nand ( n17313 , n17311 , n17312 );
not ( n17314 , n17313 );
and ( n17315 , n17306 , n17314 );
and ( n17316 , n17126 , n17313 );
nor ( n17317 , n17315 , n17316 );
not ( n17318 , n7704 );
buf ( n17319 , n5915 );
buf ( n17320 , n17319 );
not ( n17321 , n17320 );
buf ( n17322 , n5916 );
not ( n17323 , n17322 );
not ( n17324 , n17323 );
or ( n17325 , n17321 , n17324 );
not ( n17326 , n17319 );
buf ( n17327 , n17322 );
nand ( n17328 , n17326 , n17327 );
nand ( n17329 , n17325 , n17328 );
buf ( n17330 , n5917 );
buf ( n17331 , n17330 );
and ( n17332 , n17329 , n17331 );
not ( n17333 , n17329 );
not ( n17334 , n17330 );
and ( n17335 , n17333 , n17334 );
nor ( n17336 , n17332 , n17335 );
buf ( n17337 , n5918 );
nand ( n17338 , n6905 , n17337 );
buf ( n17339 , n5919 );
buf ( n17340 , n17339 );
and ( n17341 , n17338 , n17340 );
not ( n17342 , n17338 );
not ( n17343 , n17339 );
and ( n17344 , n17342 , n17343 );
nor ( n17345 , n17341 , n17344 );
xor ( n17346 , n17336 , n17345 );
buf ( n17347 , n5920 );
nand ( n17348 , n7471 , n17347 );
buf ( n17349 , n5921 );
buf ( n17350 , n17349 );
and ( n17351 , n17348 , n17350 );
not ( n17352 , n17348 );
not ( n17353 , n17349 );
and ( n17354 , n17352 , n17353 );
nor ( n17355 , n17351 , n17354 );
not ( n17356 , n17355 );
xnor ( n17357 , n17346 , n17356 );
not ( n17358 , n17357 );
or ( n17359 , n17318 , n17358 );
or ( n17360 , n17357 , n7704 );
nand ( n17361 , n17359 , n17360 );
not ( n17362 , n17361 );
not ( n17363 , n16674 );
not ( n17364 , n17363 );
not ( n17365 , n17364 );
and ( n17366 , n17362 , n17365 );
and ( n17367 , n17361 , n17364 );
nor ( n17368 , n17366 , n17367 );
nand ( n17369 , n11134 , n17368 );
xor ( n17370 , n17317 , n17369 );
not ( n17371 , n17370 );
or ( n17372 , n17305 , n17371 );
or ( n17373 , n17370 , n17304 );
nand ( n17374 , n17372 , n17373 );
buf ( n17375 , n15500 );
xor ( n17376 , n17375 , n7312 );
xnor ( n17377 , n17376 , n7336 );
not ( n17378 , n17377 );
nand ( n17379 , n17378 , n10948 );
buf ( n17380 , n5922 );
not ( n17381 , n17380 );
buf ( n17382 , n5923 );
nand ( n17383 , n6817 , n17382 );
buf ( n17384 , n17383 );
not ( n17385 , n17384 );
or ( n17386 , n17381 , n17385 );
or ( n17387 , n17384 , n17380 );
nand ( n17388 , n17386 , n17387 );
not ( n17389 , n17388 );
buf ( n17390 , n14463 );
not ( n17391 , n17390 );
or ( n17392 , n17389 , n17391 );
not ( n17393 , n17388 );
nand ( n17394 , n17393 , n14464 );
nand ( n17395 , n17392 , n17394 );
buf ( n17396 , n14430 );
not ( n17397 , n17396 );
and ( n17398 , n17395 , n17397 );
not ( n17399 , n17395 );
and ( n17400 , n17399 , n17396 );
nor ( n17401 , n17398 , n17400 );
buf ( n17402 , n17401 );
not ( n17403 , n17402 );
and ( n17404 , n17379 , n17403 );
not ( n17405 , n17379 );
and ( n17406 , n17405 , n17402 );
nor ( n17407 , n17404 , n17406 );
and ( n17408 , n17374 , n17407 );
not ( n17409 , n17374 );
not ( n17410 , n17407 );
and ( n17411 , n17409 , n17410 );
nor ( n17412 , n17408 , n17411 );
not ( n17413 , n17412 );
not ( n17414 , n17413 );
buf ( n17415 , n5924 );
not ( n17416 , n17050 );
not ( n17417 , n7888 );
not ( n17418 , n17417 );
or ( n17419 , n17416 , n17418 );
not ( n17420 , n17049 );
nand ( n17421 , n17420 , n7889 );
nand ( n17422 , n17419 , n17421 );
buf ( n17423 , n5925 );
buf ( n17424 , n17423 );
and ( n17425 , n17422 , n17424 );
not ( n17426 , n17422 );
not ( n17427 , n17423 );
and ( n17428 , n17426 , n17427 );
nor ( n17429 , n17425 , n17428 );
xor ( n17430 , n17429 , n16042 );
buf ( n17431 , n5926 );
nand ( n17432 , n6934 , n17431 );
buf ( n17433 , n5927 );
buf ( n17434 , n17433 );
and ( n17435 , n17432 , n17434 );
not ( n17436 , n17432 );
not ( n17437 , n17433 );
and ( n17438 , n17436 , n17437 );
nor ( n17439 , n17435 , n17438 );
not ( n17440 , n17439 );
xnor ( n17441 , n17430 , n17440 );
xor ( n17442 , n17415 , n17441 );
buf ( n17443 , n5928 );
buf ( n17444 , n17443 );
not ( n17445 , n17444 );
buf ( n17446 , n5929 );
not ( n17447 , n17446 );
not ( n17448 , n17447 );
or ( n17449 , n17445 , n17448 );
not ( n17450 , n17443 );
buf ( n17451 , n17446 );
nand ( n17452 , n17450 , n17451 );
nand ( n17453 , n17449 , n17452 );
buf ( n17454 , n5930 );
buf ( n17455 , n17454 );
and ( n17456 , n17453 , n17455 );
not ( n17457 , n17453 );
not ( n17458 , n17454 );
and ( n17459 , n17457 , n17458 );
nor ( n17460 , n17456 , n17459 );
buf ( n17461 , n5931 );
nand ( n17462 , n6706 , n17461 );
buf ( n17463 , n5932 );
buf ( n17464 , n17463 );
and ( n17465 , n17462 , n17464 );
not ( n17466 , n17462 );
not ( n17467 , n17463 );
and ( n17468 , n17466 , n17467 );
nor ( n17469 , n17465 , n17468 );
xor ( n17470 , n17460 , n17469 );
buf ( n17471 , n5933 );
nand ( n17472 , n7617 , n17471 );
buf ( n17473 , n5934 );
buf ( n17474 , n17473 );
and ( n17475 , n17472 , n17474 );
not ( n17476 , n17472 );
not ( n17477 , n17473 );
and ( n17478 , n17476 , n17477 );
nor ( n17479 , n17475 , n17478 );
xnor ( n17480 , n17470 , n17479 );
not ( n17481 , n17480 );
xnor ( n17482 , n17442 , n17481 );
not ( n17483 , n17482 );
not ( n17484 , n17483 );
nand ( n17485 , n17484 , n11368 );
not ( n17486 , n17485 );
buf ( n17487 , n5935 );
nand ( n17488 , n12401 , n17487 );
buf ( n17489 , n5936 );
buf ( n17490 , n17489 );
and ( n17491 , n17488 , n17490 );
not ( n17492 , n17488 );
not ( n17493 , n17489 );
and ( n17494 , n17492 , n17493 );
nor ( n17495 , n17491 , n17494 );
not ( n17496 , n17495 );
buf ( n17497 , n5937 );
buf ( n17498 , n17497 );
not ( n17499 , n17498 );
buf ( n17500 , n5938 );
not ( n17501 , n17500 );
not ( n17502 , n17501 );
or ( n17503 , n17499 , n17502 );
not ( n17504 , n17497 );
buf ( n17505 , n17500 );
nand ( n17506 , n17504 , n17505 );
nand ( n17507 , n17503 , n17506 );
buf ( n17508 , n5939 );
not ( n17509 , n17508 );
and ( n17510 , n17507 , n17509 );
not ( n17511 , n17507 );
buf ( n17512 , n17508 );
and ( n17513 , n17511 , n17512 );
nor ( n17514 , n17510 , n17513 );
buf ( n17515 , n5940 );
nand ( n17516 , n7133 , n17515 );
buf ( n17517 , n5941 );
buf ( n17518 , n17517 );
and ( n17519 , n17516 , n17518 );
not ( n17520 , n17516 );
not ( n17521 , n17517 );
and ( n17522 , n17520 , n17521 );
nor ( n17523 , n17519 , n17522 );
xor ( n17524 , n17514 , n17523 );
buf ( n17525 , n5942 );
nand ( n17526 , n6985 , n17525 );
buf ( n17527 , n5943 );
buf ( n17528 , n17527 );
and ( n17529 , n17526 , n17528 );
not ( n17530 , n17526 );
not ( n17531 , n17527 );
and ( n17532 , n17530 , n17531 );
nor ( n17533 , n17529 , n17532 );
xor ( n17534 , n17524 , n17533 );
not ( n17535 , n17534 );
not ( n17536 , n17535 );
or ( n17537 , n17496 , n17536 );
or ( n17538 , n17535 , n17495 );
nand ( n17539 , n17537 , n17538 );
not ( n17540 , n17539 );
xor ( n17541 , n14225 , n14234 );
xnor ( n17542 , n17541 , n14241 );
not ( n17543 , n17542 );
not ( n17544 , n17543 );
or ( n17545 , n17540 , n17544 );
or ( n17546 , n14243 , n17539 );
nand ( n17547 , n17545 , n17546 );
buf ( n17548 , n17547 );
not ( n17549 , n17548 );
and ( n17550 , n17486 , n17549 );
and ( n17551 , n17485 , n17548 );
nor ( n17552 , n17550 , n17551 );
not ( n17553 , n17552 );
buf ( n17554 , n9774 );
not ( n17555 , n17554 );
buf ( n17556 , n5944 );
not ( n17557 , n17556 );
buf ( n17558 , n5945 );
buf ( n17559 , n17558 );
not ( n17560 , n17559 );
buf ( n17561 , n5946 );
not ( n17562 , n17561 );
not ( n17563 , n17562 );
or ( n17564 , n17560 , n17563 );
not ( n17565 , n17558 );
buf ( n17566 , n17561 );
nand ( n17567 , n17565 , n17566 );
nand ( n17568 , n17564 , n17567 );
xor ( n17569 , n17557 , n17568 );
buf ( n17570 , n5947 );
buf ( n17571 , n5948 );
xor ( n17572 , n17570 , n17571 );
buf ( n17573 , n5949 );
nand ( n17574 , n8785 , n17573 );
xnor ( n17575 , n17572 , n17574 );
xor ( n17576 , n17569 , n17575 );
not ( n17577 , n17576 );
not ( n17578 , n17577 );
or ( n17579 , n17555 , n17578 );
or ( n17580 , n17577 , n17554 );
nand ( n17581 , n17579 , n17580 );
buf ( n17582 , n8026 );
not ( n17583 , n17582 );
and ( n17584 , n17581 , n17583 );
not ( n17585 , n17581 );
and ( n17586 , n17585 , n17582 );
nor ( n17587 , n17584 , n17586 );
not ( n17588 , n17587 );
not ( n17589 , n15371 );
not ( n17590 , n12404 );
not ( n17591 , n16948 );
not ( n17592 , n17591 );
not ( n17593 , n17592 );
or ( n17594 , n17590 , n17593 );
not ( n17595 , n12404 );
nand ( n17596 , n17591 , n17595 );
nand ( n17597 , n17594 , n17596 );
not ( n17598 , n17597 );
or ( n17599 , n17589 , n17598 );
or ( n17600 , n17597 , n16955 );
nand ( n17601 , n17599 , n17600 );
not ( n17602 , n17601 );
nand ( n17603 , n17602 , n11723 );
not ( n17604 , n17603 );
or ( n17605 , n17588 , n17604 );
or ( n17606 , n17603 , n17587 );
nand ( n17607 , n17605 , n17606 );
not ( n17608 , n17607 );
and ( n17609 , n17553 , n17608 );
and ( n17610 , n17552 , n17607 );
nor ( n17611 , n17609 , n17610 );
not ( n17612 , n17611 );
not ( n17613 , n17612 );
and ( n17614 , n17414 , n17613 );
and ( n17615 , n17413 , n17612 );
nor ( n17616 , n17614 , n17615 );
buf ( n17617 , n17616 );
and ( n17618 , n17274 , n17617 );
not ( n17619 , n17274 );
not ( n17620 , n17611 );
not ( n17621 , n17412 );
or ( n17622 , n17620 , n17621 );
not ( n17623 , n17611 );
nand ( n17624 , n17623 , n17413 );
nand ( n17625 , n17622 , n17624 );
buf ( n17626 , n17625 );
and ( n17627 , n17619 , n17626 );
nor ( n17628 , n17618 , n17627 );
buf ( n17629 , n5950 );
buf ( n17630 , n17629 );
not ( n17631 , n17630 );
buf ( n17632 , n5951 );
not ( n17633 , n17632 );
not ( n17634 , n17633 );
or ( n17635 , n17631 , n17634 );
not ( n17636 , n17629 );
buf ( n17637 , n17632 );
nand ( n17638 , n17636 , n17637 );
nand ( n17639 , n17635 , n17638 );
buf ( n17640 , n5952 );
buf ( n17641 , n17640 );
and ( n17642 , n17639 , n17641 );
not ( n17643 , n17639 );
not ( n17644 , n17640 );
and ( n17645 , n17643 , n17644 );
nor ( n17646 , n17642 , n17645 );
buf ( n17647 , n5953 );
nand ( n17648 , n7865 , n17647 );
buf ( n17649 , n5954 );
buf ( n17650 , n17649 );
and ( n17651 , n17648 , n17650 );
not ( n17652 , n17648 );
not ( n17653 , n17649 );
and ( n17654 , n17652 , n17653 );
nor ( n17655 , n17651 , n17654 );
xor ( n17656 , n17646 , n17655 );
buf ( n17657 , n5955 );
nand ( n17658 , n6706 , n17657 );
buf ( n17659 , n5956 );
buf ( n17660 , n17659 );
and ( n17661 , n17658 , n17660 );
not ( n17662 , n17658 );
not ( n17663 , n17659 );
and ( n17664 , n17662 , n17663 );
nor ( n17665 , n17661 , n17664 );
xnor ( n17666 , n17656 , n17665 );
not ( n17667 , n17666 );
and ( n17668 , n15574 , n17667 );
not ( n17669 , n15574 );
and ( n17670 , n17669 , n17666 );
or ( n17671 , n17668 , n17670 );
not ( n17672 , n13617 );
buf ( n17673 , n17672 );
and ( n17674 , n17671 , n17673 );
not ( n17675 , n17671 );
and ( n17676 , n17675 , n13618 );
nor ( n17677 , n17674 , n17676 );
buf ( n17678 , n5957 );
nand ( n17679 , n7921 , n17678 );
buf ( n17680 , n5958 );
not ( n17681 , n17680 );
and ( n17682 , n17679 , n17681 );
not ( n17683 , n17679 );
buf ( n17684 , n17680 );
and ( n17685 , n17683 , n17684 );
nor ( n17686 , n17682 , n17685 );
not ( n17687 , n17686 );
and ( n17688 , n17687 , n13319 );
not ( n17689 , n17687 );
not ( n17690 , n13298 );
xor ( n17691 , n17690 , n13317 );
xnor ( n17692 , n17691 , n13307 );
not ( n17693 , n17692 );
and ( n17694 , n17689 , n17693 );
nor ( n17695 , n17688 , n17694 );
and ( n17696 , n17695 , n13343 );
not ( n17697 , n17695 );
buf ( n17698 , n13342 );
and ( n17699 , n17697 , n17698 );
or ( n17700 , n17696 , n17699 );
nand ( n17701 , n17677 , n17700 );
not ( n17702 , n17701 );
buf ( n17703 , n5959 );
nand ( n17704 , n7230 , n17703 );
buf ( n17705 , n5960 );
not ( n17706 , n17705 );
and ( n17707 , n17704 , n17706 );
not ( n17708 , n17704 );
buf ( n17709 , n17705 );
and ( n17710 , n17708 , n17709 );
nor ( n17711 , n17707 , n17710 );
buf ( n17712 , n17711 );
not ( n17713 , n17712 );
not ( n17714 , n14641 );
or ( n17715 , n17713 , n17714 );
not ( n17716 , n17712 );
not ( n17717 , n14641 );
nand ( n17718 , n17716 , n17717 );
nand ( n17719 , n17715 , n17718 );
and ( n17720 , n17719 , n11009 );
not ( n17721 , n17719 );
and ( n17722 , n17721 , n10995 );
nor ( n17723 , n17720 , n17722 );
not ( n17724 , n17723 );
and ( n17725 , n17702 , n17724 );
and ( n17726 , n17701 , n17723 );
nor ( n17727 , n17725 , n17726 );
not ( n17728 , n17727 );
not ( n17729 , n17728 );
not ( n17730 , n12220 );
xor ( n17731 , n17730 , n12228 );
xnor ( n17732 , n17731 , n12235 );
not ( n17733 , n17732 );
not ( n17734 , n15548 );
not ( n17735 , n11991 );
and ( n17736 , n17734 , n17735 );
and ( n17737 , n15548 , n11991 );
nor ( n17738 , n17736 , n17737 );
not ( n17739 , n17738 );
not ( n17740 , n17739 );
or ( n17741 , n17733 , n17740 );
not ( n17742 , n17732 );
nand ( n17743 , n17742 , n17738 );
nand ( n17744 , n17741 , n17743 );
not ( n17745 , n17744 );
not ( n17746 , n14236 );
buf ( n17747 , n5961 );
buf ( n17748 , n17747 );
not ( n17749 , n17748 );
buf ( n17750 , n5962 );
not ( n17751 , n17750 );
not ( n17752 , n17751 );
or ( n17753 , n17749 , n17752 );
not ( n17754 , n17747 );
buf ( n17755 , n17750 );
nand ( n17756 , n17754 , n17755 );
nand ( n17757 , n17753 , n17756 );
buf ( n17758 , n5963 );
not ( n17759 , n17758 );
and ( n17760 , n17757 , n17759 );
not ( n17761 , n17757 );
buf ( n17762 , n17758 );
and ( n17763 , n17761 , n17762 );
nor ( n17764 , n17760 , n17763 );
xor ( n17765 , n17764 , n12029 );
buf ( n17766 , n5964 );
nand ( n17767 , n7785 , n17766 );
buf ( n17768 , n5965 );
buf ( n17769 , n17768 );
and ( n17770 , n17767 , n17769 );
not ( n17771 , n17767 );
not ( n17772 , n17768 );
and ( n17773 , n17771 , n17772 );
nor ( n17774 , n17770 , n17773 );
xnor ( n17775 , n17765 , n17774 );
not ( n17776 , n17775 );
not ( n17777 , n17776 );
or ( n17778 , n17746 , n17777 );
not ( n17779 , n14236 );
not ( n17780 , n17775 );
not ( n17781 , n17780 );
nand ( n17782 , n17779 , n17781 );
nand ( n17783 , n17778 , n17782 );
buf ( n17784 , n5966 );
buf ( n17785 , n17784 );
not ( n17786 , n17785 );
buf ( n17787 , n5967 );
not ( n17788 , n17787 );
not ( n17789 , n17788 );
or ( n17790 , n17786 , n17789 );
not ( n17791 , n17784 );
buf ( n17792 , n17787 );
nand ( n17793 , n17791 , n17792 );
nand ( n17794 , n17790 , n17793 );
buf ( n17795 , n5968 );
not ( n17796 , n17795 );
and ( n17797 , n17794 , n17796 );
not ( n17798 , n17794 );
buf ( n17799 , n17795 );
and ( n17800 , n17798 , n17799 );
nor ( n17801 , n17797 , n17800 );
buf ( n17802 , n5969 );
nand ( n17803 , n6706 , n17802 );
buf ( n17804 , n5970 );
buf ( n17805 , n17804 );
and ( n17806 , n17803 , n17805 );
not ( n17807 , n17803 );
not ( n17808 , n17804 );
and ( n17809 , n17807 , n17808 );
nor ( n17810 , n17806 , n17809 );
xor ( n17811 , n17801 , n17810 );
buf ( n17812 , n5971 );
nand ( n17813 , n10107 , n17812 );
buf ( n17814 , n5972 );
buf ( n17815 , n17814 );
and ( n17816 , n17813 , n17815 );
not ( n17817 , n17813 );
not ( n17818 , n17814 );
and ( n17819 , n17817 , n17818 );
nor ( n17820 , n17816 , n17819 );
not ( n17821 , n17820 );
xnor ( n17822 , n17811 , n17821 );
buf ( n17823 , n17822 );
not ( n17824 , n17823 );
and ( n17825 , n17783 , n17824 );
not ( n17826 , n17783 );
not ( n17827 , n17822 );
not ( n17828 , n17827 );
and ( n17829 , n17826 , n17828 );
nor ( n17830 , n17825 , n17829 );
nand ( n17831 , n17745 , n17830 );
not ( n17832 , n17831 );
not ( n17833 , n7693 );
not ( n17834 , n17336 );
xor ( n17835 , n17834 , n17355 );
not ( n17836 , n17345 );
xnor ( n17837 , n17835 , n17836 );
not ( n17838 , n17837 );
or ( n17839 , n17833 , n17838 );
or ( n17840 , n17837 , n7693 );
nand ( n17841 , n17839 , n17840 );
and ( n17842 , n17841 , n17239 );
not ( n17843 , n17841 );
and ( n17844 , n17843 , n17363 );
nor ( n17845 , n17842 , n17844 );
not ( n17846 , n17845 );
not ( n17847 , n17846 );
and ( n17848 , n17832 , n17847 );
and ( n17849 , n17831 , n17846 );
nor ( n17850 , n17848 , n17849 );
not ( n17851 , n17850 );
buf ( n17852 , n10006 );
not ( n17853 , n17852 );
buf ( n17854 , n5973 );
not ( n17855 , n17854 );
buf ( n17856 , n5974 );
buf ( n17857 , n17856 );
and ( n17858 , n17855 , n17857 );
not ( n17859 , n17855 );
not ( n17860 , n17856 );
and ( n17861 , n17859 , n17860 );
nor ( n17862 , n17858 , n17861 );
xor ( n17863 , n6686 , n17862 );
buf ( n17864 , n5975 );
xor ( n17865 , n14915 , n17864 );
buf ( n17866 , n5976 );
nand ( n17867 , n7134 , n17866 );
xnor ( n17868 , n17865 , n17867 );
xnor ( n17869 , n17863 , n17868 );
not ( n17870 , n17869 );
or ( n17871 , n17853 , n17870 );
xor ( n17872 , n6686 , n17862 );
xnor ( n17873 , n17872 , n17868 );
or ( n17874 , n17873 , n17852 );
nand ( n17875 , n17871 , n17874 );
and ( n17876 , n17875 , n7584 );
not ( n17877 , n17875 );
and ( n17878 , n17877 , n7580 );
nor ( n17879 , n17876 , n17878 );
not ( n17880 , n17879 );
xor ( n17881 , n9577 , n9596 );
not ( n17882 , n9586 );
xnor ( n17883 , n17881 , n17882 );
buf ( n17884 , n17883 );
not ( n17885 , n17884 );
buf ( n17886 , n5977 );
nand ( n17887 , n7750 , n17886 );
buf ( n17888 , n5978 );
buf ( n17889 , n17888 );
and ( n17890 , n17887 , n17889 );
not ( n17891 , n17887 );
not ( n17892 , n17888 );
and ( n17893 , n17891 , n17892 );
nor ( n17894 , n17890 , n17893 );
buf ( n17895 , n17894 );
not ( n17896 , n17895 );
not ( n17897 , n12364 );
not ( n17898 , n17897 );
or ( n17899 , n17896 , n17898 );
not ( n17900 , n12364 );
or ( n17901 , n17900 , n17895 );
nand ( n17902 , n17899 , n17901 );
not ( n17903 , n17902 );
or ( n17904 , n17885 , n17903 );
or ( n17905 , n17902 , n17884 );
nand ( n17906 , n17904 , n17905 );
nand ( n17907 , n17880 , n17906 );
buf ( n17908 , n5979 );
not ( n17909 , n17908 );
not ( n17910 , n17909 );
not ( n17911 , n9031 );
or ( n17912 , n17910 , n17911 );
xor ( n17913 , n9011 , n9020 );
xnor ( n17914 , n17913 , n9030 );
or ( n17915 , n17909 , n17914 );
nand ( n17916 , n17912 , n17915 );
not ( n17917 , n9074 );
buf ( n17918 , n17917 );
and ( n17919 , n17916 , n17918 );
not ( n17920 , n17916 );
and ( n17921 , n17920 , n9075 );
nor ( n17922 , n17919 , n17921 );
and ( n17923 , n17907 , n17922 );
not ( n17924 , n17907 );
not ( n17925 , n17922 );
and ( n17926 , n17924 , n17925 );
nor ( n17927 , n17923 , n17926 );
not ( n17928 , n17927 );
or ( n17929 , n17851 , n17928 );
or ( n17930 , n17927 , n17850 );
nand ( n17931 , n17929 , n17930 );
not ( n17932 , n17723 );
not ( n17933 , n17700 );
nand ( n17934 , n17932 , n17933 );
not ( n17935 , n9098 );
not ( n17936 , n8536 );
or ( n17937 , n17935 , n17936 );
not ( n17938 , n8531 );
or ( n17939 , n17938 , n9098 );
nand ( n17940 , n17937 , n17939 );
buf ( n17941 , n5980 );
buf ( n17942 , n17941 );
not ( n17943 , n17942 );
buf ( n17944 , n5981 );
not ( n17945 , n17944 );
not ( n17946 , n17945 );
or ( n17947 , n17943 , n17946 );
not ( n17948 , n17941 );
buf ( n17949 , n17944 );
nand ( n17950 , n17948 , n17949 );
nand ( n17951 , n17947 , n17950 );
buf ( n17952 , n5982 );
buf ( n17953 , n17952 );
and ( n17954 , n17951 , n17953 );
not ( n17955 , n17951 );
not ( n17956 , n17952 );
and ( n17957 , n17955 , n17956 );
nor ( n17958 , n17954 , n17957 );
buf ( n17959 , n5983 );
nand ( n17960 , n6760 , n17959 );
buf ( n17961 , n5984 );
not ( n17962 , n17961 );
and ( n17963 , n17960 , n17962 );
not ( n17964 , n17960 );
buf ( n17965 , n17961 );
and ( n17966 , n17964 , n17965 );
nor ( n17967 , n17963 , n17966 );
xor ( n17968 , n17958 , n17967 );
buf ( n17969 , n5985 );
nand ( n17970 , n6804 , n17969 );
buf ( n17971 , n5986 );
buf ( n17972 , n17971 );
and ( n17973 , n17970 , n17972 );
not ( n17974 , n17970 );
not ( n17975 , n17971 );
and ( n17976 , n17974 , n17975 );
nor ( n17977 , n17973 , n17976 );
xor ( n17978 , n17968 , n17977 );
not ( n17979 , n17978 );
not ( n17980 , n17979 );
and ( n17981 , n17940 , n17980 );
not ( n17982 , n17940 );
not ( n17983 , n17980 );
and ( n17984 , n17982 , n17983 );
nor ( n17985 , n17981 , n17984 );
and ( n17986 , n17934 , n17985 );
not ( n17987 , n17934 );
not ( n17988 , n17985 );
and ( n17989 , n17987 , n17988 );
nor ( n17990 , n17986 , n17989 );
xnor ( n17991 , n17931 , n17990 );
buf ( n17992 , n7576 );
not ( n17993 , n17992 );
not ( n17994 , n6772 );
or ( n17995 , n17993 , n17994 );
not ( n17996 , n17992 );
not ( n17997 , n6771 );
nand ( n17998 , n17996 , n17997 );
nand ( n17999 , n17995 , n17998 );
not ( n18000 , n10941 );
and ( n18001 , n17999 , n18000 );
not ( n18002 , n17999 );
and ( n18003 , n18002 , n10942 );
nor ( n18004 , n18001 , n18003 );
buf ( n18005 , n5987 );
nand ( n18006 , n6607 , n18005 );
buf ( n18007 , n5988 );
buf ( n18008 , n18007 );
and ( n18009 , n18006 , n18008 );
not ( n18010 , n18006 );
not ( n18011 , n18007 );
and ( n18012 , n18010 , n18011 );
nor ( n18013 , n18009 , n18012 );
buf ( n18014 , n18013 );
not ( n18015 , n18014 );
not ( n18016 , n9220 );
or ( n18017 , n18015 , n18016 );
not ( n18018 , n10854 );
or ( n18019 , n18018 , n18014 );
nand ( n18020 , n18017 , n18019 );
not ( n18021 , n15287 );
and ( n18022 , n18020 , n18021 );
not ( n18023 , n18020 );
not ( n18024 , n10896 );
and ( n18025 , n18023 , n18024 );
nor ( n18026 , n18022 , n18025 );
not ( n18027 , n18026 );
nand ( n18028 , n18004 , n18027 );
not ( n18029 , n18028 );
buf ( n18030 , n5989 );
buf ( n18031 , n18030 );
not ( n18032 , n18031 );
buf ( n18033 , n5990 );
not ( n18034 , n18033 );
not ( n18035 , n18034 );
or ( n18036 , n18032 , n18035 );
not ( n18037 , n18030 );
buf ( n18038 , n18033 );
nand ( n18039 , n18037 , n18038 );
nand ( n18040 , n18036 , n18039 );
buf ( n18041 , n5991 );
not ( n18042 , n18041 );
and ( n18043 , n18040 , n18042 );
not ( n18044 , n18040 );
buf ( n18045 , n18041 );
and ( n18046 , n18044 , n18045 );
nor ( n18047 , n18043 , n18046 );
buf ( n18048 , n5992 );
nand ( n18049 , n7471 , n18048 );
buf ( n18050 , n5993 );
buf ( n18051 , n18050 );
and ( n18052 , n18049 , n18051 );
not ( n18053 , n18049 );
not ( n18054 , n18050 );
and ( n18055 , n18053 , n18054 );
nor ( n18056 , n18052 , n18055 );
xor ( n18057 , n18047 , n18056 );
buf ( n18058 , n5994 );
nand ( n18059 , n7196 , n18058 );
buf ( n18060 , n5995 );
not ( n18061 , n18060 );
and ( n18062 , n18059 , n18061 );
not ( n18063 , n18059 );
buf ( n18064 , n18060 );
and ( n18065 , n18063 , n18064 );
nor ( n18066 , n18062 , n18065 );
xnor ( n18067 , n18057 , n18066 );
buf ( n18068 , n18067 );
xor ( n18069 , n10158 , n18068 );
buf ( n18070 , n5996 );
not ( n18071 , n18070 );
buf ( n18072 , n5997 );
not ( n18073 , n18072 );
buf ( n18074 , n14432 );
and ( n18075 , n18073 , n18074 );
not ( n18076 , n18073 );
and ( n18077 , n18076 , n14433 );
nor ( n18078 , n18075 , n18077 );
xor ( n18079 , n18071 , n18078 );
buf ( n18080 , n5998 );
xor ( n18081 , n18080 , n17380 );
xnor ( n18082 , n18081 , n17383 );
xnor ( n18083 , n18079 , n18082 );
buf ( n18084 , n18083 );
xnor ( n18085 , n18069 , n18084 );
not ( n18086 , n18085 );
not ( n18087 , n18086 );
or ( n18088 , n18029 , n18087 );
or ( n18089 , n18086 , n18028 );
nand ( n18090 , n18088 , n18089 );
not ( n18091 , n18090 );
not ( n18092 , n18091 );
not ( n18093 , n14520 );
not ( n18094 , n11413 );
not ( n18095 , n18094 );
not ( n18096 , n18095 );
and ( n18097 , n18093 , n18096 );
and ( n18098 , n14521 , n18095 );
nor ( n18099 , n18097 , n18098 );
buf ( n18100 , n5999 );
buf ( n18101 , n18100 );
not ( n18102 , n18101 );
buf ( n18103 , n6000 );
not ( n18104 , n18103 );
not ( n18105 , n18104 );
or ( n18106 , n18102 , n18105 );
not ( n18107 , n18100 );
buf ( n18108 , n18103 );
nand ( n18109 , n18107 , n18108 );
nand ( n18110 , n18106 , n18109 );
not ( n18111 , n18110 );
buf ( n18112 , n6001 );
buf ( n18113 , n6002 );
nand ( n18114 , n7477 , n18113 );
buf ( n18115 , n6003 );
buf ( n18116 , n18115 );
and ( n18117 , n18114 , n18116 );
not ( n18118 , n18114 );
not ( n18119 , n18115 );
and ( n18120 , n18118 , n18119 );
nor ( n18121 , n18117 , n18120 );
xor ( n18122 , n18112 , n18121 );
buf ( n18123 , n6004 );
nand ( n18124 , n7082 , n18123 );
buf ( n18125 , n6005 );
not ( n18126 , n18125 );
and ( n18127 , n18124 , n18126 );
not ( n18128 , n18124 );
buf ( n18129 , n18125 );
and ( n18130 , n18128 , n18129 );
nor ( n18131 , n18127 , n18130 );
xnor ( n18132 , n18122 , n18131 );
not ( n18133 , n18132 );
not ( n18134 , n18133 );
or ( n18135 , n18111 , n18134 );
not ( n18136 , n18110 );
nand ( n18137 , n18132 , n18136 );
nand ( n18138 , n18135 , n18137 );
not ( n18139 , n18138 );
and ( n18140 , n18099 , n18139 );
not ( n18141 , n18099 );
and ( n18142 , n18141 , n18138 );
nor ( n18143 , n18140 , n18142 );
xor ( n18144 , n7332 , n7329 );
not ( n18145 , n18144 );
not ( n18146 , n15458 );
or ( n18147 , n18145 , n18146 );
or ( n18148 , n12685 , n18144 );
nand ( n18149 , n18147 , n18148 );
not ( n18150 , n18149 );
not ( n18151 , n8296 );
buf ( n18152 , n6006 );
not ( n18153 , n18152 );
not ( n18154 , n18153 );
or ( n18155 , n18151 , n18154 );
not ( n18156 , n8295 );
buf ( n18157 , n18152 );
nand ( n18158 , n18156 , n18157 );
nand ( n18159 , n18155 , n18158 );
buf ( n18160 , n6007 );
buf ( n18161 , n18160 );
and ( n18162 , n18159 , n18161 );
not ( n18163 , n18159 );
not ( n18164 , n18160 );
and ( n18165 , n18163 , n18164 );
nor ( n18166 , n18162 , n18165 );
buf ( n18167 , n6008 );
nand ( n18168 , n6622 , n18167 );
buf ( n18169 , n6009 );
buf ( n18170 , n18169 );
and ( n18171 , n18168 , n18170 );
not ( n18172 , n18168 );
not ( n18173 , n18169 );
and ( n18174 , n18172 , n18173 );
nor ( n18175 , n18171 , n18174 );
not ( n18176 , n18175 );
xor ( n18177 , n18166 , n18176 );
buf ( n18178 , n6010 );
nand ( n18179 , n8520 , n18178 );
buf ( n18180 , n6011 );
not ( n18181 , n18180 );
and ( n18182 , n18179 , n18181 );
not ( n18183 , n18179 );
buf ( n18184 , n18180 );
and ( n18185 , n18183 , n18184 );
nor ( n18186 , n18182 , n18185 );
xnor ( n18187 , n18177 , n18186 );
buf ( n18188 , n18187 );
not ( n18189 , n18188 );
and ( n18190 , n18150 , n18189 );
not ( n18191 , n18187 );
not ( n18192 , n18191 );
and ( n18193 , n18149 , n18192 );
nor ( n18194 , n18190 , n18193 );
nand ( n18195 , n18143 , n18194 );
xor ( n18196 , n11897 , n10498 );
xnor ( n18197 , n18196 , n9725 );
not ( n18198 , n18197 );
and ( n18199 , n18195 , n18198 );
not ( n18200 , n18195 );
and ( n18201 , n18200 , n18197 );
nor ( n18202 , n18199 , n18201 );
not ( n18203 , n18202 );
not ( n18204 , n18203 );
or ( n18205 , n18092 , n18204 );
nand ( n18206 , n18202 , n18090 );
nand ( n18207 , n18205 , n18206 );
and ( n18208 , n17991 , n18207 );
not ( n18209 , n17991 );
not ( n18210 , n18207 );
and ( n18211 , n18209 , n18210 );
nor ( n18212 , n18208 , n18211 );
not ( n18213 , n18212 );
or ( n18214 , n17729 , n18213 );
not ( n18215 , n17728 );
not ( n18216 , n18212 );
nand ( n18217 , n18215 , n18216 );
nand ( n18218 , n18214 , n18217 );
not ( n18219 , n13662 );
not ( n18220 , n18219 );
not ( n18221 , n14341 );
or ( n18222 , n18220 , n18221 );
or ( n18223 , n14341 , n18219 );
nand ( n18224 , n18222 , n18223 );
and ( n18225 , n18224 , n16845 );
not ( n18226 , n18224 );
not ( n18227 , n14384 );
and ( n18228 , n18226 , n18227 );
nor ( n18229 , n18225 , n18228 );
not ( n18230 , n18229 );
not ( n18231 , n18230 );
buf ( n18232 , n6012 );
not ( n18233 , n18232 );
buf ( n18234 , n6013 );
not ( n18235 , n18234 );
and ( n18236 , n18235 , n16808 );
not ( n18237 , n18235 );
and ( n18238 , n18237 , n16804 );
nor ( n18239 , n18236 , n18238 );
xor ( n18240 , n18233 , n18239 );
buf ( n18241 , n6014 );
buf ( n18242 , n6015 );
xor ( n18243 , n18241 , n18242 );
buf ( n18244 , n6016 );
nand ( n18245 , n7288 , n18244 );
xnor ( n18246 , n18243 , n18245 );
xnor ( n18247 , n18240 , n18246 );
not ( n18248 , n18247 );
not ( n18249 , n15701 );
buf ( n18250 , n6017 );
buf ( n18251 , n18250 );
not ( n18252 , n18251 );
not ( n18253 , n14162 );
not ( n18254 , n18253 );
or ( n18255 , n18252 , n18254 );
not ( n18256 , n18250 );
nand ( n18257 , n18256 , n14163 );
nand ( n18258 , n18255 , n18257 );
buf ( n18259 , n6018 );
not ( n18260 , n18259 );
and ( n18261 , n18258 , n18260 );
not ( n18262 , n18258 );
buf ( n18263 , n18259 );
and ( n18264 , n18262 , n18263 );
nor ( n18265 , n18261 , n18264 );
buf ( n18266 , n6019 );
nand ( n18267 , n8923 , n18266 );
buf ( n18268 , n6020 );
buf ( n18269 , n18268 );
and ( n18270 , n18267 , n18269 );
not ( n18271 , n18267 );
not ( n18272 , n18268 );
and ( n18273 , n18271 , n18272 );
nor ( n18274 , n18270 , n18273 );
xor ( n18275 , n18265 , n18274 );
buf ( n18276 , n6021 );
nand ( n18277 , n7133 , n18276 );
buf ( n18278 , n6022 );
buf ( n18279 , n18278 );
and ( n18280 , n18277 , n18279 );
not ( n18281 , n18277 );
not ( n18282 , n18278 );
and ( n18283 , n18281 , n18282 );
nor ( n18284 , n18280 , n18283 );
not ( n18285 , n18284 );
xnor ( n18286 , n18275 , n18285 );
not ( n18287 , n18286 );
or ( n18288 , n18249 , n18287 );
not ( n18289 , n15701 );
not ( n18290 , n18265 );
xor ( n18291 , n18290 , n18284 );
not ( n18292 , n18274 );
xnor ( n18293 , n18291 , n18292 );
nand ( n18294 , n18289 , n18293 );
nand ( n18295 , n18288 , n18294 );
not ( n18296 , n18295 );
or ( n18297 , n18248 , n18296 );
not ( n18298 , n18247 );
not ( n18299 , n18298 );
or ( n18300 , n18299 , n18295 );
nand ( n18301 , n18297 , n18300 );
buf ( n18302 , n6023 );
not ( n18303 , n18302 );
not ( n18304 , n18303 );
not ( n18305 , n18304 );
buf ( n18306 , n6024 );
buf ( n18307 , n18306 );
not ( n18308 , n18307 );
buf ( n18309 , n6025 );
not ( n18310 , n18309 );
not ( n18311 , n18310 );
or ( n18312 , n18308 , n18311 );
not ( n18313 , n18306 );
buf ( n18314 , n18309 );
nand ( n18315 , n18313 , n18314 );
nand ( n18316 , n18312 , n18315 );
buf ( n18317 , n6026 );
not ( n18318 , n18317 );
and ( n18319 , n18316 , n18318 );
not ( n18320 , n18316 );
buf ( n18321 , n18317 );
and ( n18322 , n18320 , n18321 );
nor ( n18323 , n18319 , n18322 );
xor ( n18324 , n18323 , n17894 );
buf ( n18325 , n6027 );
nand ( n18326 , n7750 , n18325 );
buf ( n18327 , n6028 );
buf ( n18328 , n18327 );
and ( n18329 , n18326 , n18328 );
not ( n18330 , n18326 );
not ( n18331 , n18327 );
and ( n18332 , n18330 , n18331 );
nor ( n18333 , n18329 , n18332 );
xnor ( n18334 , n18324 , n18333 );
not ( n18335 , n18334 );
not ( n18336 , n18335 );
or ( n18337 , n18305 , n18336 );
not ( n18338 , n18334 );
or ( n18339 , n18338 , n18304 );
nand ( n18340 , n18337 , n18339 );
buf ( n18341 , n6029 );
buf ( n18342 , n18341 );
not ( n18343 , n18342 );
buf ( n18344 , n6030 );
not ( n18345 , n18344 );
not ( n18346 , n18345 );
or ( n18347 , n18343 , n18346 );
not ( n18348 , n18341 );
buf ( n18349 , n18344 );
nand ( n18350 , n18348 , n18349 );
nand ( n18351 , n18347 , n18350 );
buf ( n18352 , n6031 );
buf ( n18353 , n18352 );
and ( n18354 , n18351 , n18353 );
not ( n18355 , n18351 );
not ( n18356 , n18352 );
and ( n18357 , n18355 , n18356 );
nor ( n18358 , n18354 , n18357 );
xor ( n18359 , n18358 , n9557 );
buf ( n18360 , n6032 );
nand ( n18361 , n7356 , n18360 );
buf ( n18362 , n6033 );
buf ( n18363 , n18362 );
and ( n18364 , n18361 , n18363 );
not ( n18365 , n18361 );
not ( n18366 , n18362 );
and ( n18367 , n18365 , n18366 );
nor ( n18368 , n18364 , n18367 );
xnor ( n18369 , n18359 , n18368 );
buf ( n18370 , n18369 );
and ( n18371 , n18340 , n18370 );
not ( n18372 , n18340 );
not ( n18373 , n18370 );
and ( n18374 , n18372 , n18373 );
nor ( n18375 , n18371 , n18374 );
nand ( n18376 , n18301 , n18375 );
not ( n18377 , n18376 );
or ( n18378 , n18231 , n18377 );
or ( n18379 , n18376 , n18230 );
nand ( n18380 , n18378 , n18379 );
not ( n18381 , n18380 );
not ( n18382 , n16063 );
buf ( n18383 , n6034 );
buf ( n18384 , n18383 );
not ( n18385 , n18384 );
buf ( n18386 , n6035 );
not ( n18387 , n18386 );
not ( n18388 , n18387 );
or ( n18389 , n18385 , n18388 );
not ( n18390 , n18383 );
buf ( n18391 , n18386 );
nand ( n18392 , n18390 , n18391 );
nand ( n18393 , n18389 , n18392 );
xor ( n18394 , n16999 , n18393 );
buf ( n18395 , n6036 );
buf ( n18396 , n6037 );
not ( n18397 , n18396 );
xor ( n18398 , n18395 , n18397 );
buf ( n18399 , n6038 );
nand ( n18400 , n7921 , n18399 );
xnor ( n18401 , n18398 , n18400 );
xnor ( n18402 , n18394 , n18401 );
not ( n18403 , n18402 );
not ( n18404 , n18403 );
or ( n18405 , n18382 , n18404 );
or ( n18406 , n18403 , n16063 );
nand ( n18407 , n18405 , n18406 );
not ( n18408 , n17191 );
not ( n18409 , n18408 );
and ( n18410 , n18407 , n18409 );
not ( n18411 , n18407 );
and ( n18412 , n18411 , n17200 );
nor ( n18413 , n18410 , n18412 );
buf ( n18414 , n6039 );
buf ( n18415 , n18414 );
not ( n18416 , n18415 );
not ( n18417 , n14797 );
or ( n18418 , n18416 , n18417 );
not ( n18419 , n18415 );
not ( n18420 , n14786 );
xor ( n18421 , n14777 , n18420 );
xnor ( n18422 , n18421 , n14796 );
nand ( n18423 , n18419 , n18422 );
nand ( n18424 , n18418 , n18423 );
and ( n18425 , n18424 , n10810 );
not ( n18426 , n18424 );
and ( n18427 , n18426 , n10809 );
nor ( n18428 , n18425 , n18427 );
not ( n18429 , n18428 );
nand ( n18430 , n18413 , n18429 );
not ( n18431 , n18430 );
not ( n18432 , n12012 );
buf ( n18433 , n6040 );
buf ( n18434 , n18433 );
not ( n18435 , n18434 );
buf ( n18436 , n6041 );
not ( n18437 , n18436 );
not ( n18438 , n18437 );
or ( n18439 , n18435 , n18438 );
not ( n18440 , n18433 );
buf ( n18441 , n18436 );
nand ( n18442 , n18440 , n18441 );
nand ( n18443 , n18439 , n18442 );
and ( n18444 , n18443 , n12808 );
not ( n18445 , n18443 );
and ( n18446 , n18445 , n12764 );
nor ( n18447 , n18444 , n18446 );
buf ( n18448 , n6042 );
nand ( n18449 , n7195 , n18448 );
buf ( n18450 , n6043 );
buf ( n18451 , n18450 );
and ( n18452 , n18449 , n18451 );
not ( n18453 , n18449 );
not ( n18454 , n18450 );
and ( n18455 , n18453 , n18454 );
nor ( n18456 , n18452 , n18455 );
xor ( n18457 , n18447 , n18456 );
xnor ( n18458 , n18457 , n13254 );
not ( n18459 , n18458 );
or ( n18460 , n18432 , n18459 );
or ( n18461 , n18458 , n12012 );
nand ( n18462 , n18460 , n18461 );
buf ( n18463 , n6044 );
buf ( n18464 , n18463 );
not ( n18465 , n18464 );
buf ( n18466 , n6045 );
not ( n18467 , n18466 );
not ( n18468 , n18467 );
or ( n18469 , n18465 , n18468 );
not ( n18470 , n18463 );
buf ( n18471 , n18466 );
nand ( n18472 , n18470 , n18471 );
nand ( n18473 , n18469 , n18472 );
buf ( n18474 , n6046 );
buf ( n18475 , n18474 );
and ( n18476 , n18473 , n18475 );
not ( n18477 , n18473 );
not ( n18478 , n18474 );
and ( n18479 , n18477 , n18478 );
nor ( n18480 , n18476 , n18479 );
buf ( n18481 , n6047 );
nand ( n18482 , n7195 , n18481 );
buf ( n18483 , n6048 );
buf ( n18484 , n18483 );
and ( n18485 , n18482 , n18484 );
not ( n18486 , n18482 );
not ( n18487 , n18483 );
and ( n18488 , n18486 , n18487 );
nor ( n18489 , n18485 , n18488 );
xor ( n18490 , n18480 , n18489 );
xnor ( n18491 , n18490 , n7731 );
and ( n18492 , n18462 , n18491 );
not ( n18493 , n18462 );
not ( n18494 , n18489 );
xor ( n18495 , n18480 , n18494 );
xnor ( n18496 , n18495 , n7731 );
buf ( n18497 , n18496 );
and ( n18498 , n18493 , n18497 );
nor ( n18499 , n18492 , n18498 );
not ( n18500 , n18499 );
and ( n18501 , n18431 , n18500 );
not ( n18502 , n18428 );
nand ( n18503 , n18502 , n18413 );
and ( n18504 , n18503 , n18499 );
nor ( n18505 , n18501 , n18504 );
not ( n18506 , n18505 );
or ( n18507 , n18381 , n18506 );
or ( n18508 , n18505 , n18380 );
nand ( n18509 , n18507 , n18508 );
buf ( n18510 , n6049 );
buf ( n18511 , n18510 );
buf ( n18512 , n6050 );
buf ( n18513 , n18512 );
not ( n18514 , n18513 );
buf ( n18515 , n6051 );
not ( n18516 , n18515 );
not ( n18517 , n18516 );
or ( n18518 , n18514 , n18517 );
not ( n18519 , n18512 );
buf ( n18520 , n18515 );
nand ( n18521 , n18519 , n18520 );
nand ( n18522 , n18518 , n18521 );
buf ( n18523 , n6052 );
buf ( n18524 , n18523 );
and ( n18525 , n18522 , n18524 );
not ( n18526 , n18522 );
not ( n18527 , n18523 );
and ( n18528 , n18526 , n18527 );
nor ( n18529 , n18525 , n18528 );
buf ( n18530 , n6053 );
nand ( n18531 , n7471 , n18530 );
buf ( n18532 , n6054 );
buf ( n18533 , n18532 );
and ( n18534 , n18531 , n18533 );
not ( n18535 , n18531 );
not ( n18536 , n18532 );
and ( n18537 , n18535 , n18536 );
nor ( n18538 , n18534 , n18537 );
xor ( n18539 , n18529 , n18538 );
buf ( n18540 , n6055 );
nand ( n18541 , n8740 , n18540 );
buf ( n18542 , n6056 );
not ( n18543 , n18542 );
and ( n18544 , n18541 , n18543 );
not ( n18545 , n18541 );
buf ( n18546 , n18542 );
and ( n18547 , n18545 , n18546 );
nor ( n18548 , n18544 , n18547 );
xor ( n18549 , n18539 , n18548 );
buf ( n18550 , n18549 );
xor ( n18551 , n18511 , n18550 );
xnor ( n18552 , n18551 , n7521 );
not ( n18553 , n18552 );
buf ( n18554 , n6057 );
buf ( n18555 , n18554 );
not ( n18556 , n18555 );
buf ( n18557 , n6058 );
buf ( n18558 , n18557 );
not ( n18559 , n18558 );
buf ( n18560 , n6059 );
not ( n18561 , n18560 );
not ( n18562 , n18561 );
or ( n18563 , n18559 , n18562 );
not ( n18564 , n18557 );
buf ( n18565 , n18560 );
nand ( n18566 , n18564 , n18565 );
nand ( n18567 , n18563 , n18566 );
and ( n18568 , n18567 , n16247 );
not ( n18569 , n18567 );
not ( n18570 , n16246 );
and ( n18571 , n18569 , n18570 );
nor ( n18572 , n18568 , n18571 );
buf ( n18573 , n6060 );
nand ( n18574 , n8821 , n18573 );
buf ( n18575 , n6061 );
buf ( n18576 , n18575 );
and ( n18577 , n18574 , n18576 );
not ( n18578 , n18574 );
not ( n18579 , n18575 );
and ( n18580 , n18578 , n18579 );
nor ( n18581 , n18577 , n18580 );
xor ( n18582 , n18572 , n18581 );
buf ( n18583 , n6062 );
nand ( n18584 , n7196 , n18583 );
buf ( n18585 , n6063 );
buf ( n18586 , n18585 );
and ( n18587 , n18584 , n18586 );
not ( n18588 , n18584 );
not ( n18589 , n18585 );
and ( n18590 , n18588 , n18589 );
nor ( n18591 , n18587 , n18590 );
buf ( n18592 , n18591 );
xor ( n18593 , n18582 , n18592 );
not ( n18594 , n18593 );
not ( n18595 , n18594 );
or ( n18596 , n18556 , n18595 );
or ( n18597 , n18594 , n18555 );
nand ( n18598 , n18596 , n18597 );
buf ( n18599 , n6064 );
nand ( n18600 , n8740 , n18599 );
buf ( n18601 , n6065 );
buf ( n18602 , n18601 );
and ( n18603 , n18600 , n18602 );
not ( n18604 , n18600 );
not ( n18605 , n18601 );
and ( n18606 , n18604 , n18605 );
nor ( n18607 , n18603 , n18606 );
not ( n18608 , n18607 );
buf ( n18609 , n6066 );
nand ( n18610 , n7133 , n18609 );
buf ( n18611 , n6067 );
not ( n18612 , n18611 );
and ( n18613 , n18610 , n18612 );
not ( n18614 , n18610 );
buf ( n18615 , n18611 );
and ( n18616 , n18614 , n18615 );
nor ( n18617 , n18613 , n18616 );
not ( n18618 , n18617 );
or ( n18619 , n18608 , n18618 );
or ( n18620 , n18607 , n18617 );
nand ( n18621 , n18619 , n18620 );
buf ( n18622 , n6068 );
buf ( n18623 , n18622 );
not ( n18624 , n18623 );
buf ( n18625 , n6069 );
not ( n18626 , n18625 );
not ( n18627 , n18626 );
or ( n18628 , n18624 , n18627 );
not ( n18629 , n18622 );
buf ( n18630 , n18625 );
nand ( n18631 , n18629 , n18630 );
nand ( n18632 , n18628 , n18631 );
buf ( n18633 , n6070 );
not ( n18634 , n18633 );
and ( n18635 , n18632 , n18634 );
not ( n18636 , n18632 );
buf ( n18637 , n18633 );
and ( n18638 , n18636 , n18637 );
nor ( n18639 , n18635 , n18638 );
and ( n18640 , n18621 , n18639 );
not ( n18641 , n18621 );
not ( n18642 , n18639 );
and ( n18643 , n18641 , n18642 );
nor ( n18644 , n18640 , n18643 );
buf ( n18645 , n18644 );
and ( n18646 , n18598 , n18645 );
not ( n18647 , n18598 );
not ( n18648 , n18617 );
xor ( n18649 , n18639 , n18648 );
xnor ( n18650 , n18649 , n18607 );
buf ( n18651 , n18650 );
and ( n18652 , n18647 , n18651 );
nor ( n18653 , n18646 , n18652 );
nand ( n18654 , n18553 , n18653 );
not ( n18655 , n18654 );
buf ( n18656 , n10494 );
xor ( n18657 , n11916 , n18656 );
xnor ( n18658 , n18657 , n9725 );
not ( n18659 , n18658 );
and ( n18660 , n18655 , n18659 );
and ( n18661 , n18654 , n18658 );
nor ( n18662 , n18660 , n18661 );
and ( n18663 , n18509 , n18662 );
not ( n18664 , n18509 );
not ( n18665 , n18662 );
and ( n18666 , n18664 , n18665 );
nor ( n18667 , n18663 , n18666 );
not ( n18668 , n18667 );
not ( n18669 , n18668 );
buf ( n18670 , n6071 );
nand ( n18671 , n8519 , n18670 );
buf ( n18672 , n6072 );
buf ( n18673 , n18672 );
and ( n18674 , n18671 , n18673 );
not ( n18675 , n18671 );
not ( n18676 , n18672 );
and ( n18677 , n18675 , n18676 );
nor ( n18678 , n18674 , n18677 );
buf ( n18679 , n18678 );
not ( n18680 , n15394 );
and ( n18681 , n18679 , n18680 );
not ( n18682 , n18679 );
and ( n18683 , n18682 , n15395 );
nor ( n18684 , n18681 , n18683 );
buf ( n18685 , n6073 );
buf ( n18686 , n18685 );
not ( n18687 , n18686 );
buf ( n18688 , n6074 );
not ( n18689 , n18688 );
not ( n18690 , n18689 );
or ( n18691 , n18687 , n18690 );
not ( n18692 , n18685 );
buf ( n18693 , n18688 );
nand ( n18694 , n18692 , n18693 );
nand ( n18695 , n18691 , n18694 );
buf ( n18696 , n6075 );
not ( n18697 , n18696 );
and ( n18698 , n18695 , n18697 );
not ( n18699 , n18695 );
buf ( n18700 , n18696 );
and ( n18701 , n18699 , n18700 );
nor ( n18702 , n18698 , n18701 );
buf ( n18703 , n6076 );
nand ( n18704 , n7082 , n18703 );
buf ( n18705 , n6077 );
buf ( n18706 , n18705 );
and ( n18707 , n18704 , n18706 );
not ( n18708 , n18704 );
not ( n18709 , n18705 );
and ( n18710 , n18708 , n18709 );
nor ( n18711 , n18707 , n18710 );
xor ( n18712 , n18702 , n18711 );
buf ( n18713 , n6078 );
nand ( n18714 , n6608 , n18713 );
buf ( n18715 , n6079 );
buf ( n18716 , n18715 );
and ( n18717 , n18714 , n18716 );
not ( n18718 , n18714 );
not ( n18719 , n18715 );
and ( n18720 , n18718 , n18719 );
nor ( n18721 , n18717 , n18720 );
not ( n18722 , n18721 );
xnor ( n18723 , n18712 , n18722 );
buf ( n18724 , n18723 );
and ( n18725 , n18684 , n18724 );
not ( n18726 , n18684 );
xor ( n18727 , n18702 , n18721 );
not ( n18728 , n18711 );
xor ( n18729 , n18727 , n18728 );
buf ( n18730 , n18729 );
and ( n18731 , n18726 , n18730 );
nor ( n18732 , n18725 , n18731 );
not ( n18733 , n18732 );
not ( n18734 , n18733 );
xor ( n18735 , n10096 , n10116 );
buf ( n18736 , n10105 );
xnor ( n18737 , n18735 , n18736 );
not ( n18738 , n18737 );
not ( n18739 , n18738 );
xor ( n18740 , n11068 , n18739 );
buf ( n18741 , n6080 );
not ( n18742 , n18741 );
buf ( n18743 , n6081 );
nand ( n18744 , n7920 , n18743 );
buf ( n18745 , n6082 );
buf ( n18746 , n18745 );
and ( n18747 , n18744 , n18746 );
not ( n18748 , n18744 );
not ( n18749 , n18745 );
and ( n18750 , n18748 , n18749 );
nor ( n18751 , n18747 , n18750 );
xor ( n18752 , n18742 , n18751 );
buf ( n18753 , n6083 );
nand ( n18754 , n7299 , n18753 );
buf ( n18755 , n6084 );
buf ( n18756 , n18755 );
and ( n18757 , n18754 , n18756 );
not ( n18758 , n18754 );
not ( n18759 , n18755 );
and ( n18760 , n18758 , n18759 );
nor ( n18761 , n18757 , n18760 );
xnor ( n18762 , n18752 , n18761 );
not ( n18763 , n18762 );
buf ( n18764 , n6085 );
buf ( n18765 , n18764 );
not ( n18766 , n18765 );
buf ( n18767 , n6086 );
not ( n18768 , n18767 );
not ( n18769 , n18768 );
or ( n18770 , n18766 , n18769 );
not ( n18771 , n18764 );
buf ( n18772 , n18767 );
nand ( n18773 , n18771 , n18772 );
nand ( n18774 , n18770 , n18773 );
not ( n18775 , n18774 );
not ( n18776 , n18775 );
and ( n18777 , n18763 , n18776 );
and ( n18778 , n18762 , n18775 );
nor ( n18779 , n18777 , n18778 );
buf ( n18780 , n18779 );
xnor ( n18781 , n18740 , n18780 );
not ( n18782 , n18781 );
buf ( n18783 , n6087 );
buf ( n18784 , n18783 );
not ( n18785 , n18784 );
not ( n18786 , n10641 );
or ( n18787 , n18785 , n18786 );
not ( n18788 , n10641 );
not ( n18789 , n18783 );
nand ( n18790 , n18788 , n18789 );
nand ( n18791 , n18787 , n18790 );
not ( n18792 , n11542 );
buf ( n18793 , n18792 );
not ( n18794 , n18793 );
and ( n18795 , n18791 , n18794 );
not ( n18796 , n18791 );
and ( n18797 , n18796 , n18793 );
nor ( n18798 , n18795 , n18797 );
nand ( n18799 , n18782 , n18798 );
not ( n18800 , n18799 );
or ( n18801 , n18734 , n18800 );
not ( n18802 , n18798 );
not ( n18803 , n18802 );
nand ( n18804 , n18803 , n18782 );
or ( n18805 , n18804 , n18733 );
nand ( n18806 , n18801 , n18805 );
buf ( n18807 , n6088 );
buf ( n18808 , n18807 );
not ( n18809 , n18808 );
buf ( n18810 , n12688 );
not ( n18811 , n15451 );
buf ( n18812 , n6089 );
not ( n18813 , n18812 );
not ( n18814 , n18813 );
or ( n18815 , n18811 , n18814 );
not ( n18816 , n15450 );
buf ( n18817 , n18812 );
nand ( n18818 , n18816 , n18817 );
nand ( n18819 , n18815 , n18818 );
buf ( n18820 , n18819 );
xor ( n18821 , n18810 , n18820 );
buf ( n18822 , n6090 );
nand ( n18823 , n7043 , n18822 );
buf ( n18824 , n6091 );
not ( n18825 , n18824 );
and ( n18826 , n18823 , n18825 );
not ( n18827 , n18823 );
buf ( n18828 , n18824 );
and ( n18829 , n18827 , n18828 );
nor ( n18830 , n18826 , n18829 );
not ( n18831 , n18830 );
not ( n18832 , n18831 );
buf ( n18833 , n6092 );
nand ( n18834 , n7043 , n18833 );
buf ( n18835 , n6093 );
buf ( n18836 , n18835 );
and ( n18837 , n18834 , n18836 );
not ( n18838 , n18834 );
not ( n18839 , n18835 );
and ( n18840 , n18838 , n18839 );
nor ( n18841 , n18837 , n18840 );
not ( n18842 , n18841 );
not ( n18843 , n18842 );
or ( n18844 , n18832 , n18843 );
nand ( n18845 , n18841 , n18830 );
nand ( n18846 , n18844 , n18845 );
xnor ( n18847 , n18821 , n18846 );
not ( n18848 , n18847 );
or ( n18849 , n18809 , n18848 );
xor ( n18850 , n12689 , n18819 );
xor ( n18851 , n18850 , n18846 );
or ( n18852 , n18851 , n18808 );
nand ( n18853 , n18849 , n18852 );
not ( n18854 , n7336 );
and ( n18855 , n18853 , n18854 );
not ( n18856 , n18853 );
and ( n18857 , n18856 , n7336 );
nor ( n18858 , n18855 , n18857 );
not ( n18859 , n18858 );
buf ( n18860 , n8584 );
not ( n18861 , n18860 );
buf ( n18862 , n6094 );
buf ( n18863 , n18862 );
not ( n18864 , n18863 );
not ( n18865 , n16381 );
not ( n18866 , n18865 );
or ( n18867 , n18864 , n18866 );
not ( n18868 , n18862 );
nand ( n18869 , n18868 , n16382 );
nand ( n18870 , n18867 , n18869 );
buf ( n18871 , n6095 );
not ( n18872 , n18871 );
and ( n18873 , n18870 , n18872 );
not ( n18874 , n18870 );
buf ( n18875 , n18871 );
and ( n18876 , n18874 , n18875 );
nor ( n18877 , n18873 , n18876 );
buf ( n18878 , n6096 );
nand ( n18879 , n6804 , n18878 );
buf ( n18880 , n6097 );
buf ( n18881 , n18880 );
and ( n18882 , n18879 , n18881 );
not ( n18883 , n18879 );
not ( n18884 , n18880 );
and ( n18885 , n18883 , n18884 );
nor ( n18886 , n18882 , n18885 );
xor ( n18887 , n18877 , n18886 );
buf ( n18888 , n6098 );
nand ( n18889 , n7299 , n18888 );
buf ( n18890 , n6099 );
buf ( n18891 , n18890 );
and ( n18892 , n18889 , n18891 );
not ( n18893 , n18889 );
not ( n18894 , n18890 );
and ( n18895 , n18893 , n18894 );
nor ( n18896 , n18892 , n18895 );
xor ( n18897 , n18887 , n18896 );
buf ( n18898 , n18897 );
not ( n18899 , n18898 );
or ( n18900 , n18861 , n18899 );
or ( n18901 , n18898 , n18860 );
nand ( n18902 , n18900 , n18901 );
buf ( n18903 , n13005 );
and ( n18904 , n18902 , n18903 );
not ( n18905 , n18902 );
buf ( n18906 , n13010 );
and ( n18907 , n18905 , n18906 );
nor ( n18908 , n18904 , n18907 );
not ( n18909 , n18908 );
nand ( n18910 , n18859 , n18909 );
not ( n18911 , n18910 );
not ( n18912 , n6618 );
buf ( n18913 , n6100 );
buf ( n18914 , n18913 );
not ( n18915 , n18914 );
buf ( n18916 , n6101 );
not ( n18917 , n18916 );
not ( n18918 , n18917 );
or ( n18919 , n18915 , n18918 );
not ( n18920 , n18913 );
buf ( n18921 , n18916 );
nand ( n18922 , n18920 , n18921 );
nand ( n18923 , n18919 , n18922 );
buf ( n18924 , n6102 );
buf ( n18925 , n18924 );
and ( n18926 , n18923 , n18925 );
not ( n18927 , n18923 );
not ( n18928 , n18924 );
and ( n18929 , n18927 , n18928 );
nor ( n18930 , n18926 , n18929 );
buf ( n18931 , n6103 );
nand ( n18932 , n8821 , n18931 );
buf ( n18933 , n6104 );
buf ( n18934 , n18933 );
and ( n18935 , n18932 , n18934 );
not ( n18936 , n18932 );
not ( n18937 , n18933 );
and ( n18938 , n18936 , n18937 );
nor ( n18939 , n18935 , n18938 );
xor ( n18940 , n18930 , n18939 );
buf ( n18941 , n6105 );
nand ( n18942 , n6985 , n18941 );
buf ( n18943 , n6106 );
buf ( n18944 , n18943 );
and ( n18945 , n18942 , n18944 );
not ( n18946 , n18942 );
not ( n18947 , n18943 );
and ( n18948 , n18946 , n18947 );
nor ( n18949 , n18945 , n18948 );
not ( n18950 , n18949 );
xnor ( n18951 , n18940 , n18950 );
buf ( n18952 , n18951 );
not ( n18953 , n18952 );
or ( n18954 , n18912 , n18953 );
or ( n18955 , n18952 , n6618 );
nand ( n18956 , n18954 , n18955 );
not ( n18957 , n8542 );
not ( n18958 , n15846 );
not ( n18959 , n18958 );
or ( n18960 , n18957 , n18959 );
not ( n18961 , n8541 );
nand ( n18962 , n18961 , n15847 );
nand ( n18963 , n18960 , n18962 );
buf ( n18964 , n6107 );
not ( n18965 , n18964 );
and ( n18966 , n18963 , n18965 );
not ( n18967 , n18963 );
buf ( n18968 , n18964 );
and ( n18969 , n18967 , n18968 );
nor ( n18970 , n18966 , n18969 );
buf ( n18971 , n6108 );
nand ( n18972 , n7126 , n18971 );
buf ( n18973 , n6109 );
buf ( n18974 , n18973 );
and ( n18975 , n18972 , n18974 );
not ( n18976 , n18972 );
not ( n18977 , n18973 );
and ( n18978 , n18976 , n18977 );
nor ( n18979 , n18975 , n18978 );
xor ( n18980 , n18970 , n18979 );
xnor ( n18981 , n18980 , n14904 );
not ( n18982 , n18981 );
buf ( n18983 , n18982 );
not ( n18984 , n18983 );
buf ( n18985 , n18984 );
xnor ( n18986 , n18956 , n18985 );
buf ( n18987 , n18986 );
not ( n18988 , n18987 );
and ( n18989 , n18911 , n18988 );
and ( n18990 , n18910 , n18987 );
nor ( n18991 , n18989 , n18990 );
xor ( n18992 , n18806 , n18991 );
not ( n18993 , n18992 );
or ( n18994 , n18669 , n18993 );
not ( n18995 , n18992 );
nand ( n18996 , n18995 , n18667 );
nand ( n18997 , n18994 , n18996 );
buf ( n18998 , n18997 );
and ( n18999 , n18218 , n18998 );
not ( n19000 , n18218 );
not ( n19001 , n18995 );
not ( n19002 , n18667 );
and ( n19003 , n19001 , n19002 );
and ( n19004 , n18995 , n18667 );
nor ( n19005 , n19003 , n19004 );
not ( n19006 , n19005 );
not ( n19007 , n19006 );
and ( n19008 , n19000 , n19007 );
nor ( n19009 , n18999 , n19008 );
not ( n19010 , n19009 );
nand ( n19011 , n16840 , n17628 , n19010 );
not ( n19012 , n16836 );
not ( n19013 , n19012 );
not ( n19014 , n19010 );
or ( n19015 , n19013 , n19014 );
buf ( n19016 , n13752 );
nor ( n19017 , n17628 , n19016 );
nand ( n19018 , n19015 , n19017 );
buf ( n19019 , n13766 );
nand ( n19020 , n19019 , n13678 );
nand ( n19021 , n19011 , n19018 , n19020 );
buf ( n19022 , n19021 );
buf ( n19023 , n19022 );
xor ( n19024 , n15810 , n15829 );
not ( n19025 , n15819 );
xnor ( n19026 , n19024 , n19025 );
xor ( n19027 , n9272 , n19026 );
xnor ( n19028 , n19027 , n12961 );
buf ( n19029 , n6110 );
not ( n19030 , n19029 );
buf ( n19031 , n6111 );
buf ( n19032 , n19031 );
not ( n19033 , n19032 );
buf ( n19034 , n6112 );
not ( n19035 , n19034 );
not ( n19036 , n19035 );
or ( n19037 , n19033 , n19036 );
not ( n19038 , n19031 );
buf ( n19039 , n19034 );
nand ( n19040 , n19038 , n19039 );
nand ( n19041 , n19037 , n19040 );
buf ( n19042 , n6113 );
buf ( n19043 , n19042 );
and ( n19044 , n19041 , n19043 );
not ( n19045 , n19041 );
not ( n19046 , n19042 );
and ( n19047 , n19045 , n19046 );
nor ( n19048 , n19044 , n19047 );
buf ( n19049 , n6114 );
nand ( n19050 , n7133 , n19049 );
buf ( n19051 , n6115 );
xor ( n19052 , n19050 , n19051 );
xor ( n19053 , n19048 , n19052 );
buf ( n19054 , n6116 );
nand ( n19055 , n8971 , n19054 );
buf ( n19056 , n6117 );
buf ( n19057 , n19056 );
and ( n19058 , n19055 , n19057 );
not ( n19059 , n19055 );
not ( n19060 , n19056 );
and ( n19061 , n19059 , n19060 );
nor ( n19062 , n19058 , n19061 );
xnor ( n19063 , n19053 , n19062 );
not ( n19064 , n19063 );
not ( n19065 , n19064 );
not ( n19066 , n19065 );
or ( n19067 , n19030 , n19066 );
or ( n19068 , n19065 , n19029 );
nand ( n19069 , n19067 , n19068 );
not ( n19070 , n19069 );
buf ( n19071 , n6118 );
buf ( n19072 , n19071 );
not ( n19073 , n19072 );
buf ( n19074 , n6119 );
not ( n19075 , n19074 );
not ( n19076 , n19075 );
or ( n19077 , n19073 , n19076 );
not ( n19078 , n19071 );
buf ( n19079 , n19074 );
nand ( n19080 , n19078 , n19079 );
nand ( n19081 , n19077 , n19080 );
buf ( n19082 , n6120 );
buf ( n19083 , n19082 );
and ( n19084 , n19081 , n19083 );
not ( n19085 , n19081 );
not ( n19086 , n19082 );
and ( n19087 , n19085 , n19086 );
nor ( n19088 , n19084 , n19087 );
buf ( n19089 , n6121 );
nand ( n19090 , n7288 , n19089 );
buf ( n19091 , n6122 );
buf ( n19092 , n19091 );
and ( n19093 , n19090 , n19092 );
not ( n19094 , n19090 );
not ( n19095 , n19091 );
and ( n19096 , n19094 , n19095 );
nor ( n19097 , n19093 , n19096 );
xor ( n19098 , n19088 , n19097 );
buf ( n19099 , n6123 );
nand ( n19100 , n6905 , n19099 );
buf ( n19101 , n6124 );
buf ( n19102 , n19101 );
and ( n19103 , n19100 , n19102 );
not ( n19104 , n19100 );
not ( n19105 , n19101 );
and ( n19106 , n19104 , n19105 );
nor ( n19107 , n19103 , n19106 );
not ( n19108 , n19107 );
xor ( n19109 , n19098 , n19108 );
buf ( n19110 , n19109 );
not ( n19111 , n19110 );
and ( n19112 , n19070 , n19111 );
and ( n19113 , n19069 , n19110 );
nor ( n19114 , n19112 , n19113 );
not ( n19115 , n19114 );
nand ( n19116 , n19028 , n19115 );
xor ( n19117 , n16118 , n13121 );
not ( n19118 , n8193 );
xnor ( n19119 , n19117 , n19118 );
not ( n19120 , n19119 );
and ( n19121 , n19116 , n19120 );
not ( n19122 , n19116 );
and ( n19123 , n19122 , n19119 );
nor ( n19124 , n19121 , n19123 );
not ( n19125 , n19124 );
not ( n19126 , n9725 );
not ( n19127 , n10271 );
not ( n19128 , n19127 );
not ( n19129 , n9776 );
not ( n19130 , n19129 );
or ( n19131 , n19128 , n19130 );
or ( n19132 , n9780 , n19127 );
nand ( n19133 , n19131 , n19132 );
not ( n19134 , n19133 );
and ( n19135 , n19126 , n19134 );
and ( n19136 , n9725 , n19133 );
nor ( n19137 , n19135 , n19136 );
not ( n19138 , n19137 );
not ( n19139 , n19138 );
not ( n19140 , n6955 );
not ( n19141 , n19140 );
not ( n19142 , n8208 );
and ( n19143 , n19141 , n19142 );
and ( n19144 , n19140 , n8208 );
nor ( n19145 , n19143 , n19144 );
buf ( n19146 , n6125 );
buf ( n19147 , n19146 );
not ( n19148 , n19147 );
not ( n19149 , n13278 );
not ( n19150 , n19149 );
or ( n19151 , n19148 , n19150 );
not ( n19152 , n19146 );
nand ( n19153 , n19152 , n13279 );
nand ( n19154 , n19151 , n19153 );
buf ( n19155 , n6126 );
buf ( n19156 , n19155 );
and ( n19157 , n19154 , n19156 );
not ( n19158 , n19154 );
not ( n19159 , n19155 );
and ( n19160 , n19158 , n19159 );
nor ( n19161 , n19157 , n19160 );
xor ( n19162 , n19161 , n17687 );
buf ( n19163 , n6127 );
nand ( n19164 , n9257 , n19163 );
buf ( n19165 , n6128 );
buf ( n19166 , n19165 );
and ( n19167 , n19164 , n19166 );
not ( n19168 , n19164 );
not ( n19169 , n19165 );
and ( n19170 , n19168 , n19169 );
nor ( n19171 , n19167 , n19170 );
buf ( n19172 , n19171 );
xnor ( n19173 , n19162 , n19172 );
buf ( n19174 , n19173 );
and ( n19175 , n19145 , n19174 );
not ( n19176 , n19145 );
not ( n19177 , n19171 );
not ( n19178 , n17686 );
or ( n19179 , n19177 , n19178 );
or ( n19180 , n19171 , n17686 );
nand ( n19181 , n19179 , n19180 );
and ( n19182 , n19181 , n19161 );
not ( n19183 , n19181 );
not ( n19184 , n19161 );
and ( n19185 , n19183 , n19184 );
nor ( n19186 , n19182 , n19185 );
buf ( n19187 , n19186 );
and ( n19188 , n19176 , n19187 );
nor ( n19189 , n19175 , n19188 );
not ( n19190 , n19189 );
buf ( n19191 , n6129 );
buf ( n19192 , n19191 );
not ( n19193 , n19192 );
not ( n19194 , n7055 );
or ( n19195 , n19193 , n19194 );
or ( n19196 , n7055 , n19192 );
nand ( n19197 , n19195 , n19196 );
not ( n19198 , n19197 );
not ( n19199 , n13046 );
not ( n19200 , n19199 );
not ( n19201 , n13066 );
or ( n19202 , n19200 , n19201 );
nand ( n19203 , n13065 , n13046 );
nand ( n19204 , n19202 , n19203 );
not ( n19205 , n19204 );
not ( n19206 , n19205 );
or ( n19207 , n19198 , n19206 );
not ( n19208 , n19197 );
buf ( n19209 , n19204 );
nand ( n19210 , n19208 , n19209 );
nand ( n19211 , n19207 , n19210 );
nand ( n19212 , n19190 , n19211 );
not ( n19213 , n19212 );
or ( n19214 , n19139 , n19213 );
or ( n19215 , n19212 , n19138 );
nand ( n19216 , n19214 , n19215 );
not ( n19217 , n19216 );
buf ( n19218 , n6130 );
buf ( n19219 , n19218 );
not ( n19220 , n19219 );
buf ( n19221 , n6131 );
not ( n19222 , n19221 );
not ( n19223 , n19222 );
or ( n19224 , n19220 , n19223 );
not ( n19225 , n19218 );
buf ( n19226 , n19221 );
nand ( n19227 , n19225 , n19226 );
nand ( n19228 , n19224 , n19227 );
not ( n19229 , n19228 );
xor ( n19230 , n17909 , n19229 );
buf ( n19231 , n6132 );
xor ( n19232 , n19231 , n8990 );
xnor ( n19233 , n19232 , n8984 );
xnor ( n19234 , n19230 , n19233 );
not ( n19235 , n19234 );
buf ( n19236 , n6133 );
buf ( n19237 , n19236 );
not ( n19238 , n19237 );
and ( n19239 , n19235 , n19238 );
and ( n19240 , n19234 , n19237 );
nor ( n19241 , n19239 , n19240 );
buf ( n19242 , n6134 );
buf ( n19243 , n19242 );
not ( n19244 , n19243 );
buf ( n19245 , n6135 );
not ( n19246 , n19245 );
not ( n19247 , n19246 );
or ( n19248 , n19244 , n19247 );
not ( n19249 , n19242 );
buf ( n19250 , n19245 );
nand ( n19251 , n19249 , n19250 );
nand ( n19252 , n19248 , n19251 );
not ( n19253 , n19252 );
buf ( n19254 , n6136 );
not ( n19255 , n19254 );
buf ( n19256 , n6137 );
nand ( n19257 , n7093 , n19256 );
buf ( n19258 , n6138 );
buf ( n19259 , n19258 );
and ( n19260 , n19257 , n19259 );
not ( n19261 , n19257 );
not ( n19262 , n19258 );
and ( n19263 , n19261 , n19262 );
nor ( n19264 , n19260 , n19263 );
xor ( n19265 , n19255 , n19264 );
buf ( n19266 , n6139 );
nand ( n19267 , n10204 , n19266 );
buf ( n19268 , n6140 );
buf ( n19269 , n19268 );
and ( n19270 , n19267 , n19269 );
not ( n19271 , n19267 );
not ( n19272 , n19268 );
and ( n19273 , n19271 , n19272 );
nor ( n19274 , n19270 , n19273 );
xnor ( n19275 , n19265 , n19274 );
not ( n19276 , n19275 );
not ( n19277 , n19276 );
or ( n19278 , n19253 , n19277 );
not ( n19279 , n19252 );
nand ( n19280 , n19275 , n19279 );
nand ( n19281 , n19278 , n19280 );
buf ( n19282 , n19281 );
not ( n19283 , n19282 );
and ( n19284 , n19241 , n19283 );
not ( n19285 , n19241 );
and ( n19286 , n19285 , n19282 );
nor ( n19287 , n19284 , n19286 );
not ( n19288 , n19287 );
not ( n19289 , n7997 );
nand ( n19290 , n19289 , n17109 );
not ( n19291 , n19290 );
nor ( n19292 , n17109 , n8001 );
nor ( n19293 , n19291 , n19292 );
not ( n19294 , n19293 );
not ( n19295 , n12587 );
not ( n19296 , n19295 );
or ( n19297 , n19294 , n19296 );
not ( n19298 , n19293 );
nand ( n19299 , n19298 , n12587 );
nand ( n19300 , n19297 , n19299 );
nand ( n19301 , n19288 , n19300 );
not ( n19302 , n19301 );
not ( n19303 , n9482 );
buf ( n19304 , n6141 );
buf ( n19305 , n19304 );
not ( n19306 , n19305 );
buf ( n19307 , n6142 );
not ( n19308 , n19307 );
not ( n19309 , n19308 );
or ( n19310 , n19306 , n19309 );
not ( n19311 , n19304 );
buf ( n19312 , n19307 );
nand ( n19313 , n19311 , n19312 );
nand ( n19314 , n19310 , n19313 );
buf ( n19315 , n6143 );
not ( n19316 , n19315 );
and ( n19317 , n19314 , n19316 );
not ( n19318 , n19314 );
buf ( n19319 , n19315 );
and ( n19320 , n19318 , n19319 );
nor ( n19321 , n19317 , n19320 );
buf ( n19322 , n6144 );
nand ( n19323 , n8519 , n19322 );
buf ( n19324 , n6145 );
buf ( n19325 , n19324 );
and ( n19326 , n19323 , n19325 );
not ( n19327 , n19323 );
not ( n19328 , n19324 );
and ( n19329 , n19327 , n19328 );
nor ( n19330 , n19326 , n19329 );
xor ( n19331 , n19321 , n19330 );
buf ( n19332 , n6146 );
nand ( n19333 , n7413 , n19332 );
buf ( n19334 , n6147 );
buf ( n19335 , n19334 );
and ( n19336 , n19333 , n19335 );
not ( n19337 , n19333 );
not ( n19338 , n19334 );
and ( n19339 , n19337 , n19338 );
nor ( n19340 , n19336 , n19339 );
xor ( n19341 , n19331 , n19340 );
not ( n19342 , n19341 );
not ( n19343 , n19342 );
not ( n19344 , n19343 );
or ( n19345 , n19303 , n19344 );
buf ( n19346 , n19341 );
or ( n19347 , n19346 , n9482 );
nand ( n19348 , n19345 , n19347 );
not ( n19349 , n8847 );
not ( n19350 , n19349 );
and ( n19351 , n19348 , n19350 );
not ( n19352 , n19348 );
buf ( n19353 , n8846 );
and ( n19354 , n19352 , n19353 );
nor ( n19355 , n19351 , n19354 );
not ( n19356 , n19355 );
not ( n19357 , n19356 );
and ( n19358 , n19302 , n19357 );
and ( n19359 , n19301 , n19356 );
nor ( n19360 , n19358 , n19359 );
not ( n19361 , n19360 );
or ( n19362 , n19217 , n19361 );
or ( n19363 , n19360 , n19216 );
nand ( n19364 , n19362 , n19363 );
not ( n19365 , n19028 );
nand ( n19366 , n19120 , n19365 );
not ( n19367 , n7626 );
not ( n19368 , n10943 );
or ( n19369 , n19367 , n19368 );
or ( n19370 , n10943 , n7626 );
nand ( n19371 , n19369 , n19370 );
buf ( n19372 , n6148 );
buf ( n19373 , n6149 );
buf ( n19374 , n19373 );
not ( n19375 , n19374 );
buf ( n19376 , n6150 );
not ( n19377 , n19376 );
not ( n19378 , n19377 );
or ( n19379 , n19375 , n19378 );
not ( n19380 , n19373 );
buf ( n19381 , n19376 );
nand ( n19382 , n19380 , n19381 );
nand ( n19383 , n19379 , n19382 );
xor ( n19384 , n19372 , n19383 );
buf ( n19385 , n6151 );
xor ( n19386 , n16095 , n19385 );
buf ( n19387 , n6152 );
nand ( n19388 , n6817 , n19387 );
xnor ( n19389 , n19386 , n19388 );
xnor ( n19390 , n19384 , n19389 );
buf ( n19391 , n19390 );
buf ( n19392 , n19391 );
not ( n19393 , n19392 );
and ( n19394 , n19371 , n19393 );
not ( n19395 , n19371 );
and ( n19396 , n19395 , n19392 );
nor ( n19397 , n19394 , n19396 );
not ( n19398 , n19397 );
and ( n19399 , n19366 , n19398 );
not ( n19400 , n19366 );
and ( n19401 , n19400 , n19397 );
nor ( n19402 , n19399 , n19401 );
and ( n19403 , n19364 , n19402 );
not ( n19404 , n19364 );
not ( n19405 , n19402 );
and ( n19406 , n19404 , n19405 );
nor ( n19407 , n19403 , n19406 );
not ( n19408 , n19407 );
not ( n19409 , n19408 );
not ( n19410 , n12435 );
not ( n19411 , n15369 );
not ( n19412 , n19411 );
or ( n19413 , n19410 , n19412 );
or ( n19414 , n16955 , n12435 );
nand ( n19415 , n19413 , n19414 );
not ( n19416 , n18680 );
xor ( n19417 , n19415 , n19416 );
not ( n19418 , n19417 );
not ( n19419 , n10714 );
buf ( n19420 , n6153 );
buf ( n19421 , n19420 );
not ( n19422 , n19421 );
buf ( n19423 , n6154 );
not ( n19424 , n19423 );
not ( n19425 , n19424 );
or ( n19426 , n19422 , n19425 );
not ( n19427 , n19420 );
buf ( n19428 , n19423 );
nand ( n19429 , n19427 , n19428 );
nand ( n19430 , n19426 , n19429 );
buf ( n19431 , n6155 );
not ( n19432 , n19431 );
and ( n19433 , n19430 , n19432 );
not ( n19434 , n19430 );
buf ( n19435 , n19431 );
and ( n19436 , n19434 , n19435 );
nor ( n19437 , n19433 , n19436 );
not ( n19438 , n19437 );
buf ( n19439 , n6156 );
nand ( n19440 , n6706 , n19439 );
buf ( n19441 , n6157 );
buf ( n19442 , n19441 );
and ( n19443 , n19440 , n19442 );
not ( n19444 , n19440 );
not ( n19445 , n19441 );
and ( n19446 , n19444 , n19445 );
nor ( n19447 , n19443 , n19446 );
xor ( n19448 , n19438 , n19447 );
xnor ( n19449 , n19448 , n17495 );
not ( n19450 , n19449 );
or ( n19451 , n19419 , n19450 );
not ( n19452 , n19449 );
nand ( n19453 , n19452 , n10710 );
nand ( n19454 , n19451 , n19453 );
not ( n19455 , n14223 );
buf ( n19456 , n6158 );
not ( n19457 , n19456 );
not ( n19458 , n19457 );
or ( n19459 , n19455 , n19458 );
not ( n19460 , n14222 );
buf ( n19461 , n19456 );
nand ( n19462 , n19460 , n19461 );
nand ( n19463 , n19459 , n19462 );
buf ( n19464 , n6159 );
buf ( n19465 , n19464 );
and ( n19466 , n19463 , n19465 );
not ( n19467 , n19463 );
not ( n19468 , n19464 );
and ( n19469 , n19467 , n19468 );
nor ( n19470 , n19466 , n19469 );
buf ( n19471 , n6160 );
nand ( n19472 , n6660 , n19471 );
buf ( n19473 , n6161 );
buf ( n19474 , n19473 );
and ( n19475 , n19472 , n19474 );
not ( n19476 , n19472 );
not ( n19477 , n19473 );
and ( n19478 , n19476 , n19477 );
nor ( n19479 , n19475 , n19478 );
xor ( n19480 , n19470 , n19479 );
buf ( n19481 , n6162 );
nand ( n19482 , n8269 , n19481 );
buf ( n19483 , n6163 );
buf ( n19484 , n19483 );
and ( n19485 , n19482 , n19484 );
not ( n19486 , n19482 );
not ( n19487 , n19483 );
and ( n19488 , n19486 , n19487 );
nor ( n19489 , n19485 , n19488 );
xnor ( n19490 , n19480 , n19489 );
not ( n19491 , n19490 );
not ( n19492 , n19491 );
not ( n19493 , n19492 );
and ( n19494 , n19454 , n19493 );
not ( n19495 , n19454 );
buf ( n19496 , n19492 );
and ( n19497 , n19495 , n19496 );
nor ( n19498 , n19494 , n19497 );
nand ( n19499 , n19418 , n19498 );
not ( n19500 , n19499 );
buf ( n19501 , n6164 );
nand ( n19502 , n6761 , n19501 );
buf ( n19503 , n6165 );
not ( n19504 , n19503 );
and ( n19505 , n19502 , n19504 );
not ( n19506 , n19502 );
buf ( n19507 , n19503 );
and ( n19508 , n19506 , n19507 );
nor ( n19509 , n19505 , n19508 );
xor ( n19510 , n19509 , n17390 );
xnor ( n19511 , n19510 , n15254 );
not ( n19512 , n19511 );
not ( n19513 , n19512 );
or ( n19514 , n19500 , n19513 );
or ( n19515 , n19512 , n19499 );
nand ( n19516 , n19514 , n19515 );
not ( n19517 , n19516 );
not ( n19518 , n14259 );
not ( n19519 , n17823 );
or ( n19520 , n19518 , n19519 );
nand ( n19521 , n17824 , n14255 );
nand ( n19522 , n19520 , n19521 );
buf ( n19523 , n18286 );
and ( n19524 , n19522 , n19523 );
not ( n19525 , n19522 );
buf ( n19526 , n18293 );
and ( n19527 , n19525 , n19526 );
nor ( n19528 , n19524 , n19527 );
not ( n19529 , n18817 );
not ( n19530 , n12743 );
or ( n19531 , n19529 , n19530 );
buf ( n19532 , n12730 );
nand ( n19533 , n19532 , n18813 );
nand ( n19534 , n19531 , n19533 );
not ( n19535 , n12749 );
and ( n19536 , n19534 , n19535 );
not ( n19537 , n19534 );
and ( n19538 , n19537 , n12749 );
nor ( n19539 , n19536 , n19538 );
and ( n19540 , n19528 , n19539 );
buf ( n19541 , n6166 );
nand ( n19542 , n7477 , n19541 );
buf ( n19543 , n6167 );
buf ( n19544 , n19543 );
and ( n19545 , n19542 , n19544 );
not ( n19546 , n19542 );
not ( n19547 , n19543 );
and ( n19548 , n19546 , n19547 );
nor ( n19549 , n19545 , n19548 );
buf ( n19550 , n19549 );
not ( n19551 , n19550 );
not ( n19552 , n12525 );
not ( n19553 , n19552 );
or ( n19554 , n19551 , n19553 );
or ( n19555 , n19552 , n19550 );
nand ( n19556 , n19554 , n19555 );
and ( n19557 , n19556 , n12532 );
not ( n19558 , n19556 );
not ( n19559 , n12532 );
and ( n19560 , n19558 , n19559 );
nor ( n19561 , n19557 , n19560 );
not ( n19562 , n19561 );
not ( n19563 , n19562 );
and ( n19564 , n19540 , n19563 );
not ( n19565 , n19540 );
and ( n19566 , n19565 , n19562 );
nor ( n19567 , n19564 , n19566 );
not ( n19568 , n19567 );
and ( n19569 , n19517 , n19568 );
and ( n19570 , n19516 , n19567 );
nor ( n19571 , n19569 , n19570 );
not ( n19572 , n19571 );
not ( n19573 , n19572 );
and ( n19574 , n19409 , n19573 );
and ( n19575 , n19408 , n19572 );
nor ( n19576 , n19574 , n19575 );
not ( n19577 , n19576 );
or ( n19578 , n19125 , n19577 );
not ( n19579 , n19571 );
not ( n19580 , n19407 );
or ( n19581 , n19579 , n19580 );
not ( n19582 , n19407 );
nand ( n19583 , n19582 , n19572 );
nand ( n19584 , n19581 , n19583 );
not ( n19585 , n19124 );
nand ( n19586 , n19584 , n19585 );
nand ( n19587 , n19578 , n19586 );
buf ( n19588 , n6168 );
not ( n19589 , n19588 );
buf ( n19590 , n6169 );
buf ( n19591 , n19590 );
not ( n19592 , n19591 );
not ( n19593 , n19236 );
not ( n19594 , n19593 );
or ( n19595 , n19592 , n19594 );
not ( n19596 , n19590 );
nand ( n19597 , n19596 , n19237 );
nand ( n19598 , n19595 , n19597 );
buf ( n19599 , n6170 );
not ( n19600 , n19599 );
and ( n19601 , n19598 , n19600 );
not ( n19602 , n19598 );
buf ( n19603 , n19599 );
and ( n19604 , n19602 , n19603 );
nor ( n19605 , n19601 , n19604 );
buf ( n19606 , n6171 );
nand ( n19607 , n6706 , n19606 );
buf ( n19608 , n6172 );
buf ( n19609 , n19608 );
and ( n19610 , n19607 , n19609 );
not ( n19611 , n19607 );
not ( n19612 , n19608 );
and ( n19613 , n19611 , n19612 );
nor ( n19614 , n19610 , n19613 );
xor ( n19615 , n19605 , n19614 );
buf ( n19616 , n6173 );
nand ( n19617 , n7750 , n19616 );
buf ( n19618 , n6174 );
buf ( n19619 , n19618 );
and ( n19620 , n19617 , n19619 );
not ( n19621 , n19617 );
not ( n19622 , n19618 );
and ( n19623 , n19621 , n19622 );
nor ( n19624 , n19620 , n19623 );
xor ( n19625 , n19615 , n19624 );
buf ( n19626 , n19625 );
not ( n19627 , n19626 );
or ( n19628 , n19589 , n19627 );
or ( n19629 , n19626 , n19588 );
nand ( n19630 , n19628 , n19629 );
not ( n19631 , n8760 );
and ( n19632 , n19630 , n19631 );
not ( n19633 , n19630 );
buf ( n19634 , n8760 );
and ( n19635 , n19633 , n19634 );
nor ( n19636 , n19632 , n19635 );
not ( n19637 , n19636 );
not ( n19638 , n12198 );
not ( n19639 , n11058 );
or ( n19640 , n19638 , n19639 );
or ( n19641 , n11058 , n12198 );
nand ( n19642 , n19640 , n19641 );
not ( n19643 , n19642 );
xor ( n19644 , n17429 , n17439 );
xnor ( n19645 , n19644 , n16042 );
buf ( n19646 , n19645 );
not ( n19647 , n19646 );
and ( n19648 , n19643 , n19647 );
and ( n19649 , n19642 , n19646 );
nor ( n19650 , n19648 , n19649 );
not ( n19651 , n19650 );
nand ( n19652 , n19637 , n19651 );
not ( n19653 , n19652 );
xor ( n19654 , n8244 , n6957 );
not ( n19655 , n6890 );
xor ( n19656 , n19655 , n6900 );
xnor ( n19657 , n19656 , n6909 );
buf ( n19658 , n19657 );
xnor ( n19659 , n19654 , n19658 );
not ( n19660 , n19659 );
not ( n19661 , n19660 );
or ( n19662 , n19653 , n19661 );
or ( n19663 , n19660 , n19652 );
nand ( n19664 , n19662 , n19663 );
not ( n19665 , n12870 );
xor ( n19666 , n16394 , n19665 );
xnor ( n19667 , n19666 , n17229 );
not ( n19668 , n16285 );
not ( n19669 , n19668 );
not ( n19670 , n11867 );
nor ( n19671 , n19670 , n18592 );
not ( n19672 , n19671 );
nand ( n19673 , n18592 , n19670 );
nand ( n19674 , n19672 , n19673 );
not ( n19675 , n19674 );
or ( n19676 , n19669 , n19675 );
or ( n19677 , n19674 , n16289 );
nand ( n19678 , n19676 , n19677 );
nand ( n19679 , n19667 , n19678 );
not ( n19680 , n19679 );
buf ( n19681 , n6175 );
buf ( n19682 , n19681 );
not ( n19683 , n19682 );
not ( n19684 , n11261 );
or ( n19685 , n19683 , n19684 );
not ( n19686 , n19681 );
nand ( n19687 , n11260 , n19686 );
nand ( n19688 , n19685 , n19687 );
not ( n19689 , n19688 );
not ( n19690 , n11228 );
not ( n19691 , n19690 );
not ( n19692 , n19691 );
or ( n19693 , n19689 , n19692 );
or ( n19694 , n19691 , n19688 );
nand ( n19695 , n19693 , n19694 );
not ( n19696 , n19695 );
and ( n19697 , n19680 , n19696 );
and ( n19698 , n19679 , n19695 );
nor ( n19699 , n19697 , n19698 );
xor ( n19700 , n19664 , n19699 );
not ( n19701 , n19700 );
buf ( n19702 , n6176 );
buf ( n19703 , n19702 );
not ( n19704 , n19703 );
not ( n19705 , n11948 );
or ( n19706 , n19704 , n19705 );
not ( n19707 , n19703 );
nand ( n19708 , n19707 , n9948 );
nand ( n19709 , n19706 , n19708 );
not ( n19710 , n19709 );
not ( n19711 , n16737 );
and ( n19712 , n19710 , n19711 );
and ( n19713 , n19709 , n11997 );
nor ( n19714 , n19712 , n19713 );
not ( n19715 , n19714 );
not ( n19716 , n19715 );
not ( n19717 , n9244 );
nor ( n19718 , n14723 , n16971 );
not ( n19719 , n19718 );
nand ( n19720 , n14723 , n16971 );
nand ( n19721 , n19719 , n19720 );
not ( n19722 , n19721 );
and ( n19723 , n19717 , n19722 );
not ( n19724 , n15440 );
and ( n19725 , n19724 , n19721 );
nor ( n19726 , n19723 , n19725 );
not ( n19727 , n13618 );
not ( n19728 , n19727 );
buf ( n19729 , n15598 );
not ( n19730 , n19729 );
not ( n19731 , n17666 );
or ( n19732 , n19730 , n19731 );
not ( n19733 , n19729 );
nand ( n19734 , n19733 , n17667 );
nand ( n19735 , n19732 , n19734 );
not ( n19736 , n19735 );
or ( n19737 , n19728 , n19736 );
not ( n19738 , n13618 );
or ( n19739 , n19735 , n19738 );
nand ( n19740 , n19737 , n19739 );
nand ( n19741 , n19726 , n19740 );
not ( n19742 , n19741 );
or ( n19743 , n19716 , n19742 );
or ( n19744 , n19741 , n19715 );
nand ( n19745 , n19743 , n19744 );
not ( n19746 , n19745 );
not ( n19747 , n6965 );
buf ( n19748 , n6177 );
not ( n19749 , n19748 );
not ( n19750 , n19749 );
or ( n19751 , n19747 , n19750 );
not ( n19752 , n6964 );
buf ( n19753 , n19748 );
nand ( n19754 , n19752 , n19753 );
nand ( n19755 , n19751 , n19754 );
and ( n19756 , n19755 , n12095 );
not ( n19757 , n19755 );
not ( n19758 , n12094 );
and ( n19759 , n19757 , n19758 );
nor ( n19760 , n19756 , n19759 );
buf ( n19761 , n6178 );
nand ( n19762 , n7616 , n19761 );
buf ( n19763 , n6179 );
xor ( n19764 , n19762 , n19763 );
xor ( n19765 , n19760 , n19764 );
buf ( n19766 , n6180 );
nand ( n19767 , n7134 , n19766 );
buf ( n19768 , n6181 );
not ( n19769 , n19768 );
and ( n19770 , n19767 , n19769 );
not ( n19771 , n19767 );
buf ( n19772 , n19768 );
and ( n19773 , n19771 , n19772 );
nor ( n19774 , n19770 , n19773 );
xor ( n19775 , n19765 , n19774 );
xor ( n19776 , n7176 , n19775 );
buf ( n19777 , n6182 );
not ( n19778 , n19777 );
buf ( n19779 , n6183 );
buf ( n19780 , n19779 );
not ( n19781 , n19780 );
not ( n19782 , n11277 );
not ( n19783 , n19782 );
or ( n19784 , n19781 , n19783 );
not ( n19785 , n19779 );
nand ( n19786 , n19785 , n11278 );
nand ( n19787 , n19784 , n19786 );
xor ( n19788 , n19778 , n19787 );
buf ( n19789 , n6184 );
nand ( n19790 , n6816 , n19789 );
buf ( n19791 , n6185 );
buf ( n19792 , n19791 );
and ( n19793 , n19790 , n19792 );
not ( n19794 , n19790 );
not ( n19795 , n19791 );
and ( n19796 , n19794 , n19795 );
nor ( n19797 , n19793 , n19796 );
not ( n19798 , n19797 );
buf ( n19799 , n6186 );
not ( n19800 , n19799 );
and ( n19801 , n19798 , n19800 );
and ( n19802 , n19797 , n19799 );
nor ( n19803 , n19801 , n19802 );
xor ( n19804 , n19788 , n19803 );
not ( n19805 , n19804 );
xnor ( n19806 , n19776 , n19805 );
buf ( n19807 , n6187 );
nand ( n19808 , n7471 , n19807 );
buf ( n19809 , n6188 );
buf ( n19810 , n19809 );
and ( n19811 , n19808 , n19810 );
not ( n19812 , n19808 );
not ( n19813 , n19809 );
and ( n19814 , n19812 , n19813 );
nor ( n19815 , n19811 , n19814 );
buf ( n19816 , n19815 );
not ( n19817 , n19816 );
xor ( n19818 , n19048 , n19052 );
xnor ( n19819 , n19818 , n19062 );
not ( n19820 , n19819 );
not ( n19821 , n19820 );
or ( n19822 , n19817 , n19821 );
or ( n19823 , n19820 , n19816 );
nand ( n19824 , n19822 , n19823 );
xor ( n19825 , n19088 , n19107 );
not ( n19826 , n19097 );
xnor ( n19827 , n19825 , n19826 );
not ( n19828 , n19827 );
not ( n19829 , n19828 );
and ( n19830 , n19824 , n19829 );
not ( n19831 , n19824 );
and ( n19832 , n19831 , n19110 );
nor ( n19833 , n19830 , n19832 );
nand ( n19834 , n19806 , n19833 );
not ( n19835 , n14232 );
not ( n19836 , n17780 );
or ( n19837 , n19835 , n19836 );
nand ( n19838 , n17781 , n14227 );
nand ( n19839 , n19837 , n19838 );
not ( n19840 , n19839 );
not ( n19841 , n17823 );
and ( n19842 , n19840 , n19841 );
and ( n19843 , n19839 , n17828 );
nor ( n19844 , n19842 , n19843 );
not ( n19845 , n19844 );
and ( n19846 , n19834 , n19845 );
not ( n19847 , n19834 );
and ( n19848 , n19847 , n19844 );
nor ( n19849 , n19846 , n19848 );
not ( n19850 , n19849 );
or ( n19851 , n19746 , n19850 );
or ( n19852 , n19849 , n19745 );
nand ( n19853 , n19851 , n19852 );
xor ( n19854 , n9952 , n15503 );
buf ( n19855 , n6189 );
not ( n19856 , n19855 );
and ( n19857 , n19856 , n18808 );
not ( n19858 , n19856 );
not ( n19859 , n18807 );
and ( n19860 , n19858 , n19859 );
nor ( n19861 , n19857 , n19860 );
not ( n19862 , n19861 );
buf ( n19863 , n6190 );
buf ( n19864 , n6191 );
nand ( n19865 , n7412 , n19864 );
buf ( n19866 , n6192 );
buf ( n19867 , n19866 );
and ( n19868 , n19865 , n19867 );
not ( n19869 , n19865 );
not ( n19870 , n19866 );
and ( n19871 , n19869 , n19870 );
nor ( n19872 , n19868 , n19871 );
xor ( n19873 , n19863 , n19872 );
buf ( n19874 , n6193 );
nand ( n19875 , n7288 , n19874 );
buf ( n19876 , n6194 );
not ( n19877 , n19876 );
and ( n19878 , n19875 , n19877 );
not ( n19879 , n19875 );
buf ( n19880 , n19876 );
and ( n19881 , n19879 , n19880 );
nor ( n19882 , n19878 , n19881 );
xnor ( n19883 , n19873 , n19882 );
not ( n19884 , n19883 );
or ( n19885 , n19862 , n19884 );
or ( n19886 , n19883 , n19861 );
nand ( n19887 , n19885 , n19886 );
buf ( n19888 , n19887 );
not ( n19889 , n19888 );
xnor ( n19890 , n19854 , n19889 );
buf ( n19891 , n17479 );
not ( n19892 , n19891 );
not ( n19893 , n7977 );
or ( n19894 , n19892 , n19893 );
or ( n19895 , n7977 , n19891 );
nand ( n19896 , n19894 , n19895 );
buf ( n19897 , n6195 );
not ( n19898 , n19897 );
buf ( n19899 , n6196 );
buf ( n19900 , n19899 );
and ( n19901 , n19898 , n19900 );
not ( n19902 , n19898 );
not ( n19903 , n19899 );
and ( n19904 , n19902 , n19903 );
nor ( n19905 , n19901 , n19904 );
not ( n19906 , n19905 );
not ( n19907 , n19906 );
xor ( n19908 , n19029 , n19815 );
buf ( n19909 , n6197 );
nand ( n19910 , n8785 , n19909 );
buf ( n19911 , n6198 );
not ( n19912 , n19911 );
and ( n19913 , n19910 , n19912 );
not ( n19914 , n19910 );
buf ( n19915 , n19911 );
and ( n19916 , n19914 , n19915 );
nor ( n19917 , n19913 , n19916 );
xnor ( n19918 , n19908 , n19917 );
not ( n19919 , n19918 );
not ( n19920 , n19919 );
or ( n19921 , n19907 , n19920 );
nand ( n19922 , n19918 , n19905 );
nand ( n19923 , n19921 , n19922 );
buf ( n19924 , n19923 );
and ( n19925 , n19896 , n19924 );
not ( n19926 , n19896 );
not ( n19927 , n19918 );
not ( n19928 , n19905 );
and ( n19929 , n19927 , n19928 );
and ( n19930 , n19918 , n19905 );
nor ( n19931 , n19929 , n19930 );
buf ( n19932 , n19931 );
and ( n19933 , n19926 , n19932 );
nor ( n19934 , n19925 , n19933 );
nand ( n19935 , n19890 , n19934 );
buf ( n19936 , n6199 );
buf ( n19937 , n19936 );
not ( n19938 , n19937 );
not ( n19939 , n8887 );
not ( n19940 , n19939 );
not ( n19941 , n19940 );
or ( n19942 , n19938 , n19941 );
not ( n19943 , n8888 );
or ( n19944 , n19943 , n19937 );
nand ( n19945 , n19942 , n19944 );
not ( n19946 , n19945 );
buf ( n19947 , n6200 );
buf ( n19948 , n19947 );
buf ( n19949 , n6201 );
not ( n19950 , n19949 );
buf ( n19951 , n6202 );
buf ( n19952 , n19951 );
nand ( n19953 , n19950 , n19952 );
not ( n19954 , n19951 );
buf ( n19955 , n19949 );
nand ( n19956 , n19954 , n19955 );
and ( n19957 , n19953 , n19956 );
xor ( n19958 , n19948 , n19957 );
buf ( n19959 , n6203 );
buf ( n19960 , n6204 );
xor ( n19961 , n19959 , n19960 );
buf ( n19962 , n6205 );
nand ( n19963 , n6761 , n19962 );
xnor ( n19964 , n19961 , n19963 );
xnor ( n19965 , n19958 , n19964 );
not ( n19966 , n19965 );
not ( n19967 , n19966 );
or ( n19968 , n19946 , n19967 );
not ( n19969 , n19965 );
not ( n19970 , n19969 );
not ( n19971 , n19970 );
or ( n19972 , n19971 , n19945 );
nand ( n19973 , n19968 , n19972 );
not ( n19974 , n19973 );
and ( n19975 , n19935 , n19974 );
not ( n19976 , n19935 );
and ( n19977 , n19976 , n19973 );
nor ( n19978 , n19975 , n19977 );
and ( n19979 , n19853 , n19978 );
not ( n19980 , n19853 );
not ( n19981 , n19978 );
and ( n19982 , n19980 , n19981 );
nor ( n19983 , n19979 , n19982 );
not ( n19984 , n19983 );
or ( n19985 , n19701 , n19984 );
not ( n19986 , n19983 );
not ( n19987 , n19700 );
nand ( n19988 , n19986 , n19987 );
nand ( n19989 , n19985 , n19988 );
buf ( n19990 , n19989 );
and ( n19991 , n19587 , n19990 );
not ( n19992 , n19587 );
and ( n19993 , n19983 , n19700 );
not ( n19994 , n19983 );
and ( n19995 , n19994 , n19987 );
nor ( n19996 , n19993 , n19995 );
buf ( n19997 , n19996 );
and ( n19998 , n19992 , n19997 );
nor ( n19999 , n19991 , n19998 );
not ( n20000 , n19999 );
not ( n20001 , n16838 );
nor ( n20002 , n20000 , n20001 );
not ( n20003 , n20002 );
buf ( n20004 , n6206 );
nand ( n20005 , n8387 , n20004 );
buf ( n20006 , n6207 );
buf ( n20007 , n20006 );
and ( n20008 , n20005 , n20007 );
not ( n20009 , n20005 );
not ( n20010 , n20006 );
and ( n20011 , n20009 , n20010 );
nor ( n20012 , n20008 , n20011 );
not ( n20013 , n20012 );
and ( n20014 , n20013 , n7796 );
not ( n20015 , n20013 );
not ( n20016 , n7795 );
and ( n20017 , n20015 , n20016 );
or ( n20018 , n20014 , n20017 );
buf ( n20019 , n6208 );
buf ( n20020 , n20019 );
not ( n20021 , n20020 );
buf ( n20022 , n6209 );
not ( n20023 , n20022 );
not ( n20024 , n20023 );
or ( n20025 , n20021 , n20024 );
not ( n20026 , n20019 );
buf ( n20027 , n20022 );
nand ( n20028 , n20026 , n20027 );
nand ( n20029 , n20025 , n20028 );
buf ( n20030 , n6210 );
buf ( n20031 , n20030 );
and ( n20032 , n20029 , n20031 );
not ( n20033 , n20029 );
not ( n20034 , n20030 );
and ( n20035 , n20033 , n20034 );
nor ( n20036 , n20032 , n20035 );
buf ( n20037 , n6211 );
nand ( n20038 , n7981 , n20037 );
buf ( n20039 , n6212 );
not ( n20040 , n20039 );
and ( n20041 , n20038 , n20040 );
not ( n20042 , n20038 );
buf ( n20043 , n20039 );
and ( n20044 , n20042 , n20043 );
nor ( n20045 , n20041 , n20044 );
xor ( n20046 , n20036 , n20045 );
buf ( n20047 , n6213 );
nand ( n20048 , n6608 , n20047 );
buf ( n20049 , n6214 );
not ( n20050 , n20049 );
and ( n20051 , n20048 , n20050 );
not ( n20052 , n20048 );
buf ( n20053 , n20049 );
and ( n20054 , n20052 , n20053 );
nor ( n20055 , n20051 , n20054 );
xnor ( n20056 , n20046 , n20055 );
buf ( n20057 , n20056 );
not ( n20058 , n20057 );
buf ( n20059 , n20058 );
and ( n20060 , n20018 , n20059 );
not ( n20061 , n20018 );
not ( n20062 , n20056 );
not ( n20063 , n20062 );
not ( n20064 , n20063 );
not ( n20065 , n20064 );
and ( n20066 , n20061 , n20065 );
nor ( n20067 , n20060 , n20066 );
not ( n20068 , n20067 );
buf ( n20069 , n6215 );
xor ( n20070 , n20069 , n14820 );
buf ( n20071 , n6216 );
nand ( n20072 , n7865 , n20071 );
buf ( n20073 , n6217 );
not ( n20074 , n20073 );
and ( n20075 , n20072 , n20074 );
not ( n20076 , n20072 );
buf ( n20077 , n20073 );
and ( n20078 , n20076 , n20077 );
nor ( n20079 , n20075 , n20078 );
xnor ( n20080 , n20070 , n20079 );
not ( n20081 , n20080 );
buf ( n20082 , n6218 );
not ( n20083 , n20082 );
buf ( n20084 , n6219 );
buf ( n20085 , n20084 );
and ( n20086 , n20083 , n20085 );
not ( n20087 , n20083 );
not ( n20088 , n20084 );
and ( n20089 , n20087 , n20088 );
nor ( n20090 , n20086 , n20089 );
not ( n20091 , n20090 );
and ( n20092 , n20081 , n20091 );
and ( n20093 , n20080 , n20090 );
nor ( n20094 , n20092 , n20093 );
buf ( n20095 , n20094 );
xor ( n20096 , n14934 , n20095 );
buf ( n20097 , n6220 );
not ( n20098 , n20097 );
buf ( n20099 , n6221 );
buf ( n20100 , n20099 );
nand ( n20101 , n20098 , n20100 );
not ( n20102 , n20099 );
buf ( n20103 , n20097 );
nand ( n20104 , n20102 , n20103 );
and ( n20105 , n20101 , n20104 );
xor ( n20106 , n12281 , n20105 );
buf ( n20107 , n6222 );
buf ( n20108 , n6223 );
xor ( n20109 , n20107 , n20108 );
buf ( n20110 , n6224 );
nand ( n20111 , n9159 , n20110 );
xnor ( n20112 , n20109 , n20111 );
xor ( n20113 , n20106 , n20112 );
and ( n20114 , n20096 , n20113 );
not ( n20115 , n20096 );
xor ( n20116 , n12281 , n20105 );
xnor ( n20117 , n20116 , n20112 );
buf ( n20118 , n20117 );
and ( n20119 , n20115 , n20118 );
nor ( n20120 , n20114 , n20119 );
not ( n20121 , n20120 );
nand ( n20122 , n20068 , n20121 );
buf ( n20123 , n6225 );
nand ( n20124 , n7909 , n20123 );
buf ( n20125 , n6226 );
buf ( n20126 , n20125 );
and ( n20127 , n20124 , n20126 );
not ( n20128 , n20124 );
not ( n20129 , n20125 );
and ( n20130 , n20128 , n20129 );
nor ( n20131 , n20127 , n20130 );
not ( n20132 , n20131 );
buf ( n20133 , n10131 );
xor ( n20134 , n10163 , n20133 );
xnor ( n20135 , n20134 , n10141 );
buf ( n20136 , n20135 );
not ( n20137 , n20136 );
or ( n20138 , n20132 , n20137 );
or ( n20139 , n20136 , n20131 );
nand ( n20140 , n20138 , n20139 );
not ( n20141 , n17534 );
not ( n20142 , n20141 );
and ( n20143 , n20140 , n20142 );
not ( n20144 , n20140 );
not ( n20145 , n20142 );
and ( n20146 , n20144 , n20145 );
nor ( n20147 , n20143 , n20146 );
and ( n20148 , n20122 , n20147 );
not ( n20149 , n20122 );
not ( n20150 , n20147 );
and ( n20151 , n20149 , n20150 );
nor ( n20152 , n20148 , n20151 );
not ( n20153 , n20152 );
buf ( n20154 , n6227 );
buf ( n20155 , n20154 );
not ( n20156 , n20155 );
not ( n20157 , n9790 );
not ( n20158 , n20157 );
or ( n20159 , n20156 , n20158 );
not ( n20160 , n20154 );
nand ( n20161 , n20160 , n9791 );
nand ( n20162 , n20159 , n20161 );
buf ( n20163 , n6228 );
not ( n20164 , n20163 );
and ( n20165 , n20162 , n20164 );
not ( n20166 , n20162 );
buf ( n20167 , n20163 );
and ( n20168 , n20166 , n20167 );
nor ( n20169 , n20165 , n20168 );
buf ( n20170 , n6229 );
nand ( n20171 , n7288 , n20170 );
buf ( n20172 , n6230 );
buf ( n20173 , n20172 );
and ( n20174 , n20171 , n20173 );
not ( n20175 , n20171 );
not ( n20176 , n20172 );
and ( n20177 , n20175 , n20176 );
nor ( n20178 , n20174 , n20177 );
xor ( n20179 , n20169 , n20178 );
xor ( n20180 , n20179 , n8720 );
xor ( n20181 , n19083 , n20180 );
buf ( n20182 , n6231 );
nand ( n20183 , n6863 , n20182 );
buf ( n20184 , n6232 );
buf ( n20185 , n20184 );
and ( n20186 , n20183 , n20185 );
not ( n20187 , n20183 );
not ( n20188 , n20184 );
and ( n20189 , n20187 , n20188 );
nor ( n20190 , n20186 , n20189 );
xor ( n20191 , n19588 , n20190 );
buf ( n20192 , n6233 );
nand ( n20193 , n6608 , n20192 );
buf ( n20194 , n6234 );
not ( n20195 , n20194 );
and ( n20196 , n20193 , n20195 );
not ( n20197 , n20193 );
buf ( n20198 , n20194 );
and ( n20199 , n20197 , n20198 );
nor ( n20200 , n20196 , n20199 );
xnor ( n20201 , n20191 , n20200 );
not ( n20202 , n20201 );
buf ( n20203 , n6235 );
buf ( n20204 , n20203 );
not ( n20205 , n20204 );
buf ( n20206 , n6236 );
not ( n20207 , n20206 );
not ( n20208 , n20207 );
or ( n20209 , n20205 , n20208 );
not ( n20210 , n20203 );
buf ( n20211 , n20206 );
nand ( n20212 , n20210 , n20211 );
nand ( n20213 , n20209 , n20212 );
not ( n20214 , n20213 );
not ( n20215 , n20214 );
and ( n20216 , n20202 , n20215 );
and ( n20217 , n20201 , n20214 );
nor ( n20218 , n20216 , n20217 );
xnor ( n20219 , n20181 , n20218 );
not ( n20220 , n20219 );
not ( n20221 , n18368 );
not ( n20222 , n9597 );
or ( n20223 , n20221 , n20222 );
or ( n20224 , n9597 , n18368 );
nand ( n20225 , n20223 , n20224 );
not ( n20226 , n20225 );
not ( n20227 , n9630 );
and ( n20228 , n20226 , n20227 );
and ( n20229 , n20225 , n9630 );
nor ( n20230 , n20228 , n20229 );
not ( n20231 , n15388 );
not ( n20232 , n13456 );
not ( n20233 , n20232 );
or ( n20234 , n20231 , n20233 );
not ( n20235 , n15388 );
not ( n20236 , n13435 );
xor ( n20237 , n20236 , n13454 );
xnor ( n20238 , n20237 , n13444 );
nand ( n20239 , n20235 , n20238 );
nand ( n20240 , n20234 , n20239 );
buf ( n20241 , n6237 );
buf ( n20242 , n20241 );
not ( n20243 , n20242 );
buf ( n20244 , n6238 );
not ( n20245 , n20244 );
not ( n20246 , n20245 );
or ( n20247 , n20243 , n20246 );
not ( n20248 , n20241 );
buf ( n20249 , n20244 );
nand ( n20250 , n20248 , n20249 );
nand ( n20251 , n20247 , n20250 );
buf ( n20252 , n6239 );
not ( n20253 , n20252 );
and ( n20254 , n20251 , n20253 );
not ( n20255 , n20251 );
buf ( n20256 , n20252 );
and ( n20257 , n20255 , n20256 );
nor ( n20258 , n20254 , n20257 );
buf ( n20259 , n6240 );
nand ( n20260 , n6760 , n20259 );
buf ( n20261 , n6241 );
not ( n20262 , n20261 );
and ( n20263 , n20260 , n20262 );
not ( n20264 , n20260 );
buf ( n20265 , n20261 );
and ( n20266 , n20264 , n20265 );
nor ( n20267 , n20263 , n20266 );
xor ( n20268 , n20258 , n20267 );
buf ( n20269 , n6242 );
nand ( n20270 , n7094 , n20269 );
buf ( n20271 , n6243 );
not ( n20272 , n20271 );
and ( n20273 , n20270 , n20272 );
not ( n20274 , n20270 );
buf ( n20275 , n20271 );
and ( n20276 , n20274 , n20275 );
nor ( n20277 , n20273 , n20276 );
xnor ( n20278 , n20268 , n20277 );
not ( n20279 , n20278 );
not ( n20280 , n20279 );
and ( n20281 , n20240 , n20280 );
not ( n20282 , n20240 );
not ( n20283 , n20278 );
buf ( n20284 , n20283 );
and ( n20285 , n20282 , n20284 );
nor ( n20286 , n20281 , n20285 );
nand ( n20287 , n20230 , n20286 );
not ( n20288 , n20287 );
or ( n20289 , n20220 , n20288 );
or ( n20290 , n20287 , n20219 );
nand ( n20291 , n20289 , n20290 );
not ( n20292 , n20291 );
not ( n20293 , n17836 );
not ( n20294 , n20293 );
buf ( n20295 , n6244 );
buf ( n20296 , n20295 );
not ( n20297 , n20296 );
buf ( n20298 , n6245 );
not ( n20299 , n20298 );
not ( n20300 , n20299 );
or ( n20301 , n20297 , n20300 );
not ( n20302 , n20295 );
buf ( n20303 , n20298 );
nand ( n20304 , n20302 , n20303 );
nand ( n20305 , n20301 , n20304 );
and ( n20306 , n20305 , n14608 );
not ( n20307 , n20305 );
not ( n20308 , n14607 );
and ( n20309 , n20307 , n20308 );
nor ( n20310 , n20306 , n20309 );
buf ( n20311 , n6246 );
nand ( n20312 , n10204 , n20311 );
buf ( n20313 , n6247 );
not ( n20314 , n20313 );
and ( n20315 , n20312 , n20314 );
not ( n20316 , n20312 );
buf ( n20317 , n20313 );
and ( n20318 , n20316 , n20317 );
nor ( n20319 , n20315 , n20318 );
xor ( n20320 , n20310 , n20319 );
buf ( n20321 , n6248 );
nand ( n20322 , n7516 , n20321 );
buf ( n20323 , n6249 );
not ( n20324 , n20323 );
and ( n20325 , n20322 , n20324 );
not ( n20326 , n20322 );
buf ( n20327 , n20323 );
and ( n20328 , n20326 , n20327 );
nor ( n20329 , n20325 , n20328 );
xnor ( n20330 , n20320 , n20329 );
not ( n20331 , n20330 );
not ( n20332 , n20331 );
or ( n20333 , n20294 , n20332 );
or ( n20334 , n20331 , n20293 );
nand ( n20335 , n20333 , n20334 );
buf ( n20336 , n6250 );
buf ( n20337 , n20336 );
not ( n20338 , n20337 );
buf ( n20339 , n6251 );
not ( n20340 , n20339 );
not ( n20341 , n20340 );
or ( n20342 , n20338 , n20341 );
not ( n20343 , n20336 );
buf ( n20344 , n20339 );
nand ( n20345 , n20343 , n20344 );
nand ( n20346 , n20342 , n20345 );
buf ( n20347 , n6252 );
buf ( n20348 , n20347 );
and ( n20349 , n20346 , n20348 );
not ( n20350 , n20346 );
not ( n20351 , n20347 );
and ( n20352 , n20350 , n20351 );
nor ( n20353 , n20349 , n20352 );
xor ( n20354 , n20353 , n17711 );
buf ( n20355 , n6253 );
nand ( n20356 , n9619 , n20355 );
buf ( n20357 , n6254 );
not ( n20358 , n20357 );
and ( n20359 , n20356 , n20358 );
not ( n20360 , n20356 );
buf ( n20361 , n20357 );
and ( n20362 , n20360 , n20361 );
nor ( n20363 , n20359 , n20362 );
xnor ( n20364 , n20354 , n20363 );
buf ( n20365 , n20364 );
and ( n20366 , n20335 , n20365 );
not ( n20367 , n20335 );
not ( n20368 , n17711 );
xor ( n20369 , n20353 , n20368 );
xnor ( n20370 , n20369 , n20363 );
not ( n20371 , n20370 );
not ( n20372 , n20371 );
and ( n20373 , n20367 , n20372 );
nor ( n20374 , n20366 , n20373 );
not ( n20375 , n20374 );
buf ( n20376 , n6255 );
nand ( n20377 , n8821 , n20376 );
buf ( n20378 , n6256 );
not ( n20379 , n20378 );
and ( n20380 , n20377 , n20379 );
not ( n20381 , n20377 );
buf ( n20382 , n20378 );
and ( n20383 , n20381 , n20382 );
nor ( n20384 , n20380 , n20383 );
not ( n20385 , n20384 );
not ( n20386 , n11129 );
or ( n20387 , n20385 , n20386 );
not ( n20388 , n20384 );
buf ( n20389 , n11114 );
xor ( n20390 , n20389 , n11124 );
xnor ( n20391 , n20390 , n11128 );
nand ( n20392 , n20388 , n20391 );
nand ( n20393 , n20387 , n20392 );
not ( n20394 , n20131 );
buf ( n20395 , n6257 );
nand ( n20396 , n7230 , n20395 );
buf ( n20397 , n6258 );
not ( n20398 , n20397 );
and ( n20399 , n20396 , n20398 );
not ( n20400 , n20396 );
buf ( n20401 , n20397 );
and ( n20402 , n20400 , n20401 );
nor ( n20403 , n20399 , n20402 );
not ( n20404 , n20403 );
or ( n20405 , n20394 , n20404 );
or ( n20406 , n20131 , n20403 );
nand ( n20407 , n20405 , n20406 );
buf ( n20408 , n6259 );
buf ( n20409 , n20408 );
not ( n20410 , n20409 );
buf ( n20411 , n6260 );
not ( n20412 , n20411 );
not ( n20413 , n20412 );
or ( n20414 , n20410 , n20413 );
not ( n20415 , n20408 );
buf ( n20416 , n20411 );
nand ( n20417 , n20415 , n20416 );
nand ( n20418 , n20414 , n20417 );
buf ( n20419 , n6261 );
buf ( n20420 , n20419 );
and ( n20421 , n20418 , n20420 );
not ( n20422 , n20418 );
not ( n20423 , n20419 );
and ( n20424 , n20422 , n20423 );
nor ( n20425 , n20421 , n20424 );
not ( n20426 , n20425 );
and ( n20427 , n20407 , n20426 );
not ( n20428 , n20407 );
and ( n20429 , n20428 , n20425 );
nor ( n20430 , n20427 , n20429 );
buf ( n20431 , n20430 );
and ( n20432 , n20393 , n20431 );
not ( n20433 , n20393 );
xor ( n20434 , n20425 , n20131 );
buf ( n20435 , n20403 );
xnor ( n20436 , n20434 , n20435 );
buf ( n20437 , n20436 );
and ( n20438 , n20433 , n20437 );
nor ( n20439 , n20432 , n20438 );
nand ( n20440 , n20375 , n20439 );
not ( n20441 , n20440 );
buf ( n20442 , n9470 );
not ( n20443 , n20442 );
not ( n20444 , n19346 );
or ( n20445 , n20443 , n20444 );
not ( n20446 , n20442 );
nand ( n20447 , n20446 , n19342 );
nand ( n20448 , n20445 , n20447 );
and ( n20449 , n20448 , n19349 );
not ( n20450 , n20448 );
not ( n20451 , n19353 );
and ( n20452 , n20450 , n20451 );
nor ( n20453 , n20449 , n20452 );
not ( n20454 , n20453 );
and ( n20455 , n20441 , n20454 );
not ( n20456 , n20374 );
nand ( n20457 , n20456 , n20439 );
and ( n20458 , n20457 , n20453 );
nor ( n20459 , n20455 , n20458 );
not ( n20460 , n20459 );
or ( n20461 , n20292 , n20460 );
or ( n20462 , n20459 , n20291 );
nand ( n20463 , n20461 , n20462 );
buf ( n20464 , n8749 );
buf ( n20465 , n6262 );
buf ( n20466 , n20465 );
not ( n20467 , n20466 );
not ( n20468 , n11110 );
or ( n20469 , n20467 , n20468 );
not ( n20470 , n20465 );
nand ( n20471 , n20470 , n11065 );
nand ( n20472 , n20469 , n20471 );
buf ( n20473 , n6263 );
not ( n20474 , n20473 );
and ( n20475 , n20472 , n20474 );
not ( n20476 , n20472 );
buf ( n20477 , n20473 );
and ( n20478 , n20476 , n20477 );
nor ( n20479 , n20475 , n20478 );
buf ( n20480 , n6264 );
nand ( n20481 , n7299 , n20480 );
buf ( n20482 , n6265 );
buf ( n20483 , n20482 );
and ( n20484 , n20481 , n20483 );
not ( n20485 , n20481 );
not ( n20486 , n20482 );
and ( n20487 , n20485 , n20486 );
nor ( n20488 , n20484 , n20487 );
xor ( n20489 , n20479 , n20488 );
buf ( n20490 , n6266 );
nand ( n20491 , n6660 , n20490 );
buf ( n20492 , n6267 );
buf ( n20493 , n20492 );
and ( n20494 , n20491 , n20493 );
not ( n20495 , n20491 );
not ( n20496 , n20492 );
and ( n20497 , n20495 , n20496 );
nor ( n20498 , n20494 , n20497 );
xnor ( n20499 , n20489 , n20498 );
buf ( n20500 , n20499 );
xor ( n20501 , n20464 , n20500 );
not ( n20502 , n19282 );
xnor ( n20503 , n20501 , n20502 );
buf ( n20504 , n18979 );
buf ( n20505 , n8580 );
and ( n20506 , n20504 , n20505 );
not ( n20507 , n20504 );
and ( n20508 , n20507 , n15850 );
nor ( n20509 , n20506 , n20508 );
not ( n20510 , n20509 );
not ( n20511 , n20510 );
not ( n20512 , n11061 );
or ( n20513 , n20511 , n20512 );
nand ( n20514 , n8612 , n20509 );
nand ( n20515 , n20513 , n20514 );
nand ( n20516 , n20503 , n20515 );
not ( n20517 , n20516 );
buf ( n20518 , n12080 );
not ( n20519 , n20518 );
not ( n20520 , n18045 );
not ( n20521 , n14471 );
not ( n20522 , n20521 );
or ( n20523 , n20520 , n20522 );
not ( n20524 , n18045 );
nand ( n20525 , n20524 , n14471 );
nand ( n20526 , n20523 , n20525 );
not ( n20527 , n20526 );
or ( n20528 , n20519 , n20527 );
or ( n20529 , n20526 , n20518 );
nand ( n20530 , n20528 , n20529 );
not ( n20531 , n20530 );
not ( n20532 , n20531 );
not ( n20533 , n20532 );
and ( n20534 , n20517 , n20533 );
and ( n20535 , n20516 , n20532 );
nor ( n20536 , n20534 , n20535 );
and ( n20537 , n20463 , n20536 );
not ( n20538 , n20463 );
not ( n20539 , n20536 );
and ( n20540 , n20538 , n20539 );
nor ( n20541 , n20537 , n20540 );
not ( n20542 , n16926 );
buf ( n20543 , n6268 );
buf ( n20544 , n6269 );
buf ( n20545 , n20544 );
not ( n20546 , n20545 );
buf ( n20547 , n6270 );
not ( n20548 , n20547 );
not ( n20549 , n20548 );
or ( n20550 , n20546 , n20549 );
not ( n20551 , n20544 );
buf ( n20552 , n20547 );
nand ( n20553 , n20551 , n20552 );
nand ( n20554 , n20550 , n20553 );
xor ( n20555 , n20543 , n20554 );
buf ( n20556 , n6271 );
not ( n20557 , n20556 );
buf ( n20558 , n6272 );
xor ( n20559 , n20557 , n20558 );
buf ( n20560 , n6273 );
nand ( n20561 , n8821 , n20560 );
xnor ( n20562 , n20559 , n20561 );
xnor ( n20563 , n20555 , n20562 );
buf ( n20564 , n20563 );
not ( n20565 , n20564 );
not ( n20566 , n20565 );
or ( n20567 , n20542 , n20566 );
not ( n20568 , n20564 );
or ( n20569 , n20568 , n16926 );
nand ( n20570 , n20567 , n20569 );
and ( n20571 , n20570 , n13500 );
not ( n20572 , n20570 );
and ( n20573 , n20572 , n13499 );
nor ( n20574 , n20571 , n20573 );
not ( n20575 , n20574 );
not ( n20576 , n20575 );
nand ( n20577 , n20067 , n20147 );
not ( n20578 , n20577 );
or ( n20579 , n20576 , n20578 );
or ( n20580 , n20575 , n20577 );
nand ( n20581 , n20579 , n20580 );
not ( n20582 , n20581 );
not ( n20583 , n20582 );
not ( n20584 , n19140 );
xor ( n20585 , n8278 , n20584 );
xor ( n20586 , n20585 , n19658 );
not ( n20587 , n20586 );
buf ( n20588 , n8968 );
and ( n20589 , n8973 , n20588 );
not ( n20590 , n8973 );
and ( n20591 , n20590 , n8969 );
nor ( n20592 , n20589 , n20591 );
not ( n20593 , n20592 );
buf ( n20594 , n6274 );
buf ( n20595 , n20594 );
not ( n20596 , n20595 );
buf ( n20597 , n6275 );
not ( n20598 , n20597 );
not ( n20599 , n20598 );
or ( n20600 , n20596 , n20599 );
not ( n20601 , n20594 );
buf ( n20602 , n20597 );
nand ( n20603 , n20601 , n20602 );
nand ( n20604 , n20600 , n20603 );
buf ( n20605 , n6276 );
not ( n20606 , n20605 );
and ( n20607 , n20604 , n20606 );
not ( n20608 , n20604 );
buf ( n20609 , n20605 );
and ( n20610 , n20608 , n20609 );
nor ( n20611 , n20607 , n20610 );
buf ( n20612 , n6277 );
nand ( n20613 , n8344 , n20612 );
buf ( n20614 , n6278 );
buf ( n20615 , n20614 );
and ( n20616 , n20613 , n20615 );
not ( n20617 , n20613 );
not ( n20618 , n20614 );
and ( n20619 , n20617 , n20618 );
nor ( n20620 , n20616 , n20619 );
xor ( n20621 , n20611 , n20620 );
buf ( n20622 , n6279 );
nand ( n20623 , n9619 , n20622 );
buf ( n20624 , n6280 );
not ( n20625 , n20624 );
and ( n20626 , n20623 , n20625 );
not ( n20627 , n20623 );
buf ( n20628 , n20624 );
and ( n20629 , n20627 , n20628 );
nor ( n20630 , n20626 , n20629 );
xnor ( n20631 , n20621 , n20630 );
not ( n20632 , n20631 );
not ( n20633 , n20632 );
or ( n20634 , n20593 , n20633 );
buf ( n20635 , n20631 );
not ( n20636 , n20635 );
or ( n20637 , n20636 , n20592 );
nand ( n20638 , n20634 , n20637 );
buf ( n20639 , n14337 );
and ( n20640 , n20638 , n20639 );
not ( n20641 , n20638 );
and ( n20642 , n20641 , n14343 );
nor ( n20643 , n20640 , n20642 );
nand ( n20644 , n20587 , n20643 );
not ( n20645 , n18875 );
not ( n20646 , n16420 );
or ( n20647 , n20645 , n20646 );
or ( n20648 , n16420 , n18875 );
nand ( n20649 , n20647 , n20648 );
and ( n20650 , n20649 , n16443 );
not ( n20651 , n20649 );
and ( n20652 , n20651 , n16446 );
nor ( n20653 , n20650 , n20652 );
not ( n20654 , n20653 );
and ( n20655 , n20644 , n20654 );
not ( n20656 , n20644 );
and ( n20657 , n20656 , n20653 );
nor ( n20658 , n20655 , n20657 );
not ( n20659 , n20658 );
or ( n20660 , n20583 , n20659 );
not ( n20661 , n20658 );
nand ( n20662 , n20661 , n20581 );
nand ( n20663 , n20660 , n20662 );
and ( n20664 , n20541 , n20663 );
not ( n20665 , n20541 );
not ( n20666 , n20663 );
and ( n20667 , n20665 , n20666 );
nor ( n20668 , n20664 , n20667 );
not ( n20669 , n20668 );
or ( n20670 , n20153 , n20669 );
not ( n20671 , n20152 );
not ( n20672 , n20541 );
not ( n20673 , n20663 );
and ( n20674 , n20672 , n20673 );
and ( n20675 , n20541 , n20663 );
nor ( n20676 , n20674 , n20675 );
not ( n20677 , n20676 );
nand ( n20678 , n20671 , n20677 );
nand ( n20679 , n20670 , n20678 );
not ( n20680 , n17788 );
not ( n20681 , n12088 );
or ( n20682 , n20680 , n20681 );
not ( n20683 , n17788 );
nand ( n20684 , n20683 , n12018 );
nand ( n20685 , n20682 , n20684 );
not ( n20686 , n14160 );
not ( n20687 , n20686 );
and ( n20688 , n20685 , n20687 );
not ( n20689 , n20685 );
and ( n20690 , n20689 , n20686 );
nor ( n20691 , n20688 , n20690 );
not ( n20692 , n15146 );
not ( n20693 , n17246 );
or ( n20694 , n20692 , n20693 );
or ( n20695 , n17246 , n15146 );
nand ( n20696 , n20694 , n20695 );
not ( n20697 , n14101 );
buf ( n20698 , n20697 );
not ( n20699 , n20698 );
and ( n20700 , n20696 , n20699 );
not ( n20701 , n20696 );
not ( n20702 , n14113 );
not ( n20703 , n20702 );
and ( n20704 , n20701 , n20703 );
nor ( n20705 , n20700 , n20704 );
not ( n20706 , n20705 );
nand ( n20707 , n20691 , n20706 );
not ( n20708 , n20707 );
buf ( n20709 , n6281 );
not ( n20710 , n20709 );
not ( n20711 , n13390 );
or ( n20712 , n20710 , n20711 );
not ( n20713 , n20709 );
nand ( n20714 , n20713 , n13395 );
nand ( n20715 , n20712 , n20714 );
and ( n20716 , n20715 , n13403 );
not ( n20717 , n20715 );
and ( n20718 , n20717 , n11823 );
nor ( n20719 , n20716 , n20718 );
buf ( n20720 , n20719 );
not ( n20721 , n20720 );
and ( n20722 , n20708 , n20721 );
nand ( n20723 , n20691 , n20706 );
and ( n20724 , n20723 , n20720 );
nor ( n20725 , n20722 , n20724 );
buf ( n20726 , n6282 );
buf ( n20727 , n20726 );
not ( n20728 , n20727 );
not ( n20729 , n18554 );
not ( n20730 , n20729 );
or ( n20731 , n20728 , n20730 );
not ( n20732 , n20726 );
nand ( n20733 , n20732 , n18555 );
nand ( n20734 , n20731 , n20733 );
buf ( n20735 , n20734 );
not ( n20736 , n20735 );
buf ( n20737 , n6283 );
buf ( n20738 , n6284 );
not ( n20739 , n20738 );
xor ( n20740 , n20737 , n20739 );
buf ( n20741 , n6285 );
nand ( n20742 , n6934 , n20741 );
buf ( n20743 , n6286 );
not ( n20744 , n20743 );
and ( n20745 , n20742 , n20744 );
not ( n20746 , n20742 );
buf ( n20747 , n20743 );
and ( n20748 , n20746 , n20747 );
nor ( n20749 , n20745 , n20748 );
xnor ( n20750 , n20740 , n20749 );
not ( n20751 , n20750 );
not ( n20752 , n20751 );
or ( n20753 , n20736 , n20752 );
or ( n20754 , n20751 , n20735 );
nand ( n20755 , n20753 , n20754 );
not ( n20756 , n20755 );
buf ( n20757 , n6287 );
buf ( n20758 , n20757 );
not ( n20759 , n20758 );
buf ( n20760 , n6288 );
not ( n20761 , n20760 );
not ( n20762 , n20761 );
or ( n20763 , n20759 , n20762 );
not ( n20764 , n20757 );
buf ( n20765 , n20760 );
nand ( n20766 , n20764 , n20765 );
nand ( n20767 , n20763 , n20766 );
buf ( n20768 , n6289 );
not ( n20769 , n20768 );
and ( n20770 , n20767 , n20769 );
not ( n20771 , n20767 );
buf ( n20772 , n20768 );
and ( n20773 , n20771 , n20772 );
nor ( n20774 , n20770 , n20773 );
buf ( n20775 , n6290 );
nand ( n20776 , n8223 , n20775 );
buf ( n20777 , n6291 );
not ( n20778 , n20777 );
and ( n20779 , n20776 , n20778 );
not ( n20780 , n20776 );
buf ( n20781 , n20777 );
and ( n20782 , n20780 , n20781 );
nor ( n20783 , n20779 , n20782 );
xor ( n20784 , n20774 , n20783 );
buf ( n20785 , n6292 );
nand ( n20786 , n6934 , n20785 );
buf ( n20787 , n6293 );
buf ( n20788 , n20787 );
and ( n20789 , n20786 , n20788 );
not ( n20790 , n20786 );
not ( n20791 , n20787 );
and ( n20792 , n20790 , n20791 );
nor ( n20793 , n20789 , n20792 );
xor ( n20794 , n20784 , n20793 );
not ( n20795 , n20794 );
not ( n20796 , n20795 );
buf ( n20797 , n17630 );
not ( n20798 , n20797 );
and ( n20799 , n20796 , n20798 );
and ( n20800 , n20795 , n20797 );
nor ( n20801 , n20799 , n20800 );
not ( n20802 , n20801 );
and ( n20803 , n20756 , n20802 );
not ( n20804 , n20735 );
not ( n20805 , n20751 );
or ( n20806 , n20804 , n20805 );
not ( n20807 , n20735 );
nand ( n20808 , n20807 , n20750 );
nand ( n20809 , n20806 , n20808 );
and ( n20810 , n20809 , n20801 );
nor ( n20811 , n20803 , n20810 );
not ( n20812 , n20811 );
not ( n20813 , n7686 );
not ( n20814 , n17837 );
or ( n20815 , n20813 , n20814 );
not ( n20816 , n7686 );
nand ( n20817 , n20816 , n17357 );
nand ( n20818 , n20815 , n20817 );
and ( n20819 , n20818 , n17363 );
not ( n20820 , n20818 );
and ( n20821 , n20820 , n17239 );
nor ( n20822 , n20819 , n20821 );
not ( n20823 , n20822 );
nand ( n20824 , n20812 , n20823 );
buf ( n20825 , n14640 );
not ( n20826 , n20825 );
buf ( n20827 , n6294 );
buf ( n20828 , n20827 );
not ( n20829 , n20828 );
buf ( n20830 , n6295 );
not ( n20831 , n20830 );
not ( n20832 , n20831 );
or ( n20833 , n20829 , n20832 );
not ( n20834 , n20827 );
buf ( n20835 , n20830 );
nand ( n20836 , n20834 , n20835 );
nand ( n20837 , n20833 , n20836 );
not ( n20838 , n15143 );
and ( n20839 , n20837 , n20838 );
not ( n20840 , n20837 );
and ( n20841 , n20840 , n15144 );
nor ( n20842 , n20839 , n20841 );
buf ( n20843 , n6296 );
nand ( n20844 , n6660 , n20843 );
buf ( n20845 , n6297 );
buf ( n20846 , n20845 );
and ( n20847 , n20844 , n20846 );
not ( n20848 , n20844 );
not ( n20849 , n20845 );
and ( n20850 , n20848 , n20849 );
nor ( n20851 , n20847 , n20850 );
xor ( n20852 , n20842 , n20851 );
buf ( n20853 , n6298 );
nand ( n20854 , n6934 , n20853 );
buf ( n20855 , n6299 );
not ( n20856 , n20855 );
and ( n20857 , n20854 , n20856 );
not ( n20858 , n20854 );
buf ( n20859 , n20855 );
and ( n20860 , n20858 , n20859 );
nor ( n20861 , n20857 , n20860 );
xor ( n20862 , n20852 , n20861 );
not ( n20863 , n20862 );
not ( n20864 , n20863 );
or ( n20865 , n20826 , n20864 );
not ( n20866 , n20825 );
nand ( n20867 , n20866 , n20862 );
nand ( n20868 , n20865 , n20867 );
not ( n20869 , n16293 );
buf ( n20870 , n6300 );
not ( n20871 , n20870 );
not ( n20872 , n20871 );
or ( n20873 , n20869 , n20872 );
not ( n20874 , n16292 );
buf ( n20875 , n20870 );
nand ( n20876 , n20874 , n20875 );
nand ( n20877 , n20873 , n20876 );
buf ( n20878 , n6301 );
buf ( n20879 , n20878 );
and ( n20880 , n20877 , n20879 );
not ( n20881 , n20877 );
not ( n20882 , n20878 );
and ( n20883 , n20881 , n20882 );
nor ( n20884 , n20880 , n20883 );
buf ( n20885 , n6302 );
nand ( n20886 , n8923 , n20885 );
buf ( n20887 , n6303 );
xor ( n20888 , n20886 , n20887 );
xor ( n20889 , n20884 , n20888 );
buf ( n20890 , n6304 );
nand ( n20891 , n10577 , n20890 );
buf ( n20892 , n6305 );
not ( n20893 , n20892 );
and ( n20894 , n20891 , n20893 );
not ( n20895 , n20891 );
buf ( n20896 , n20892 );
and ( n20897 , n20895 , n20896 );
nor ( n20898 , n20894 , n20897 );
xor ( n20899 , n20889 , n20898 );
buf ( n20900 , n20899 );
and ( n20901 , n20868 , n20900 );
not ( n20902 , n20868 );
xor ( n20903 , n20884 , n20888 );
xnor ( n20904 , n20903 , n20898 );
buf ( n20905 , n20904 );
and ( n20906 , n20902 , n20905 );
nor ( n20907 , n20901 , n20906 );
and ( n20908 , n20824 , n20907 );
not ( n20909 , n20824 );
not ( n20910 , n20907 );
and ( n20911 , n20909 , n20910 );
nor ( n20912 , n20908 , n20911 );
or ( n20913 , n20725 , n20912 );
nand ( n20914 , n20912 , n20725 );
nand ( n20915 , n20913 , n20914 );
xor ( n20916 , n10483 , n14056 );
xnor ( n20917 , n20916 , n8074 );
not ( n20918 , n20917 );
not ( n20919 , n9855 );
not ( n20920 , n20919 );
xor ( n20921 , n7807 , n20920 );
buf ( n20922 , n6306 );
buf ( n20923 , n6307 );
buf ( n20924 , n20923 );
not ( n20925 , n20924 );
not ( n20926 , n9398 );
or ( n20927 , n20925 , n20926 );
not ( n20928 , n20923 );
nand ( n20929 , n20928 , n9353 );
nand ( n20930 , n20927 , n20929 );
xor ( n20931 , n20922 , n20930 );
buf ( n20932 , n6308 );
buf ( n20933 , n6309 );
not ( n20934 , n20933 );
xor ( n20935 , n20932 , n20934 );
buf ( n20936 , n6310 );
nand ( n20937 , n7413 , n20936 );
xnor ( n20938 , n20935 , n20937 );
xnor ( n20939 , n20931 , n20938 );
buf ( n20940 , n20939 );
not ( n20941 , n20940 );
xnor ( n20942 , n20921 , n20941 );
nand ( n20943 , n20918 , n20942 );
not ( n20944 , n20943 );
not ( n20945 , n16446 );
buf ( n20946 , n18896 );
and ( n20947 , n20946 , n16420 );
not ( n20948 , n20946 );
not ( n20949 , n16420 );
and ( n20950 , n20948 , n20949 );
nor ( n20951 , n20947 , n20950 );
not ( n20952 , n20951 );
or ( n20953 , n20945 , n20952 );
or ( n20954 , n20951 , n16446 );
nand ( n20955 , n20953 , n20954 );
buf ( n20956 , n20955 );
not ( n20957 , n20956 );
and ( n20958 , n20944 , n20957 );
and ( n20959 , n20943 , n20956 );
nor ( n20960 , n20958 , n20959 );
and ( n20961 , n20915 , n20960 );
not ( n20962 , n20915 );
not ( n20963 , n20960 );
and ( n20964 , n20962 , n20963 );
nor ( n20965 , n20961 , n20964 );
not ( n20966 , n20965 );
not ( n20967 , n8976 );
not ( n20968 , n20967 );
not ( n20969 , n20968 );
not ( n20970 , n12291 );
not ( n20971 , n8945 );
not ( n20972 , n20971 );
or ( n20973 , n20970 , n20972 );
or ( n20974 , n8947 , n12291 );
nand ( n20975 , n20973 , n20974 );
not ( n20976 , n20975 );
or ( n20977 , n20969 , n20976 );
or ( n20978 , n20975 , n8977 );
nand ( n20979 , n20977 , n20978 );
not ( n20980 , n20979 );
not ( n20981 , n15507 );
xor ( n20982 , n9954 , n20981 );
xor ( n20983 , n20982 , n19889 );
not ( n20984 , n20983 );
nand ( n20985 , n20980 , n20984 );
not ( n20986 , n20985 );
buf ( n20987 , n6311 );
nand ( n20988 , n7515 , n20987 );
buf ( n20989 , n6312 );
buf ( n20990 , n20989 );
and ( n20991 , n20988 , n20990 );
not ( n20992 , n20988 );
not ( n20993 , n20989 );
and ( n20994 , n20992 , n20993 );
nor ( n20995 , n20991 , n20994 );
not ( n20996 , n20995 );
not ( n20997 , n20996 );
not ( n20998 , n13863 );
buf ( n20999 , n6313 );
not ( n21000 , n20999 );
not ( n21001 , n21000 );
or ( n21002 , n20998 , n21001 );
not ( n21003 , n13862 );
buf ( n21004 , n20999 );
nand ( n21005 , n21003 , n21004 );
nand ( n21006 , n21002 , n21005 );
buf ( n21007 , n6314 );
not ( n21008 , n21007 );
and ( n21009 , n21006 , n21008 );
not ( n21010 , n21006 );
buf ( n21011 , n21007 );
and ( n21012 , n21010 , n21011 );
nor ( n21013 , n21009 , n21012 );
xor ( n21014 , n21013 , n15048 );
buf ( n21015 , n6315 );
nand ( n21016 , n7134 , n21015 );
buf ( n21017 , n6316 );
not ( n21018 , n21017 );
and ( n21019 , n21016 , n21018 );
not ( n21020 , n21016 );
buf ( n21021 , n21017 );
and ( n21022 , n21020 , n21021 );
nor ( n21023 , n21019 , n21022 );
xnor ( n21024 , n21014 , n21023 );
not ( n21025 , n21024 );
not ( n21026 , n21025 );
not ( n21027 , n21026 );
or ( n21028 , n20997 , n21027 );
not ( n21029 , n20996 );
buf ( n21030 , n21024 );
not ( n21031 , n21030 );
nand ( n21032 , n21029 , n21031 );
nand ( n21033 , n21028 , n21032 );
not ( n21034 , n7425 );
and ( n21035 , n21033 , n21034 );
not ( n21036 , n21033 );
buf ( n21037 , n7428 );
and ( n21038 , n21036 , n21037 );
nor ( n21039 , n21035 , n21038 );
not ( n21040 , n21039 );
and ( n21041 , n20986 , n21040 );
buf ( n21042 , n20979 );
not ( n21043 , n21042 );
nand ( n21044 , n21043 , n20984 );
and ( n21045 , n21044 , n21039 );
nor ( n21046 , n21041 , n21045 );
not ( n21047 , n21046 );
xor ( n21048 , n8851 , n10463 );
not ( n21049 , n11185 );
xnor ( n21050 , n21048 , n21049 );
not ( n21051 , n21050 );
not ( n21052 , n7278 );
not ( n21053 , n18187 );
or ( n21054 , n21052 , n21053 );
xor ( n21055 , n18166 , n18175 );
xnor ( n21056 , n21055 , n18186 );
buf ( n21057 , n21056 );
nand ( n21058 , n21057 , n7274 );
nand ( n21059 , n21054 , n21058 );
buf ( n21060 , n6317 );
buf ( n21061 , n21060 );
not ( n21062 , n21061 );
not ( n21063 , n6782 );
not ( n21064 , n21063 );
or ( n21065 , n21062 , n21064 );
not ( n21066 , n21060 );
nand ( n21067 , n21066 , n6783 );
nand ( n21068 , n21065 , n21067 );
buf ( n21069 , n6318 );
not ( n21070 , n21069 );
and ( n21071 , n21068 , n21070 );
not ( n21072 , n21068 );
buf ( n21073 , n21069 );
and ( n21074 , n21072 , n21073 );
nor ( n21075 , n21071 , n21074 );
buf ( n21076 , n6319 );
nand ( n21077 , n6905 , n21076 );
buf ( n21078 , n6320 );
buf ( n21079 , n21078 );
and ( n21080 , n21077 , n21079 );
not ( n21081 , n21077 );
not ( n21082 , n21078 );
and ( n21083 , n21081 , n21082 );
nor ( n21084 , n21080 , n21083 );
xor ( n21085 , n21075 , n21084 );
buf ( n21086 , n6321 );
nand ( n21087 , n6816 , n21086 );
buf ( n21088 , n6322 );
buf ( n21089 , n21088 );
and ( n21090 , n21087 , n21089 );
not ( n21091 , n21087 );
not ( n21092 , n21088 );
and ( n21093 , n21091 , n21092 );
nor ( n21094 , n21090 , n21093 );
not ( n21095 , n21094 );
xor ( n21096 , n21085 , n21095 );
not ( n21097 , n21096 );
not ( n21098 , n21097 );
and ( n21099 , n21059 , n21098 );
not ( n21100 , n21059 );
xor ( n21101 , n21075 , n21094 );
not ( n21102 , n21084 );
xnor ( n21103 , n21101 , n21102 );
buf ( n21104 , n21103 );
buf ( n21105 , n21104 );
and ( n21106 , n21100 , n21105 );
nor ( n21107 , n21099 , n21106 );
not ( n21108 , n21107 );
nand ( n21109 , n21051 , n21108 );
buf ( n21110 , n6323 );
nand ( n21111 , n10577 , n21110 );
buf ( n21112 , n6324 );
not ( n21113 , n21112 );
and ( n21114 , n21111 , n21113 );
not ( n21115 , n21111 );
buf ( n21116 , n21112 );
and ( n21117 , n21115 , n21116 );
nor ( n21118 , n21114 , n21117 );
not ( n21119 , n10273 );
xor ( n21120 , n21118 , n21119 );
xnor ( n21121 , n21120 , n10237 );
not ( n21122 , n21121 );
and ( n21123 , n21109 , n21122 );
not ( n21124 , n21109 );
and ( n21125 , n21124 , n21121 );
nor ( n21126 , n21123 , n21125 );
not ( n21127 , n21126 );
or ( n21128 , n21047 , n21127 );
or ( n21129 , n21046 , n21126 );
nand ( n21130 , n21128 , n21129 );
not ( n21131 , n21130 );
and ( n21132 , n20966 , n21131 );
and ( n21133 , n20965 , n21130 );
nor ( n21134 , n21132 , n21133 );
not ( n21135 , n21134 );
not ( n21136 , n21135 );
and ( n21137 , n20679 , n21136 );
not ( n21138 , n20679 );
buf ( n21139 , n21134 );
not ( n21140 , n21139 );
and ( n21141 , n21138 , n21140 );
nor ( n21142 , n21137 , n21141 );
not ( n21143 , n17177 );
buf ( n21144 , n17037 );
not ( n21145 , n21144 );
or ( n21146 , n21143 , n21145 );
nand ( n21147 , n17044 , n17173 );
nand ( n21148 , n21146 , n21147 );
not ( n21149 , n10852 );
buf ( n21150 , n6325 );
not ( n21151 , n21150 );
not ( n21152 , n21151 );
or ( n21153 , n21149 , n21152 );
not ( n21154 , n10851 );
buf ( n21155 , n21150 );
nand ( n21156 , n21154 , n21155 );
nand ( n21157 , n21153 , n21156 );
buf ( n21158 , n6326 );
not ( n21159 , n21158 );
and ( n21160 , n21157 , n21159 );
not ( n21161 , n21157 );
buf ( n21162 , n21158 );
and ( n21163 , n21161 , n21162 );
nor ( n21164 , n21160 , n21163 );
xor ( n21165 , n21164 , n18013 );
buf ( n21166 , n6327 );
nand ( n21167 , n7471 , n21166 );
buf ( n21168 , n6328 );
not ( n21169 , n21168 );
and ( n21170 , n21167 , n21169 );
not ( n21171 , n21167 );
buf ( n21172 , n21168 );
and ( n21173 , n21171 , n21172 );
nor ( n21174 , n21170 , n21173 );
not ( n21175 , n21174 );
xnor ( n21176 , n21165 , n21175 );
not ( n21177 , n21176 );
not ( n21178 , n21177 );
and ( n21179 , n21148 , n21178 );
not ( n21180 , n21148 );
not ( n21181 , n18013 );
not ( n21182 , n21174 );
or ( n21183 , n21181 , n21182 );
or ( n21184 , n18013 , n21174 );
nand ( n21185 , n21183 , n21184 );
buf ( n21186 , n21164 );
and ( n21187 , n21185 , n21186 );
not ( n21188 , n21185 );
not ( n21189 , n21186 );
and ( n21190 , n21188 , n21189 );
nor ( n21191 , n21187 , n21190 );
not ( n21192 , n21191 );
not ( n21193 , n21192 );
buf ( n21194 , n21193 );
and ( n21195 , n21180 , n21194 );
nor ( n21196 , n21179 , n21195 );
not ( n21197 , n21196 );
not ( n21198 , n12170 );
not ( n21199 , n11038 );
xor ( n21200 , n21199 , n11047 );
xnor ( n21201 , n21200 , n11057 );
not ( n21202 , n21201 );
or ( n21203 , n21198 , n21202 );
nand ( n21204 , n11059 , n12166 );
nand ( n21205 , n21203 , n21204 );
buf ( n21206 , n17441 );
and ( n21207 , n21205 , n21206 );
not ( n21208 , n21205 );
and ( n21209 , n21208 , n19646 );
nor ( n21210 , n21207 , n21209 );
nand ( n21211 , n21197 , n21210 );
not ( n21212 , n21211 );
xor ( n21213 , n9446 , n9456 );
xnor ( n21214 , n21213 , n9466 );
buf ( n21215 , n21214 );
xor ( n21216 , n7005 , n21215 );
xnor ( n21217 , n21216 , n9489 );
not ( n21218 , n21217 );
not ( n21219 , n21218 );
or ( n21220 , n21212 , n21219 );
or ( n21221 , n21218 , n21211 );
nand ( n21222 , n21220 , n21221 );
not ( n21223 , n21222 );
not ( n21224 , n17755 );
not ( n21225 , n12080 );
or ( n21226 , n21224 , n21225 );
buf ( n21227 , n12076 );
nand ( n21228 , n21227 , n17751 );
nand ( n21229 , n21226 , n21228 );
and ( n21230 , n21229 , n12089 );
not ( n21231 , n21229 );
and ( n21232 , n21231 , n12019 );
nor ( n21233 , n21230 , n21232 );
buf ( n21234 , n10048 );
and ( n21235 , n21234 , n7579 );
not ( n21236 , n21234 );
not ( n21237 , n7578 );
and ( n21238 , n21236 , n21237 );
or ( n21239 , n21235 , n21238 );
and ( n21240 , n21239 , n7629 );
not ( n21241 , n21239 );
not ( n21242 , n7629 );
and ( n21243 , n21241 , n21242 );
nor ( n21244 , n21240 , n21243 );
nand ( n21245 , n21233 , n21244 );
and ( n21246 , n9849 , n9404 );
not ( n21247 , n9849 );
and ( n21248 , n21247 , n9403 );
nor ( n21249 , n21246 , n21248 );
not ( n21250 , n21249 );
not ( n21251 , n7715 );
not ( n21252 , n21251 );
and ( n21253 , n21250 , n21252 );
and ( n21254 , n21249 , n7716 );
nor ( n21255 , n21253 , n21254 );
and ( n21256 , n21245 , n21255 );
not ( n21257 , n21245 );
not ( n21258 , n21255 );
and ( n21259 , n21257 , n21258 );
nor ( n21260 , n21256 , n21259 );
not ( n21261 , n21260 );
not ( n21262 , n21261 );
buf ( n21263 , n7747 );
not ( n21264 , n21263 );
not ( n21265 , n7752 );
or ( n21266 , n21264 , n21265 );
or ( n21267 , n7752 , n21263 );
nand ( n21268 , n21266 , n21267 );
and ( n21269 , n15743 , n21268 );
not ( n21270 , n21269 );
or ( n21271 , n21268 , n15743 );
nand ( n21272 , n21270 , n21271 );
not ( n21273 , n15748 );
and ( n21274 , n21272 , n21273 );
not ( n21275 , n21272 );
and ( n21276 , n21275 , n15697 );
nor ( n21277 , n21274 , n21276 );
not ( n21278 , n21277 );
nand ( n21279 , n21217 , n21196 );
not ( n21280 , n21279 );
or ( n21281 , n21278 , n21280 );
not ( n21282 , n21197 );
nand ( n21283 , n21282 , n21217 );
or ( n21284 , n21283 , n21277 );
nand ( n21285 , n21281 , n21284 );
not ( n21286 , n21285 );
or ( n21287 , n21262 , n21286 );
or ( n21288 , n21285 , n21261 );
nand ( n21289 , n21287 , n21288 );
not ( n21290 , n21289 );
not ( n21291 , n15630 );
not ( n21292 , n18723 );
or ( n21293 , n21291 , n21292 );
or ( n21294 , n18723 , n15630 );
nand ( n21295 , n21293 , n21294 );
buf ( n21296 , n17666 );
not ( n21297 , n21296 );
and ( n21298 , n21295 , n21297 );
not ( n21299 , n21295 );
and ( n21300 , n21299 , n21296 );
nor ( n21301 , n21298 , n21300 );
buf ( n21302 , n6329 );
nand ( n21303 , n7515 , n21302 );
buf ( n21304 , n6330 );
buf ( n21305 , n21304 );
and ( n21306 , n21303 , n21305 );
not ( n21307 , n21303 );
not ( n21308 , n21304 );
and ( n21309 , n21307 , n21308 );
nor ( n21310 , n21306 , n21309 );
not ( n21311 , n21310 );
not ( n21312 , n21311 );
not ( n21313 , n21312 );
not ( n21314 , n11821 );
not ( n21315 , n21314 );
or ( n21316 , n21313 , n21315 );
or ( n21317 , n11822 , n21312 );
nand ( n21318 , n21316 , n21317 );
and ( n21319 , n21318 , n11868 );
not ( n21320 , n21318 );
not ( n21321 , n11868 );
and ( n21322 , n21320 , n21321 );
nor ( n21323 , n21319 , n21322 );
nand ( n21324 , n21301 , n21323 );
not ( n21325 , n21324 );
not ( n21326 , n7832 );
not ( n21327 , n20939 );
or ( n21328 , n21326 , n21327 );
or ( n21329 , n20939 , n7832 );
nand ( n21330 , n21328 , n21329 );
and ( n21331 , n21330 , n20920 );
not ( n21332 , n21330 );
buf ( n21333 , n9850 );
and ( n21334 , n21332 , n21333 );
nor ( n21335 , n21331 , n21334 );
not ( n21336 , n21335 );
and ( n21337 , n21325 , n21336 );
and ( n21338 , n21324 , n21335 );
nor ( n21339 , n21337 , n21338 );
not ( n21340 , n21339 );
not ( n21341 , n20835 );
not ( n21342 , n15196 );
xor ( n21343 , n16676 , n21342 );
xnor ( n21344 , n21343 , n15203 );
not ( n21345 , n21344 );
or ( n21346 , n21341 , n21345 );
or ( n21347 , n15204 , n20835 );
nand ( n21348 , n21346 , n21347 );
not ( n21349 , n16295 );
and ( n21350 , n21348 , n21349 );
not ( n21351 , n21348 );
and ( n21352 , n21351 , n16295 );
nor ( n21353 , n21350 , n21352 );
buf ( n21354 , n6331 );
not ( n21355 , n21354 );
xor ( n21356 , n20169 , n8719 );
not ( n21357 , n20178 );
xnor ( n21358 , n21356 , n21357 );
not ( n21359 , n21358 );
or ( n21360 , n21355 , n21359 );
not ( n21361 , n21354 );
nand ( n21362 , n21361 , n20180 );
nand ( n21363 , n21360 , n21362 );
buf ( n21364 , n6332 );
buf ( n21365 , n21364 );
not ( n21366 , n21365 );
buf ( n21367 , n6333 );
not ( n21368 , n21367 );
not ( n21369 , n21368 );
or ( n21370 , n21366 , n21369 );
not ( n21371 , n21364 );
buf ( n21372 , n21367 );
nand ( n21373 , n21371 , n21372 );
nand ( n21374 , n21370 , n21373 );
buf ( n21375 , n6334 );
not ( n21376 , n21375 );
and ( n21377 , n21374 , n21376 );
not ( n21378 , n21374 );
buf ( n21379 , n21375 );
and ( n21380 , n21378 , n21379 );
nor ( n21381 , n21377 , n21380 );
xor ( n21382 , n21381 , n15265 );
buf ( n21383 , n6335 );
nand ( n21384 , n10577 , n21383 );
buf ( n21385 , n6336 );
buf ( n21386 , n21385 );
and ( n21387 , n21384 , n21386 );
not ( n21388 , n21384 );
not ( n21389 , n21385 );
and ( n21390 , n21388 , n21389 );
nor ( n21391 , n21387 , n21390 );
xnor ( n21392 , n21382 , n21391 );
buf ( n21393 , n21392 );
not ( n21394 , n21393 );
and ( n21395 , n21363 , n21394 );
not ( n21396 , n21363 );
not ( n21397 , n21392 );
buf ( n21398 , n21397 );
not ( n21399 , n21398 );
and ( n21400 , n21396 , n21399 );
nor ( n21401 , n21395 , n21400 );
nand ( n21402 , n21353 , n21401 );
buf ( n21403 , n6337 );
buf ( n21404 , n21403 );
not ( n21405 , n21404 );
buf ( n21406 , n6338 );
not ( n21407 , n21406 );
not ( n21408 , n21407 );
or ( n21409 , n21405 , n21408 );
not ( n21410 , n21403 );
buf ( n21411 , n21406 );
nand ( n21412 , n21410 , n21411 );
nand ( n21413 , n21409 , n21412 );
not ( n21414 , n21413 );
not ( n21415 , n21414 );
buf ( n21416 , n6339 );
buf ( n21417 , n6340 );
not ( n21418 , n21417 );
xor ( n21419 , n21416 , n21418 );
buf ( n21420 , n6341 );
nand ( n21421 , n6934 , n21420 );
buf ( n21422 , n6342 );
not ( n21423 , n21422 );
and ( n21424 , n21421 , n21423 );
not ( n21425 , n21421 );
buf ( n21426 , n21422 );
and ( n21427 , n21425 , n21426 );
nor ( n21428 , n21424 , n21427 );
xnor ( n21429 , n21419 , n21428 );
not ( n21430 , n21429 );
or ( n21431 , n21415 , n21430 );
or ( n21432 , n21429 , n21414 );
nand ( n21433 , n21431 , n21432 );
not ( n21434 , n21433 );
not ( n21435 , n21434 );
not ( n21436 , n14195 );
not ( n21437 , n21436 );
buf ( n21438 , n6343 );
buf ( n21439 , n21438 );
not ( n21440 , n21439 );
buf ( n21441 , n6344 );
not ( n21442 , n21441 );
not ( n21443 , n21442 );
or ( n21444 , n21440 , n21443 );
not ( n21445 , n21438 );
buf ( n21446 , n21441 );
nand ( n21447 , n21445 , n21446 );
nand ( n21448 , n21444 , n21447 );
buf ( n21449 , n6345 );
buf ( n21450 , n21449 );
and ( n21451 , n21448 , n21450 );
not ( n21452 , n21448 );
not ( n21453 , n21449 );
and ( n21454 , n21452 , n21453 );
nor ( n21455 , n21451 , n21454 );
xor ( n21456 , n21455 , n20012 );
buf ( n21457 , n6346 );
nand ( n21458 , n8387 , n21457 );
buf ( n21459 , n6347 );
buf ( n21460 , n21459 );
and ( n21461 , n21458 , n21460 );
not ( n21462 , n21458 );
not ( n21463 , n21459 );
and ( n21464 , n21462 , n21463 );
nor ( n21465 , n21461 , n21464 );
not ( n21466 , n21465 );
xor ( n21467 , n21456 , n21466 );
not ( n21468 , n21467 );
or ( n21469 , n21437 , n21468 );
xor ( n21470 , n21455 , n21465 );
xnor ( n21471 , n21470 , n20013 );
nand ( n21472 , n21471 , n14195 );
nand ( n21473 , n21469 , n21472 );
not ( n21474 , n21473 );
and ( n21475 , n21435 , n21474 );
and ( n21476 , n21434 , n21473 );
nor ( n21477 , n21475 , n21476 );
and ( n21478 , n21402 , n21477 );
not ( n21479 , n21402 );
not ( n21480 , n21477 );
and ( n21481 , n21479 , n21480 );
nor ( n21482 , n21478 , n21481 );
not ( n21483 , n21482 );
or ( n21484 , n21340 , n21483 );
or ( n21485 , n21482 , n21339 );
nand ( n21486 , n21484 , n21485 );
buf ( n21487 , n8175 );
not ( n21488 , n21487 );
buf ( n21489 , n6348 );
buf ( n21490 , n6349 );
not ( n21491 , n21490 );
buf ( n21492 , n6350 );
buf ( n21493 , n21492 );
nand ( n21494 , n21491 , n21493 );
not ( n21495 , n21492 );
buf ( n21496 , n21490 );
nand ( n21497 , n21495 , n21496 );
and ( n21498 , n21494 , n21497 );
xor ( n21499 , n21489 , n21498 );
not ( n21500 , n15079 );
buf ( n21501 , n6351 );
nand ( n21502 , n6760 , n21501 );
buf ( n21503 , n6352 );
not ( n21504 , n21503 );
and ( n21505 , n21502 , n21504 );
not ( n21506 , n21502 );
buf ( n21507 , n21503 );
and ( n21508 , n21506 , n21507 );
nor ( n21509 , n21505 , n21508 );
not ( n21510 , n21509 );
or ( n21511 , n21500 , n21510 );
or ( n21512 , n15079 , n21509 );
nand ( n21513 , n21511 , n21512 );
xnor ( n21514 , n21499 , n21513 );
buf ( n21515 , n21514 );
not ( n21516 , n21515 );
or ( n21517 , n21488 , n21516 );
or ( n21518 , n21515 , n21487 );
nand ( n21519 , n21517 , n21518 );
not ( n21520 , n16555 );
buf ( n21521 , n21520 );
not ( n21522 , n21521 );
not ( n21523 , n21522 );
and ( n21524 , n21519 , n21523 );
not ( n21525 , n21519 );
and ( n21526 , n21525 , n21522 );
nor ( n21527 , n21524 , n21526 );
not ( n21528 , n17591 );
not ( n21529 , n21528 );
not ( n21530 , n19952 );
not ( n21531 , n10463 );
or ( n21532 , n21530 , n21531 );
or ( n21533 , n10463 , n19952 );
nand ( n21534 , n21532 , n21533 );
not ( n21535 , n21534 );
or ( n21536 , n21529 , n21535 );
or ( n21537 , n21534 , n21528 );
nand ( n21538 , n21536 , n21537 );
nand ( n21539 , n21527 , n21538 );
not ( n21540 , n12580 );
not ( n21541 , n15995 );
not ( n21542 , n19686 );
or ( n21543 , n21541 , n21542 );
not ( n21544 , n15994 );
nand ( n21545 , n21544 , n19682 );
nand ( n21546 , n21543 , n21545 );
not ( n21547 , n11263 );
and ( n21548 , n21546 , n21547 );
not ( n21549 , n21546 );
and ( n21550 , n21549 , n11264 );
nor ( n21551 , n21548 , n21550 );
buf ( n21552 , n6353 );
nand ( n21553 , n7412 , n21552 );
buf ( n21554 , n6354 );
buf ( n21555 , n21554 );
and ( n21556 , n21553 , n21555 );
not ( n21557 , n21553 );
not ( n21558 , n21554 );
and ( n21559 , n21557 , n21558 );
nor ( n21560 , n21556 , n21559 );
xor ( n21561 , n21551 , n21560 );
buf ( n21562 , n6355 );
nand ( n21563 , n9257 , n21562 );
buf ( n21564 , n6356 );
not ( n21565 , n21564 );
and ( n21566 , n21563 , n21565 );
not ( n21567 , n21563 );
buf ( n21568 , n21564 );
and ( n21569 , n21567 , n21568 );
nor ( n21570 , n21566 , n21569 );
xnor ( n21571 , n21561 , n21570 );
buf ( n21572 , n21571 );
not ( n21573 , n21572 );
or ( n21574 , n21540 , n21573 );
not ( n21575 , n12580 );
not ( n21576 , n21571 );
buf ( n21577 , n21576 );
nand ( n21578 , n21575 , n21577 );
nand ( n21579 , n21574 , n21578 );
not ( n21580 , n7886 );
and ( n21581 , n21579 , n21580 );
not ( n21582 , n21579 );
buf ( n21583 , n7886 );
and ( n21584 , n21582 , n21583 );
nor ( n21585 , n21581 , n21584 );
not ( n21586 , n21585 );
and ( n21587 , n21539 , n21586 );
not ( n21588 , n21539 );
and ( n21589 , n21588 , n21585 );
nor ( n21590 , n21587 , n21589 );
not ( n21591 , n21590 );
and ( n21592 , n21486 , n21591 );
not ( n21593 , n21486 );
and ( n21594 , n21593 , n21590 );
nor ( n21595 , n21592 , n21594 );
not ( n21596 , n21595 );
or ( n21597 , n21290 , n21596 );
not ( n21598 , n21595 );
not ( n21599 , n21289 );
nand ( n21600 , n21598 , n21599 );
nand ( n21601 , n21597 , n21600 );
not ( n21602 , n21601 );
not ( n21603 , n21602 );
or ( n21604 , n21223 , n21603 );
not ( n21605 , n21222 );
nand ( n21606 , n21605 , n21601 );
nand ( n21607 , n21604 , n21606 );
not ( n21608 , n16426 );
not ( n21609 , n10587 );
or ( n21610 , n21608 , n21609 );
or ( n21611 , n10587 , n16426 );
nand ( n21612 , n21610 , n21611 );
and ( n21613 , n21612 , n10644 );
not ( n21614 , n21612 );
and ( n21615 , n21614 , n10641 );
nor ( n21616 , n21613 , n21615 );
not ( n21617 , n18084 );
not ( n21618 , n10080 );
buf ( n21619 , n6357 );
buf ( n21620 , n21619 );
not ( n21621 , n21620 );
buf ( n21622 , n6358 );
not ( n21623 , n21622 );
not ( n21624 , n21623 );
or ( n21625 , n21621 , n21624 );
not ( n21626 , n21619 );
buf ( n21627 , n21622 );
nand ( n21628 , n21626 , n21627 );
nand ( n21629 , n21625 , n21628 );
buf ( n21630 , n6359 );
buf ( n21631 , n21630 );
and ( n21632 , n21629 , n21631 );
not ( n21633 , n21629 );
not ( n21634 , n21630 );
and ( n21635 , n21633 , n21634 );
nor ( n21636 , n21632 , n21635 );
buf ( n21637 , n6360 );
nand ( n21638 , n7477 , n21637 );
buf ( n21639 , n6361 );
buf ( n21640 , n21639 );
and ( n21641 , n21638 , n21640 );
not ( n21642 , n21638 );
not ( n21643 , n21639 );
and ( n21644 , n21642 , n21643 );
nor ( n21645 , n21641 , n21644 );
not ( n21646 , n21645 );
xor ( n21647 , n21636 , n21646 );
xnor ( n21648 , n21647 , n19509 );
not ( n21649 , n21648 );
or ( n21650 , n21618 , n21649 );
or ( n21651 , n21648 , n10080 );
nand ( n21652 , n21650 , n21651 );
not ( n21653 , n21652 );
and ( n21654 , n21617 , n21653 );
and ( n21655 , n18084 , n21652 );
nor ( n21656 , n21654 , n21655 );
nand ( n21657 , n21616 , n21656 );
not ( n21658 , n21657 );
not ( n21659 , n20765 );
buf ( n21660 , n6362 );
buf ( n21661 , n21660 );
not ( n21662 , n21661 );
not ( n21663 , n11826 );
or ( n21664 , n21662 , n21663 );
not ( n21665 , n21660 );
nand ( n21666 , n21665 , n11782 );
nand ( n21667 , n21664 , n21666 );
buf ( n21668 , n6363 );
buf ( n21669 , n21668 );
and ( n21670 , n21667 , n21669 );
not ( n21671 , n21667 );
not ( n21672 , n21668 );
and ( n21673 , n21671 , n21672 );
nor ( n21674 , n21670 , n21673 );
not ( n21675 , n21674 );
xor ( n21676 , n21675 , n21310 );
buf ( n21677 , n6364 );
nand ( n21678 , n6706 , n21677 );
buf ( n21679 , n6365 );
buf ( n21680 , n21679 );
and ( n21681 , n21678 , n21680 );
not ( n21682 , n21678 );
not ( n21683 , n21679 );
and ( n21684 , n21682 , n21683 );
nor ( n21685 , n21681 , n21684 );
buf ( n21686 , n21685 );
xnor ( n21687 , n21676 , n21686 );
not ( n21688 , n21687 );
not ( n21689 , n21688 );
or ( n21690 , n21659 , n21689 );
not ( n21691 , n20765 );
nand ( n21692 , n21691 , n21687 );
nand ( n21693 , n21690 , n21692 );
not ( n21694 , n18594 );
and ( n21695 , n21693 , n21694 );
not ( n21696 , n21693 );
and ( n21697 , n21696 , n18594 );
nor ( n21698 , n21695 , n21697 );
not ( n21699 , n21698 );
and ( n21700 , n21658 , n21699 );
and ( n21701 , n21657 , n21698 );
nor ( n21702 , n21700 , n21701 );
not ( n21703 , n21702 );
not ( n21704 , n20095 );
nor ( n21705 , n18644 , n14974 );
not ( n21706 , n21705 );
nand ( n21707 , n18644 , n14974 );
nand ( n21708 , n21706 , n21707 );
not ( n21709 , n21708 );
and ( n21710 , n21704 , n21709 );
and ( n21711 , n20095 , n21708 );
nor ( n21712 , n21710 , n21711 );
not ( n21713 , n17119 );
not ( n21714 , n21571 );
or ( n21715 , n21713 , n21714 );
or ( n21716 , n21571 , n17119 );
nand ( n21717 , n21715 , n21716 );
not ( n21718 , n21717 );
not ( n21719 , n21718 );
not ( n21720 , n21580 );
or ( n21721 , n21719 , n21720 );
nand ( n21722 , n7886 , n21717 );
nand ( n21723 , n21721 , n21722 );
nand ( n21724 , n21712 , n21723 );
not ( n21725 , n16689 );
buf ( n21726 , n6366 );
buf ( n21727 , n6367 );
buf ( n21728 , n21727 );
and ( n21729 , n11010 , n21728 );
not ( n21730 , n11010 );
not ( n21731 , n21727 );
and ( n21732 , n21730 , n21731 );
nor ( n21733 , n21729 , n21732 );
xor ( n21734 , n21726 , n21733 );
buf ( n21735 , n6368 );
buf ( n21736 , n6369 );
xor ( n21737 , n21735 , n21736 );
buf ( n21738 , n6370 );
nand ( n21739 , n7478 , n21738 );
xnor ( n21740 , n21737 , n21739 );
xnor ( n21741 , n21734 , n21740 );
not ( n21742 , n21741 );
not ( n21743 , n21742 );
or ( n21744 , n21725 , n21743 );
or ( n21745 , n21742 , n16689 );
nand ( n21746 , n21744 , n21745 );
buf ( n21747 , n6371 );
buf ( n21748 , n6372 );
nand ( n21749 , n8134 , n21748 );
buf ( n21750 , n6373 );
buf ( n21751 , n21750 );
and ( n21752 , n21749 , n21751 );
not ( n21753 , n21749 );
not ( n21754 , n21750 );
and ( n21755 , n21753 , n21754 );
nor ( n21756 , n21752 , n21755 );
xor ( n21757 , n21747 , n21756 );
buf ( n21758 , n6374 );
nand ( n21759 , n7515 , n21758 );
buf ( n21760 , n6375 );
not ( n21761 , n21760 );
and ( n21762 , n21759 , n21761 );
not ( n21763 , n21759 );
buf ( n21764 , n21760 );
and ( n21765 , n21763 , n21764 );
nor ( n21766 , n21762 , n21765 );
xnor ( n21767 , n21757 , n21766 );
not ( n21768 , n21767 );
buf ( n21769 , n6376 );
not ( n21770 , n21769 );
and ( n21771 , n21770 , n9978 );
not ( n21772 , n21770 );
not ( n21773 , n9977 );
and ( n21774 , n21772 , n21773 );
nor ( n21775 , n21771 , n21774 );
not ( n21776 , n21775 );
and ( n21777 , n21768 , n21776 );
and ( n21778 , n21767 , n21775 );
nor ( n21779 , n21777 , n21778 );
buf ( n21780 , n21779 );
and ( n21781 , n21746 , n21780 );
not ( n21782 , n21746 );
not ( n21783 , n21779 );
and ( n21784 , n21782 , n21783 );
nor ( n21785 , n21781 , n21784 );
and ( n21786 , n21724 , n21785 );
not ( n21787 , n21724 );
not ( n21788 , n21785 );
and ( n21789 , n21787 , n21788 );
nor ( n21790 , n21786 , n21789 );
not ( n21791 , n21790 );
or ( n21792 , n21703 , n21791 );
or ( n21793 , n21790 , n21702 );
nand ( n21794 , n21792 , n21793 );
buf ( n21795 , n6377 );
not ( n21796 , n21795 );
not ( n21797 , n21796 );
not ( n21798 , n15395 );
or ( n21799 , n21797 , n21798 );
not ( n21800 , n21796 );
nand ( n21801 , n21800 , n18680 );
nand ( n21802 , n21799 , n21801 );
and ( n21803 , n21802 , n18730 );
not ( n21804 , n21802 );
and ( n21805 , n21804 , n18724 );
nor ( n21806 , n21803 , n21805 );
not ( n21807 , n21806 );
not ( n21808 , n14624 );
not ( n21809 , n20862 );
not ( n21810 , n21809 );
or ( n21811 , n21808 , n21810 );
not ( n21812 , n20862 );
or ( n21813 , n21812 , n14624 );
nand ( n21814 , n21811 , n21813 );
and ( n21815 , n21814 , n20900 );
not ( n21816 , n21814 );
and ( n21817 , n21816 , n20905 );
nor ( n21818 , n21815 , n21817 );
not ( n21819 , n21818 );
nand ( n21820 , n21807 , n21819 );
not ( n21821 , n20552 );
xor ( n21822 , n11696 , n11705 );
xnor ( n21823 , n21822 , n11715 );
not ( n21824 , n21823 );
or ( n21825 , n21821 , n21824 );
or ( n21826 , n11716 , n20552 );
nand ( n21827 , n21825 , n21826 );
buf ( n21828 , n11425 );
and ( n21829 , n21827 , n21828 );
not ( n21830 , n21827 );
xor ( n21831 , n11404 , n11423 );
xnor ( n21832 , n21831 , n18094 );
not ( n21833 , n21832 );
not ( n21834 , n21833 );
and ( n21835 , n21830 , n21834 );
nor ( n21836 , n21829 , n21835 );
xor ( n21837 , n21820 , n21836 );
and ( n21838 , n21794 , n21837 );
not ( n21839 , n21794 );
not ( n21840 , n21837 );
and ( n21841 , n21839 , n21840 );
nor ( n21842 , n21838 , n21841 );
buf ( n21843 , n21842 );
not ( n21844 , n13760 );
buf ( n21845 , n6378 );
buf ( n21846 , n21845 );
not ( n21847 , n21846 );
buf ( n21848 , n6379 );
not ( n21849 , n21848 );
not ( n21850 , n21849 );
or ( n21851 , n21847 , n21850 );
not ( n21852 , n21845 );
buf ( n21853 , n21848 );
nand ( n21854 , n21852 , n21853 );
nand ( n21855 , n21851 , n21854 );
and ( n21856 , n21855 , n11371 );
not ( n21857 , n21855 );
not ( n21858 , n11370 );
and ( n21859 , n21857 , n21858 );
nor ( n21860 , n21856 , n21859 );
not ( n21861 , n21860 );
xor ( n21862 , n21861 , n9644 );
buf ( n21863 , n6380 );
nand ( n21864 , n7617 , n21863 );
buf ( n21865 , n6381 );
not ( n21866 , n21865 );
and ( n21867 , n21864 , n21866 );
not ( n21868 , n21864 );
buf ( n21869 , n21865 );
and ( n21870 , n21868 , n21869 );
nor ( n21871 , n21867 , n21870 );
xnor ( n21872 , n21862 , n21871 );
buf ( n21873 , n21872 );
not ( n21874 , n21873 );
or ( n21875 , n21844 , n21874 );
or ( n21876 , n21873 , n13760 );
nand ( n21877 , n21875 , n21876 );
not ( n21878 , n19658 );
and ( n21879 , n21877 , n21878 );
not ( n21880 , n21877 );
and ( n21881 , n21880 , n19658 );
nor ( n21882 , n21879 , n21881 );
not ( n21883 , n11545 );
buf ( n21884 , n6382 );
not ( n21885 , n21884 );
not ( n21886 , n21885 );
or ( n21887 , n21883 , n21886 );
not ( n21888 , n11544 );
buf ( n21889 , n21884 );
nand ( n21890 , n21888 , n21889 );
nand ( n21891 , n21887 , n21890 );
buf ( n21892 , n6383 );
buf ( n21893 , n21892 );
and ( n21894 , n21891 , n21893 );
not ( n21895 , n21891 );
not ( n21896 , n21892 );
and ( n21897 , n21895 , n21896 );
nor ( n21898 , n21894 , n21897 );
buf ( n21899 , n6384 );
nand ( n21900 , n7133 , n21899 );
buf ( n21901 , n6385 );
buf ( n21902 , n21901 );
and ( n21903 , n21900 , n21902 );
not ( n21904 , n21900 );
not ( n21905 , n21901 );
and ( n21906 , n21904 , n21905 );
nor ( n21907 , n21903 , n21906 );
xor ( n21908 , n21898 , n21907 );
buf ( n21909 , n6386 );
nand ( n21910 , n7082 , n21909 );
buf ( n21911 , n6387 );
buf ( n21912 , n21911 );
and ( n21913 , n21910 , n21912 );
not ( n21914 , n21910 );
not ( n21915 , n21911 );
and ( n21916 , n21914 , n21915 );
nor ( n21917 , n21913 , n21916 );
xnor ( n21918 , n21908 , n21917 );
not ( n21919 , n21918 );
not ( n21920 , n21919 );
not ( n21921 , n21920 );
not ( n21922 , n7892 );
not ( n21923 , n13026 );
not ( n21924 , n18789 );
or ( n21925 , n21923 , n21924 );
not ( n21926 , n13025 );
nand ( n21927 , n21926 , n18784 );
nand ( n21928 , n21925 , n21927 );
buf ( n21929 , n6388 );
not ( n21930 , n21929 );
and ( n21931 , n21928 , n21930 );
not ( n21932 , n21928 );
buf ( n21933 , n21929 );
and ( n21934 , n21932 , n21933 );
nor ( n21935 , n21931 , n21934 );
buf ( n21936 , n6389 );
nand ( n21937 , n7616 , n21936 );
buf ( n21938 , n6390 );
buf ( n21939 , n21938 );
and ( n21940 , n21937 , n21939 );
not ( n21941 , n21937 );
not ( n21942 , n21938 );
and ( n21943 , n21941 , n21942 );
nor ( n21944 , n21940 , n21943 );
xor ( n21945 , n21935 , n21944 );
buf ( n21946 , n6391 );
nand ( n21947 , n8519 , n21946 );
buf ( n21948 , n6392 );
buf ( n21949 , n21948 );
and ( n21950 , n21947 , n21949 );
not ( n21951 , n21947 );
not ( n21952 , n21948 );
and ( n21953 , n21951 , n21952 );
nor ( n21954 , n21950 , n21953 );
xor ( n21955 , n21945 , n21954 );
not ( n21956 , n21955 );
or ( n21957 , n21922 , n21956 );
xor ( n21958 , n21935 , n21954 );
xor ( n21959 , n21958 , n21944 );
not ( n21960 , n21959 );
not ( n21961 , n21960 );
or ( n21962 , n21961 , n7892 );
nand ( n21963 , n21957 , n21962 );
not ( n21964 , n21963 );
or ( n21965 , n21921 , n21964 );
not ( n21966 , n21919 );
or ( n21967 , n21963 , n21966 );
nand ( n21968 , n21965 , n21967 );
not ( n21969 , n21968 );
nand ( n21970 , n21882 , n21969 );
not ( n21971 , n21970 );
not ( n21972 , n9190 );
not ( n21973 , n13236 );
or ( n21974 , n21972 , n21973 );
or ( n21975 , n13236 , n9190 );
nand ( n21976 , n21974 , n21975 );
not ( n21977 , n6638 );
and ( n21978 , n21976 , n21977 );
not ( n21979 , n21976 );
not ( n21980 , n21977 );
and ( n21981 , n21979 , n21980 );
nor ( n21982 , n21978 , n21981 );
not ( n21983 , n21982 );
not ( n21984 , n21983 );
and ( n21985 , n21971 , n21984 );
and ( n21986 , n21970 , n21983 );
nor ( n21987 , n21985 , n21986 );
buf ( n21988 , n17908 );
xor ( n21989 , n21988 , n19228 );
xnor ( n21990 , n21989 , n19233 );
buf ( n21991 , n21990 );
not ( n21992 , n21991 );
not ( n21993 , n19603 );
and ( n21994 , n21992 , n21993 );
and ( n21995 , n21991 , n19603 );
nor ( n21996 , n21994 , n21995 );
not ( n21997 , n19282 );
and ( n21998 , n21996 , n21997 );
not ( n21999 , n21996 );
not ( n22000 , n20502 );
and ( n22001 , n21999 , n22000 );
nor ( n22002 , n21998 , n22001 );
not ( n22003 , n18391 );
not ( n22004 , n16997 );
or ( n22005 , n22003 , n22004 );
not ( n22006 , n16997 );
nand ( n22007 , n22006 , n18387 );
nand ( n22008 , n22005 , n22007 );
and ( n22009 , n22008 , n17044 );
not ( n22010 , n22008 );
buf ( n22011 , n21144 );
and ( n22012 , n22010 , n22011 );
nor ( n22013 , n22009 , n22012 );
not ( n22014 , n22013 );
nand ( n22015 , n22002 , n22014 );
not ( n22016 , n7756 );
not ( n22017 , n18441 );
not ( n22018 , n12804 );
or ( n22019 , n22017 , n22018 );
or ( n22020 , n12804 , n18441 );
nand ( n22021 , n22019 , n22020 );
not ( n22022 , n22021 );
and ( n22023 , n22016 , n22022 );
and ( n22024 , n7756 , n22021 );
nor ( n22025 , n22023 , n22024 );
and ( n22026 , n22015 , n22025 );
not ( n22027 , n22015 );
not ( n22028 , n22025 );
and ( n22029 , n22027 , n22028 );
nor ( n22030 , n22026 , n22029 );
and ( n22031 , n21987 , n22030 );
not ( n22032 , n21987 );
not ( n22033 , n22030 );
and ( n22034 , n22032 , n22033 );
nor ( n22035 , n22031 , n22034 );
and ( n22036 , n21843 , n22035 );
not ( n22037 , n21843 );
not ( n22038 , n22035 );
and ( n22039 , n22037 , n22038 );
nor ( n22040 , n22036 , n22039 );
buf ( n22041 , n22040 );
and ( n22042 , n21607 , n22041 );
not ( n22043 , n21607 );
not ( n22044 , n22035 );
not ( n22045 , n21842 );
or ( n22046 , n22044 , n22045 );
not ( n22047 , n21842 );
nand ( n22048 , n22047 , n22038 );
nand ( n22049 , n22046 , n22048 );
buf ( n22050 , n22049 );
and ( n22051 , n22043 , n22050 );
nor ( n22052 , n22042 , n22051 );
nand ( n22053 , n21142 , n22052 );
or ( n22054 , n20003 , n22053 );
not ( n22055 , n22052 );
not ( n22056 , n19999 );
or ( n22057 , n22055 , n22056 );
buf ( n22058 , n13752 );
buf ( n22059 , n22058 );
nor ( n22060 , n21142 , n22059 );
nand ( n22061 , n22057 , n22060 );
buf ( n22062 , n13766 );
nand ( n22063 , n22062 , n19092 );
nand ( n22064 , n22054 , n22061 , n22063 );
buf ( n22065 , n22064 );
buf ( n22066 , n22065 );
not ( n22067 , n18780 );
not ( n22068 , n22067 );
buf ( n22069 , n6393 );
buf ( n22070 , n6394 );
buf ( n22071 , n22070 );
not ( n22072 , n22071 );
buf ( n22073 , n6395 );
not ( n22074 , n22073 );
not ( n22075 , n22074 );
or ( n22076 , n22072 , n22075 );
not ( n22077 , n22070 );
buf ( n22078 , n22073 );
nand ( n22079 , n22077 , n22078 );
nand ( n22080 , n22076 , n22079 );
xor ( n22081 , n22069 , n22080 );
buf ( n22082 , n6396 );
not ( n22083 , n22082 );
xor ( n22084 , n21354 , n22083 );
buf ( n22085 , n6397 );
nand ( n22086 , n8134 , n22085 );
xnor ( n22087 , n22084 , n22086 );
xnor ( n22088 , n22081 , n22087 );
not ( n22089 , n22088 );
not ( n22090 , n22089 );
not ( n22091 , n9045 );
and ( n22092 , n22090 , n22091 );
xor ( n22093 , n22069 , n22080 );
xnor ( n22094 , n22093 , n22087 );
not ( n22095 , n22094 );
and ( n22096 , n22095 , n9045 );
nor ( n22097 , n22092 , n22096 );
not ( n22098 , n22097 );
and ( n22099 , n22068 , n22098 );
and ( n22100 , n22067 , n22097 );
nor ( n22101 , n22099 , n22100 );
nand ( n22102 , n22101 , n19695 );
not ( n22103 , n22102 );
not ( n22104 , n11167 );
not ( n22105 , n19192 );
buf ( n22106 , n6398 );
not ( n22107 , n22106 );
not ( n22108 , n22107 );
or ( n22109 , n22105 , n22108 );
not ( n22110 , n19191 );
buf ( n22111 , n22106 );
nand ( n22112 , n22110 , n22111 );
nand ( n22113 , n22109 , n22112 );
buf ( n22114 , n6399 );
buf ( n22115 , n22114 );
and ( n22116 , n22113 , n22115 );
not ( n22117 , n22113 );
not ( n22118 , n22114 );
and ( n22119 , n22117 , n22118 );
nor ( n22120 , n22116 , n22119 );
buf ( n22121 , n6400 );
nand ( n22122 , n7195 , n22121 );
buf ( n22123 , n6401 );
buf ( n22124 , n22123 );
and ( n22125 , n22122 , n22124 );
not ( n22126 , n22122 );
not ( n22127 , n22123 );
and ( n22128 , n22126 , n22127 );
nor ( n22129 , n22125 , n22128 );
xor ( n22130 , n22120 , n22129 );
buf ( n22131 , n6402 );
nand ( n22132 , n13379 , n22131 );
buf ( n22133 , n6403 );
buf ( n22134 , n22133 );
and ( n22135 , n22132 , n22134 );
not ( n22136 , n22132 );
not ( n22137 , n22133 );
and ( n22138 , n22136 , n22137 );
nor ( n22139 , n22135 , n22138 );
xnor ( n22140 , n22130 , n22139 );
buf ( n22141 , n22140 );
not ( n22142 , n22141 );
or ( n22143 , n22104 , n22142 );
not ( n22144 , n11167 );
not ( n22145 , n22140 );
nand ( n22146 , n22144 , n22145 );
nand ( n22147 , n22143 , n22146 );
buf ( n22148 , n6404 );
buf ( n22149 , n22148 );
not ( n22150 , n22149 );
not ( n22151 , n13035 );
not ( n22152 , n22151 );
or ( n22153 , n22150 , n22152 );
not ( n22154 , n22148 );
nand ( n22155 , n22154 , n13036 );
nand ( n22156 , n22153 , n22155 );
buf ( n22157 , n6405 );
not ( n22158 , n22157 );
and ( n22159 , n22156 , n22158 );
not ( n22160 , n22156 );
buf ( n22161 , n22157 );
and ( n22162 , n22160 , n22161 );
nor ( n22163 , n22159 , n22162 );
buf ( n22164 , n6406 );
nand ( n22165 , n7477 , n22164 );
buf ( n22166 , n6407 );
not ( n22167 , n22166 );
and ( n22168 , n22165 , n22167 );
not ( n22169 , n22165 );
buf ( n22170 , n22166 );
and ( n22171 , n22169 , n22170 );
nor ( n22172 , n22168 , n22171 );
xor ( n22173 , n22163 , n22172 );
buf ( n22174 , n6408 );
nand ( n22175 , n7516 , n22174 );
buf ( n22176 , n6409 );
not ( n22177 , n22176 );
and ( n22178 , n22175 , n22177 );
not ( n22179 , n22175 );
buf ( n22180 , n22176 );
and ( n22181 , n22179 , n22180 );
nor ( n22182 , n22178 , n22181 );
xnor ( n22183 , n22173 , n22182 );
not ( n22184 , n22183 );
not ( n22185 , n22184 );
and ( n22186 , n22147 , n22185 );
not ( n22187 , n22147 );
not ( n22188 , n22183 );
buf ( n22189 , n22188 );
and ( n22190 , n22187 , n22189 );
nor ( n22191 , n22186 , n22190 );
not ( n22192 , n22191 );
and ( n22193 , n22103 , n22192 );
and ( n22194 , n22102 , n22191 );
nor ( n22195 , n22193 , n22194 );
not ( n22196 , n22195 );
not ( n22197 , n22196 );
buf ( n22198 , n6410 );
not ( n22199 , n13349 );
buf ( n22200 , n6411 );
not ( n22201 , n22200 );
not ( n22202 , n22201 );
or ( n22203 , n22199 , n22202 );
not ( n22204 , n13348 );
buf ( n22205 , n22200 );
nand ( n22206 , n22204 , n22205 );
nand ( n22207 , n22203 , n22206 );
xor ( n22208 , n22198 , n22207 );
buf ( n22209 , n6412 );
xor ( n22210 , n20709 , n22209 );
buf ( n22211 , n6413 );
nand ( n22212 , n7196 , n22211 );
xnor ( n22213 , n22210 , n22212 );
xnor ( n22214 , n22208 , n22213 );
buf ( n22215 , n22214 );
not ( n22216 , n22215 );
not ( n22217 , n13426 );
not ( n22218 , n11473 );
or ( n22219 , n22217 , n22218 );
nand ( n22220 , n11469 , n13422 );
nand ( n22221 , n22219 , n22220 );
not ( n22222 , n22221 );
or ( n22223 , n22216 , n22222 );
or ( n22224 , n22215 , n22221 );
nand ( n22225 , n22223 , n22224 );
not ( n22226 , n10695 );
not ( n22227 , n20430 );
or ( n22228 , n22226 , n22227 );
not ( n22229 , n10695 );
nand ( n22230 , n22229 , n20436 );
nand ( n22231 , n22228 , n22230 );
buf ( n22232 , n19449 );
not ( n22233 , n22232 );
and ( n22234 , n22231 , n22233 );
not ( n22235 , n22231 );
and ( n22236 , n22235 , n22232 );
nor ( n22237 , n22234 , n22236 );
not ( n22238 , n22237 );
nand ( n22239 , n22225 , n22238 );
buf ( n22240 , n19833 );
not ( n22241 , n22240 );
and ( n22242 , n22239 , n22241 );
not ( n22243 , n22239 );
and ( n22244 , n22243 , n22240 );
nor ( n22245 , n22242 , n22244 );
not ( n22246 , n22245 );
not ( n22247 , n22246 );
not ( n22248 , n18403 );
not ( n22249 , n9168 );
not ( n22250 , n17978 );
or ( n22251 , n22249 , n22250 );
not ( n22252 , n9168 );
nand ( n22253 , n22252 , n17979 );
nand ( n22254 , n22251 , n22253 );
not ( n22255 , n22254 );
and ( n22256 , n22248 , n22255 );
buf ( n22257 , n18403 );
and ( n22258 , n22257 , n22254 );
nor ( n22259 , n22256 , n22258 );
not ( n22260 , n8360 );
not ( n22261 , n14592 );
or ( n22262 , n22260 , n22261 );
not ( n22263 , n8360 );
nand ( n22264 , n22263 , n14596 );
nand ( n22265 , n22262 , n22264 );
and ( n22266 , n22265 , n14600 );
not ( n22267 , n22265 );
and ( n22268 , n22267 , n14603 );
nor ( n22269 , n22266 , n22268 );
nand ( n22270 , n22259 , n22269 );
not ( n22271 , n22270 );
not ( n22272 , n19651 );
and ( n22273 , n22271 , n22272 );
and ( n22274 , n22270 , n19651 );
nor ( n22275 , n22273 , n22274 );
not ( n22276 , n22275 );
not ( n22277 , n22276 );
or ( n22278 , n22247 , n22277 );
nand ( n22279 , n22275 , n22245 );
nand ( n22280 , n22278 , n22279 );
buf ( n22281 , n15886 );
buf ( n22282 , n10844 );
or ( n22283 , n22281 , n22282 );
nand ( n22284 , n10846 , n22281 );
nand ( n22285 , n22283 , n22284 );
not ( n22286 , n22285 );
not ( n22287 , n8145 );
not ( n22288 , n22287 );
buf ( n22289 , n22288 );
not ( n22290 , n22289 );
and ( n22291 , n22286 , n22290 );
and ( n22292 , n22285 , n22289 );
nor ( n22293 , n22291 , n22292 );
not ( n22294 , n14131 );
not ( n22295 , n18496 );
or ( n22296 , n22294 , n22295 );
not ( n22297 , n14131 );
nand ( n22298 , n22297 , n18491 );
nand ( n22299 , n22296 , n22298 );
not ( n22300 , n21471 );
not ( n22301 , n22300 );
and ( n22302 , n22299 , n22301 );
not ( n22303 , n22299 );
not ( n22304 , n21467 );
not ( n22305 , n22304 );
and ( n22306 , n22303 , n22305 );
nor ( n22307 , n22302 , n22306 );
nand ( n22308 , n22293 , n22307 );
not ( n22309 , n19740 );
and ( n22310 , n22308 , n22309 );
not ( n22311 , n22308 );
and ( n22312 , n22311 , n19740 );
nor ( n22313 , n22310 , n22312 );
not ( n22314 , n22313 );
and ( n22315 , n22280 , n22314 );
not ( n22316 , n22280 );
and ( n22317 , n22316 , n22313 );
nor ( n22318 , n22315 , n22317 );
not ( n22319 , n22191 );
not ( n22320 , n22101 );
nand ( n22321 , n22319 , n22320 );
not ( n22322 , n22321 );
not ( n22323 , n19678 );
and ( n22324 , n22322 , n22323 );
and ( n22325 , n22321 , n19678 );
nor ( n22326 , n22324 , n22325 );
not ( n22327 , n22326 );
not ( n22328 , n22327 );
not ( n22329 , n17126 );
buf ( n22330 , n8024 );
not ( n22331 , n22330 );
not ( n22332 , n17112 );
or ( n22333 , n22331 , n22332 );
not ( n22334 , n22330 );
nand ( n22335 , n22334 , n17309 );
nand ( n22336 , n22333 , n22335 );
not ( n22337 , n22336 );
and ( n22338 , n22329 , n22337 );
not ( n22339 , n17127 );
and ( n22340 , n22339 , n22336 );
nor ( n22341 , n22338 , n22340 );
not ( n22342 , n11924 );
not ( n22343 , n13289 );
not ( n22344 , n10278 );
or ( n22345 , n22343 , n22344 );
or ( n22346 , n10278 , n13289 );
nand ( n22347 , n22345 , n22346 );
not ( n22348 , n22347 );
and ( n22349 , n22342 , n22348 );
and ( n22350 , n16374 , n22347 );
nor ( n22351 , n22349 , n22350 );
not ( n22352 , n22351 );
nand ( n22353 , n22341 , n22352 );
not ( n22354 , n19934 );
and ( n22355 , n22353 , n22354 );
not ( n22356 , n22353 );
and ( n22357 , n22356 , n19934 );
nor ( n22358 , n22355 , n22357 );
not ( n22359 , n22358 );
not ( n22360 , n22359 );
or ( n22361 , n22328 , n22360 );
nand ( n22362 , n22358 , n22326 );
nand ( n22363 , n22361 , n22362 );
and ( n22364 , n22318 , n22363 );
not ( n22365 , n22318 );
not ( n22366 , n22363 );
and ( n22367 , n22365 , n22366 );
nor ( n22368 , n22364 , n22367 );
not ( n22369 , n22368 );
or ( n22370 , n22197 , n22369 );
not ( n22371 , n22196 );
not ( n22372 , n22366 );
not ( n22373 , n22318 );
not ( n22374 , n22373 );
or ( n22375 , n22372 , n22374 );
nand ( n22376 , n22318 , n22363 );
nand ( n22377 , n22375 , n22376 );
nand ( n22378 , n22371 , n22377 );
nand ( n22379 , n22370 , n22378 );
not ( n22380 , n21365 );
not ( n22381 , n8790 );
or ( n22382 , n22380 , n22381 );
buf ( n22383 , n8789 );
not ( n22384 , n22383 );
or ( n22385 , n22384 , n21365 );
nand ( n22386 , n22382 , n22385 );
not ( n22387 , n22386 );
not ( n22388 , n15273 );
and ( n22389 , n22387 , n22388 );
and ( n22390 , n22386 , n15254 );
nor ( n22391 , n22389 , n22390 );
not ( n22392 , n22391 );
not ( n22393 , n22392 );
not ( n22394 , n12174 );
not ( n22395 , n21201 );
or ( n22396 , n22394 , n22395 );
nand ( n22397 , n11058 , n12177 );
nand ( n22398 , n22396 , n22397 );
not ( n22399 , n22398 );
not ( n22400 , n19645 );
and ( n22401 , n22399 , n22400 );
and ( n22402 , n22398 , n19645 );
nor ( n22403 , n22401 , n22402 );
not ( n22404 , n22403 );
not ( n22405 , n10502 );
buf ( n22406 , n14054 );
not ( n22407 , n22406 );
or ( n22408 , n22405 , n22407 );
not ( n22409 , n10502 );
nand ( n22410 , n22409 , n14055 );
nand ( n22411 , n22408 , n22410 );
and ( n22412 , n22411 , n16363 );
not ( n22413 , n22411 );
and ( n22414 , n22413 , n16357 );
nor ( n22415 , n22412 , n22414 );
nand ( n22416 , n22404 , n22415 );
not ( n22417 , n22416 );
and ( n22418 , n22393 , n22417 );
and ( n22419 , n22392 , n22416 );
nor ( n22420 , n22418 , n22419 );
not ( n22421 , n22420 );
not ( n22422 , n22421 );
not ( n22423 , n8073 );
not ( n22424 , n9716 );
not ( n22425 , n8026 );
or ( n22426 , n22424 , n22425 );
or ( n22427 , n8026 , n9716 );
nand ( n22428 , n22426 , n22427 );
not ( n22429 , n22428 );
and ( n22430 , n22423 , n22429 );
and ( n22431 , n8074 , n22428 );
nor ( n22432 , n22430 , n22431 );
not ( n22433 , n22432 );
not ( n22434 , n22433 );
not ( n22435 , n20565 );
not ( n22436 , n10432 );
not ( n22437 , n11641 );
buf ( n22438 , n6414 );
not ( n22439 , n22438 );
not ( n22440 , n22439 );
or ( n22441 , n22437 , n22440 );
not ( n22442 , n11640 );
buf ( n22443 , n22438 );
nand ( n22444 , n22442 , n22443 );
nand ( n22445 , n22441 , n22444 );
buf ( n22446 , n6415 );
buf ( n22447 , n22446 );
and ( n22448 , n22445 , n22447 );
not ( n22449 , n22445 );
not ( n22450 , n22446 );
and ( n22451 , n22449 , n22450 );
nor ( n22452 , n22448 , n22451 );
not ( n22453 , n22452 );
buf ( n22454 , n6416 );
nand ( n22455 , n7921 , n22454 );
buf ( n22456 , n6417 );
buf ( n22457 , n22456 );
and ( n22458 , n22455 , n22457 );
not ( n22459 , n22455 );
not ( n22460 , n22456 );
and ( n22461 , n22459 , n22460 );
nor ( n22462 , n22458 , n22461 );
buf ( n22463 , n22462 );
xor ( n22464 , n22453 , n22463 );
buf ( n22465 , n6418 );
nand ( n22466 , n13379 , n22465 );
buf ( n22467 , n6419 );
not ( n22468 , n22467 );
and ( n22469 , n22466 , n22468 );
not ( n22470 , n22466 );
buf ( n22471 , n22467 );
and ( n22472 , n22470 , n22471 );
nor ( n22473 , n22469 , n22472 );
xnor ( n22474 , n22464 , n22473 );
not ( n22475 , n22474 );
or ( n22476 , n22436 , n22475 );
xor ( n22477 , n22452 , n22462 );
xnor ( n22478 , n22477 , n22473 );
nand ( n22479 , n22478 , n10428 );
nand ( n22480 , n22476 , n22479 );
not ( n22481 , n22480 );
and ( n22482 , n22435 , n22481 );
and ( n22483 , n20565 , n22480 );
nor ( n22484 , n22482 , n22483 );
not ( n22485 , n18192 );
not ( n22486 , n7315 );
not ( n22487 , n12748 );
or ( n22488 , n22486 , n22487 );
not ( n22489 , n7314 );
nand ( n22490 , n15458 , n22489 );
nand ( n22491 , n22488 , n22490 );
not ( n22492 , n22491 );
or ( n22493 , n22485 , n22492 );
or ( n22494 , n22491 , n18188 );
nand ( n22495 , n22493 , n22494 );
nand ( n22496 , n22484 , n22495 );
not ( n22497 , n22496 );
or ( n22498 , n22434 , n22497 );
or ( n22499 , n22496 , n22433 );
nand ( n22500 , n22498 , n22499 );
not ( n22501 , n22500 );
not ( n22502 , n22501 );
or ( n22503 , n22422 , n22502 );
nand ( n22504 , n22500 , n22420 );
nand ( n22505 , n22503 , n22504 );
not ( n22506 , n22505 );
buf ( n22507 , n6420 );
buf ( n22508 , n22507 );
not ( n22509 , n10273 );
xor ( n22510 , n22508 , n22509 );
xnor ( n22511 , n22510 , n10237 );
not ( n22512 , n22511 );
buf ( n22513 , n19254 );
not ( n22514 , n22513 );
not ( n22515 , n17918 );
or ( n22516 , n22514 , n22515 );
nand ( n22517 , n9075 , n19255 );
nand ( n22518 , n22516 , n22517 );
buf ( n22519 , n11104 );
and ( n22520 , n22518 , n22519 );
not ( n22521 , n22518 );
not ( n22522 , n11109 );
not ( n22523 , n22522 );
buf ( n22524 , n22523 );
and ( n22525 , n22521 , n22524 );
nor ( n22526 , n22520 , n22525 );
not ( n22527 , n22526 );
nand ( n22528 , n22512 , n22527 );
not ( n22529 , n22528 );
not ( n22530 , n12878 );
not ( n22531 , n16902 );
or ( n22532 , n22530 , n22531 );
or ( n22533 , n16902 , n12878 );
nand ( n22534 , n22532 , n22533 );
not ( n22535 , n8280 );
and ( n22536 , n22534 , n22535 );
not ( n22537 , n22534 );
and ( n22538 , n22537 , n8280 );
nor ( n22539 , n22536 , n22538 );
not ( n22540 , n22539 );
not ( n22541 , n22540 );
not ( n22542 , n22541 );
and ( n22543 , n22529 , n22542 );
and ( n22544 , n22528 , n22541 );
nor ( n22545 , n22543 , n22544 );
not ( n22546 , n22545 );
and ( n22547 , n22506 , n22546 );
and ( n22548 , n22505 , n22545 );
nor ( n22549 , n22547 , n22548 );
buf ( n22550 , n16625 );
and ( n22551 , n11609 , n22550 );
not ( n22552 , n11609 );
not ( n22553 , n22550 );
and ( n22554 , n22552 , n22553 );
nor ( n22555 , n22551 , n22554 );
not ( n22556 , n16585 );
not ( n22557 , n22556 );
not ( n22558 , n22557 );
and ( n22559 , n22555 , n22558 );
not ( n22560 , n22555 );
and ( n22561 , n22560 , n22557 );
nor ( n22562 , n22559 , n22561 );
not ( n22563 , n15519 );
not ( n22564 , n7310 );
not ( n22565 , n22564 );
or ( n22566 , n22563 , n22565 );
not ( n22567 , n22564 );
nand ( n22568 , n22567 , n15515 );
nand ( n22569 , n22566 , n22568 );
buf ( n22570 , n9531 );
not ( n22571 , n22570 );
buf ( n22572 , n22571 );
not ( n22573 , n22572 );
and ( n22574 , n22569 , n22573 );
not ( n22575 , n22569 );
and ( n22576 , n22575 , n22572 );
nor ( n22577 , n22574 , n22576 );
not ( n22578 , n22577 );
nand ( n22579 , n22562 , n22578 );
not ( n22580 , n7770 );
not ( n22581 , n15697 );
or ( n22582 , n22580 , n22581 );
not ( n22583 , n15748 );
nand ( n22584 , n22583 , n7766 );
nand ( n22585 , n22582 , n22584 );
buf ( n22586 , n6421 );
buf ( n22587 , n22586 );
not ( n22588 , n22587 );
buf ( n22589 , n6422 );
not ( n22590 , n22589 );
not ( n22591 , n22590 );
or ( n22592 , n22588 , n22591 );
not ( n22593 , n22586 );
buf ( n22594 , n22589 );
nand ( n22595 , n22593 , n22594 );
nand ( n22596 , n22592 , n22595 );
buf ( n22597 , n6423 );
not ( n22598 , n22597 );
and ( n22599 , n22596 , n22598 );
not ( n22600 , n22596 );
buf ( n22601 , n22597 );
and ( n22602 , n22600 , n22601 );
nor ( n22603 , n22599 , n22602 );
buf ( n22604 , n6424 );
nand ( n22605 , n7401 , n22604 );
buf ( n22606 , n6425 );
buf ( n22607 , n22606 );
and ( n22608 , n22605 , n22607 );
not ( n22609 , n22605 );
not ( n22610 , n22606 );
and ( n22611 , n22609 , n22610 );
nor ( n22612 , n22608 , n22611 );
xor ( n22613 , n22603 , n22612 );
xnor ( n22614 , n22613 , n20996 );
buf ( n22615 , n22614 );
and ( n22616 , n22585 , n22615 );
not ( n22617 , n22585 );
xor ( n22618 , n22603 , n20995 );
xnor ( n22619 , n22618 , n22612 );
buf ( n22620 , n22619 );
and ( n22621 , n22617 , n22620 );
nor ( n22622 , n22616 , n22621 );
xnor ( n22623 , n22579 , n22622 );
not ( n22624 , n22623 );
not ( n22625 , n18497 );
buf ( n22626 , n12002 );
not ( n22627 , n22626 );
not ( n22628 , n18456 );
not ( n22629 , n13253 );
or ( n22630 , n22628 , n22629 );
or ( n22631 , n18456 , n13253 );
nand ( n22632 , n22630 , n22631 );
xor ( n22633 , n22632 , n18447 );
buf ( n22634 , n22633 );
not ( n22635 , n22634 );
or ( n22636 , n22627 , n22635 );
or ( n22637 , n22634 , n22626 );
nand ( n22638 , n22636 , n22637 );
not ( n22639 , n22638 );
or ( n22640 , n22625 , n22639 );
or ( n22641 , n22638 , n18497 );
nand ( n22642 , n22640 , n22641 );
not ( n22643 , n22642 );
xor ( n22644 , n6982 , n21215 );
xnor ( n22645 , n22644 , n9489 );
not ( n22646 , n22645 );
nand ( n22647 , n22643 , n22646 );
not ( n22648 , n22647 );
xor ( n22649 , n15646 , n15614 );
buf ( n22650 , n15624 );
xnor ( n22651 , n22649 , n22650 );
nand ( n22652 , n22651 , n13352 );
not ( n22653 , n22652 );
nor ( n22654 , n22651 , n13352 );
nor ( n22655 , n22653 , n22654 );
not ( n22656 , n22655 );
not ( n22657 , n15604 );
or ( n22658 , n22656 , n22657 );
or ( n22659 , n15604 , n22655 );
nand ( n22660 , n22658 , n22659 );
not ( n22661 , n22660 );
not ( n22662 , n22661 );
not ( n22663 , n22662 );
and ( n22664 , n22648 , n22663 );
not ( n22665 , n22642 );
nand ( n22666 , n22665 , n22646 );
and ( n22667 , n22666 , n22662 );
nor ( n22668 , n22664 , n22667 );
not ( n22669 , n22668 );
not ( n22670 , n22669 );
or ( n22671 , n22624 , n22670 );
not ( n22672 , n22623 );
nand ( n22673 , n22672 , n22668 );
nand ( n22674 , n22671 , n22673 );
and ( n22675 , n22549 , n22674 );
not ( n22676 , n22549 );
not ( n22677 , n22674 );
and ( n22678 , n22676 , n22677 );
nor ( n22679 , n22675 , n22678 );
buf ( n22680 , n22679 );
and ( n22681 , n22379 , n22680 );
not ( n22682 , n22379 );
and ( n22683 , n22549 , n22677 );
not ( n22684 , n22549 );
and ( n22685 , n22684 , n22674 );
nor ( n22686 , n22683 , n22685 );
buf ( n22687 , n22686 );
and ( n22688 , n22682 , n22687 );
nor ( n22689 , n22681 , n22688 );
not ( n22690 , n22689 );
not ( n22691 , n22690 );
not ( n22692 , n19498 );
xor ( n22693 , n16471 , n12271 );
xnor ( n22694 , n22693 , n17732 );
not ( n22695 , n22694 );
nand ( n22696 , n22692 , n22695 );
not ( n22697 , n22696 );
not ( n22698 , n19417 );
and ( n22699 , n22697 , n22698 );
and ( n22700 , n22696 , n19417 );
nor ( n22701 , n22699 , n22700 );
not ( n22702 , n22701 );
not ( n22703 , n22702 );
not ( n22704 , n19576 );
or ( n22705 , n22703 , n22704 );
not ( n22706 , n22702 );
nand ( n22707 , n22706 , n19584 );
nand ( n22708 , n22705 , n22707 );
and ( n22709 , n22708 , n19990 );
not ( n22710 , n22708 );
and ( n22711 , n22710 , n19997 );
nor ( n22712 , n22709 , n22711 );
nand ( n22713 , n22691 , n22712 );
not ( n22714 , n22713 );
buf ( n22715 , n16838 );
not ( n22716 , n22715 );
not ( n22717 , n7899 );
not ( n22718 , n21955 );
or ( n22719 , n22717 , n22718 );
not ( n22720 , n7895 );
or ( n22721 , n21955 , n22720 );
nand ( n22722 , n22719 , n22721 );
and ( n22723 , n22722 , n21966 );
not ( n22724 , n22722 );
buf ( n22725 , n21918 );
not ( n22726 , n22725 );
and ( n22727 , n22724 , n22726 );
nor ( n22728 , n22723 , n22727 );
not ( n22729 , n22728 );
buf ( n22730 , n6426 );
nand ( n22731 , n7195 , n22730 );
buf ( n22732 , n6427 );
buf ( n22733 , n22732 );
and ( n22734 , n22731 , n22733 );
not ( n22735 , n22731 );
not ( n22736 , n22732 );
and ( n22737 , n22735 , n22736 );
nor ( n22738 , n22734 , n22737 );
not ( n22739 , n22738 );
not ( n22740 , n17481 );
or ( n22741 , n22739 , n22740 );
or ( n22742 , n17481 , n22738 );
nand ( n22743 , n22741 , n22742 );
buf ( n22744 , n6428 );
buf ( n22745 , n22744 );
not ( n22746 , n22745 );
buf ( n22747 , n6429 );
not ( n22748 , n22747 );
not ( n22749 , n22748 );
or ( n22750 , n22746 , n22749 );
not ( n22751 , n22744 );
buf ( n22752 , n22747 );
nand ( n22753 , n22751 , n22752 );
nand ( n22754 , n22750 , n22753 );
buf ( n22755 , n6430 );
buf ( n22756 , n22755 );
and ( n22757 , n22754 , n22756 );
not ( n22758 , n22754 );
not ( n22759 , n22755 );
and ( n22760 , n22758 , n22759 );
nor ( n22761 , n22757 , n22760 );
buf ( n22762 , n6431 );
nand ( n22763 , n8923 , n22762 );
buf ( n22764 , n6432 );
buf ( n22765 , n22764 );
and ( n22766 , n22763 , n22765 );
not ( n22767 , n22763 );
not ( n22768 , n22764 );
and ( n22769 , n22767 , n22768 );
nor ( n22770 , n22766 , n22769 );
xor ( n22771 , n22761 , n22770 );
buf ( n22772 , n6433 );
nand ( n22773 , n6761 , n22772 );
buf ( n22774 , n6434 );
buf ( n22775 , n22774 );
and ( n22776 , n22773 , n22775 );
not ( n22777 , n22773 );
not ( n22778 , n22774 );
and ( n22779 , n22777 , n22778 );
nor ( n22780 , n22776 , n22779 );
xnor ( n22781 , n22771 , n22780 );
not ( n22782 , n22781 );
not ( n22783 , n22782 );
buf ( n22784 , n22783 );
xor ( n22785 , n22743 , n22784 );
nand ( n22786 , n22729 , n22785 );
not ( n22787 , n22786 );
buf ( n22788 , n8830 );
not ( n22789 , n22788 );
not ( n22790 , n11173 );
not ( n22791 , n22790 );
or ( n22792 , n22789 , n22791 );
not ( n22793 , n22788 );
nand ( n22794 , n22793 , n11173 );
nand ( n22795 , n22792 , n22794 );
and ( n22796 , n22795 , n11185 );
not ( n22797 , n22795 );
and ( n22798 , n22797 , n21049 );
nor ( n22799 , n22796 , n22798 );
not ( n22800 , n22799 );
or ( n22801 , n22787 , n22800 );
or ( n22802 , n22799 , n22786 );
nand ( n22803 , n22801 , n22802 );
not ( n22804 , n22803 );
not ( n22805 , n22804 );
not ( n22806 , n14663 );
buf ( n22807 , n6435 );
nand ( n22808 , n6608 , n22807 );
buf ( n22809 , n6436 );
not ( n22810 , n22809 );
and ( n22811 , n22808 , n22810 );
not ( n22812 , n22808 );
buf ( n22813 , n22809 );
and ( n22814 , n22812 , n22813 );
nor ( n22815 , n22811 , n22814 );
not ( n22816 , n22815 );
buf ( n22817 , n6437 );
buf ( n22818 , n22817 );
not ( n22819 , n22818 );
buf ( n22820 , n6438 );
not ( n22821 , n22820 );
not ( n22822 , n22821 );
or ( n22823 , n22819 , n22822 );
not ( n22824 , n22817 );
buf ( n22825 , n22820 );
nand ( n22826 , n22824 , n22825 );
nand ( n22827 , n22823 , n22826 );
buf ( n22828 , n6439 );
buf ( n22829 , n22828 );
and ( n22830 , n22827 , n22829 );
not ( n22831 , n22827 );
not ( n22832 , n22828 );
and ( n22833 , n22831 , n22832 );
nor ( n22834 , n22830 , n22833 );
xor ( n22835 , n22834 , n9811 );
buf ( n22836 , n6440 );
nand ( n22837 , n7413 , n22836 );
buf ( n22838 , n6441 );
not ( n22839 , n22838 );
and ( n22840 , n22837 , n22839 );
not ( n22841 , n22837 );
buf ( n22842 , n22838 );
and ( n22843 , n22841 , n22842 );
nor ( n22844 , n22840 , n22843 );
xnor ( n22845 , n22835 , n22844 );
not ( n22846 , n22845 );
not ( n22847 , n22846 );
or ( n22848 , n22816 , n22847 );
not ( n22849 , n22815 );
nand ( n22850 , n22849 , n22845 );
nand ( n22851 , n22848 , n22850 );
not ( n22852 , n22851 );
and ( n22853 , n22806 , n22852 );
and ( n22854 , n14663 , n22851 );
nor ( n22855 , n22853 , n22854 );
not ( n22856 , n14534 );
not ( n22857 , n12895 );
not ( n22858 , n16901 );
or ( n22859 , n22857 , n22858 );
not ( n22860 , n12895 );
not ( n22861 , n16901 );
nand ( n22862 , n22860 , n22861 );
nand ( n22863 , n22859 , n22862 );
not ( n22864 , n22863 );
or ( n22865 , n22856 , n22864 );
or ( n22866 , n22863 , n8280 );
nand ( n22867 , n22865 , n22866 );
nand ( n22868 , n22855 , n22867 );
not ( n22869 , n22868 );
not ( n22870 , n21073 );
not ( n22871 , n6828 );
or ( n22872 , n22870 , n22871 );
or ( n22873 , n6828 , n21073 );
nand ( n22874 , n22872 , n22873 );
and ( n22875 , n22874 , n6874 );
not ( n22876 , n22874 );
not ( n22877 , n11281 );
and ( n22878 , n22876 , n22877 );
nor ( n22879 , n22875 , n22878 );
not ( n22880 , n22879 );
not ( n22881 , n22880 );
and ( n22882 , n22869 , n22881 );
and ( n22883 , n22868 , n22880 );
nor ( n22884 , n22882 , n22883 );
buf ( n22885 , n16521 );
not ( n22886 , n22885 );
not ( n22887 , n12270 );
or ( n22888 , n22886 , n22887 );
not ( n22889 , n22885 );
nand ( n22890 , n22889 , n12276 );
nand ( n22891 , n22888 , n22890 );
not ( n22892 , n22891 );
not ( n22893 , n19343 );
and ( n22894 , n22892 , n22893 );
buf ( n22895 , n19346 );
and ( n22896 , n22891 , n22895 );
nor ( n22897 , n22894 , n22896 );
buf ( n22898 , n21433 );
not ( n22899 , n22898 );
buf ( n22900 , n14205 );
not ( n22901 , n22900 );
not ( n22902 , n21467 );
or ( n22903 , n22901 , n22902 );
not ( n22904 , n22900 );
nand ( n22905 , n22904 , n21471 );
nand ( n22906 , n22903 , n22905 );
not ( n22907 , n22906 );
not ( n22908 , n22907 );
or ( n22909 , n22899 , n22908 );
not ( n22910 , n22898 );
nand ( n22911 , n22910 , n22906 );
nand ( n22912 , n22909 , n22911 );
nand ( n22913 , n22897 , n22912 );
not ( n22914 , n22913 );
not ( n22915 , n11658 );
not ( n22916 , n10331 );
or ( n22917 , n22915 , n22916 );
xor ( n22918 , n10310 , n10319 );
xor ( n22919 , n22918 , n10329 );
not ( n22920 , n22919 );
or ( n22921 , n22920 , n11658 );
nand ( n22922 , n22917 , n22921 );
and ( n22923 , n22922 , n14493 );
not ( n22924 , n22922 );
and ( n22925 , n22924 , n10376 );
nor ( n22926 , n22923 , n22925 );
not ( n22927 , n22926 );
and ( n22928 , n22914 , n22927 );
and ( n22929 , n22913 , n22926 );
nor ( n22930 , n22928 , n22929 );
xor ( n22931 , n22884 , n22930 );
not ( n22932 , n22799 );
not ( n22933 , n22785 );
nand ( n22934 , n22932 , n22933 );
not ( n22935 , n9605 );
not ( n22936 , n13708 );
or ( n22937 , n22935 , n22936 );
not ( n22938 , n9605 );
nand ( n22939 , n22938 , n15568 );
nand ( n22940 , n22937 , n22939 );
buf ( n22941 , n6442 );
buf ( n22942 , n22941 );
not ( n22943 , n22942 );
buf ( n22944 , n6443 );
not ( n22945 , n22944 );
not ( n22946 , n22945 );
or ( n22947 , n22943 , n22946 );
not ( n22948 , n22941 );
buf ( n22949 , n22944 );
nand ( n22950 , n22948 , n22949 );
nand ( n22951 , n22947 , n22950 );
not ( n22952 , n12518 );
and ( n22953 , n22951 , n22952 );
not ( n22954 , n22951 );
and ( n22955 , n22954 , n12519 );
nor ( n22956 , n22953 , n22955 );
xor ( n22957 , n22956 , n19549 );
xor ( n22958 , n22957 , n16207 );
not ( n22959 , n22958 );
buf ( n22960 , n22959 );
and ( n22961 , n22940 , n22960 );
not ( n22962 , n22940 );
buf ( n22963 , n22959 );
not ( n22964 , n22963 );
and ( n22965 , n22962 , n22964 );
nor ( n22966 , n22961 , n22965 );
and ( n22967 , n22934 , n22966 );
not ( n22968 , n22934 );
not ( n22969 , n22966 );
and ( n22970 , n22968 , n22969 );
nor ( n22971 , n22967 , n22970 );
xnor ( n22972 , n22931 , n22971 );
buf ( n22973 , n10416 );
not ( n22974 , n22973 );
not ( n22975 , n22188 );
not ( n22976 , n22975 );
or ( n22977 , n22974 , n22976 );
or ( n22978 , n22185 , n22973 );
nand ( n22979 , n22977 , n22978 );
buf ( n22980 , n22478 );
buf ( n22981 , n22980 );
and ( n22982 , n22979 , n22981 );
not ( n22983 , n22979 );
buf ( n22984 , n22474 );
buf ( n22985 , n22984 );
and ( n22986 , n22983 , n22985 );
nor ( n22987 , n22982 , n22986 );
not ( n22988 , n22987 );
not ( n22989 , n22650 );
not ( n22990 , n18724 );
or ( n22991 , n22989 , n22990 );
not ( n22992 , n22650 );
nand ( n22993 , n22992 , n18730 );
nand ( n22994 , n22991 , n22993 );
buf ( n22995 , n21296 );
and ( n22996 , n22994 , n22995 );
not ( n22997 , n22994 );
buf ( n22998 , n21297 );
and ( n22999 , n22997 , n22998 );
nor ( n23000 , n22996 , n22999 );
not ( n23001 , n23000 );
nand ( n23002 , n22988 , n23001 );
not ( n23003 , n23002 );
not ( n23004 , n12613 );
buf ( n23005 , n16142 );
not ( n23006 , n23005 );
or ( n23007 , n23004 , n23006 );
or ( n23008 , n23005 , n12613 );
nand ( n23009 , n23007 , n23008 );
not ( n23010 , n16183 );
and ( n23011 , n23009 , n23010 );
not ( n23012 , n23009 );
and ( n23013 , n23012 , n16183 );
nor ( n23014 , n23011 , n23013 );
not ( n23015 , n23014 );
not ( n23016 , n23015 );
and ( n23017 , n23003 , n23016 );
and ( n23018 , n23002 , n23015 );
nor ( n23019 , n23017 , n23018 );
not ( n23020 , n23019 );
buf ( n23021 , n16091 );
xor ( n23022 , n23021 , n17192 );
xnor ( n23023 , n23022 , n22257 );
not ( n23024 , n23023 );
and ( n23025 , n20937 , n20934 );
not ( n23026 , n20937 );
buf ( n23027 , n20933 );
and ( n23028 , n23026 , n23027 );
nor ( n23029 , n23025 , n23028 );
not ( n23030 , n23029 );
not ( n23031 , n9397 );
not ( n23032 , n23031 );
or ( n23033 , n23030 , n23032 );
not ( n23034 , n23029 );
nand ( n23035 , n23034 , n14489 );
nand ( n23036 , n23033 , n23035 );
and ( n23037 , n23036 , n9405 );
not ( n23038 , n23036 );
and ( n23039 , n23038 , n7672 );
nor ( n23040 , n23037 , n23039 );
not ( n23041 , n23040 );
nand ( n23042 , n23024 , n23041 );
not ( n23043 , n20031 );
not ( n23044 , n22615 );
or ( n23045 , n23043 , n23044 );
or ( n23046 , n22615 , n20031 );
nand ( n23047 , n23045 , n23046 );
not ( n23048 , n16782 );
and ( n23049 , n23047 , n23048 );
not ( n23050 , n23047 );
and ( n23051 , n23050 , n16782 );
nor ( n23052 , n23049 , n23051 );
and ( n23053 , n23042 , n23052 );
not ( n23054 , n23042 );
not ( n23055 , n23052 );
and ( n23056 , n23054 , n23055 );
nor ( n23057 , n23053 , n23056 );
not ( n23058 , n23057 );
or ( n23059 , n23020 , n23058 );
or ( n23060 , n23057 , n23019 );
nand ( n23061 , n23059 , n23060 );
xor ( n23062 , n22972 , n23061 );
not ( n23063 , n23062 );
not ( n23064 , n23063 );
or ( n23065 , n22805 , n23064 );
or ( n23066 , n23063 , n22804 );
nand ( n23067 , n23065 , n23066 );
not ( n23068 , n19917 );
buf ( n23069 , n19063 );
not ( n23070 , n23069 );
or ( n23071 , n23068 , n23070 );
not ( n23072 , n19917 );
nand ( n23073 , n23072 , n19064 );
nand ( n23074 , n23071 , n23073 );
and ( n23075 , n23074 , n19829 );
not ( n23076 , n23074 );
and ( n23077 , n23076 , n19110 );
nor ( n23078 , n23075 , n23077 );
not ( n23079 , n23078 );
not ( n23080 , n15760 );
buf ( n23081 , n8198 );
xor ( n23082 , n23081 , n8210 );
xnor ( n23083 , n23082 , n8236 );
not ( n23084 , n23083 );
or ( n23085 , n23080 , n23084 );
or ( n23086 , n23083 , n15760 );
nand ( n23087 , n23085 , n23086 );
buf ( n23088 , n17556 );
xor ( n23089 , n23088 , n17568 );
xnor ( n23090 , n23089 , n17575 );
not ( n23091 , n23090 );
and ( n23092 , n23087 , n23091 );
not ( n23093 , n23087 );
and ( n23094 , n23093 , n23090 );
nor ( n23095 , n23092 , n23094 );
not ( n23096 , n11513 );
buf ( n23097 , n6444 );
buf ( n23098 , n23097 );
not ( n23099 , n23098 );
buf ( n23100 , n6445 );
not ( n23101 , n23100 );
not ( n23102 , n23101 );
or ( n23103 , n23099 , n23102 );
not ( n23104 , n23097 );
buf ( n23105 , n23100 );
nand ( n23106 , n23104 , n23105 );
nand ( n23107 , n23103 , n23106 );
not ( n23108 , n23107 );
not ( n23109 , n23108 );
or ( n23110 , n23096 , n23109 );
nand ( n23111 , n23107 , n11509 );
nand ( n23112 , n23110 , n23111 );
not ( n23113 , n23112 );
buf ( n23114 , n6446 );
buf ( n23115 , n23114 );
xor ( n23116 , n23115 , n22738 );
buf ( n23117 , n6447 );
nand ( n23118 , n7413 , n23117 );
buf ( n23119 , n6448 );
not ( n23120 , n23119 );
and ( n23121 , n23118 , n23120 );
not ( n23122 , n23118 );
buf ( n23123 , n23119 );
and ( n23124 , n23122 , n23123 );
nor ( n23125 , n23121 , n23124 );
xnor ( n23126 , n23116 , n23125 );
not ( n23127 , n23126 );
not ( n23128 , n23127 );
or ( n23129 , n23113 , n23128 );
or ( n23130 , n23127 , n23112 );
nand ( n23131 , n23129 , n23130 );
buf ( n23132 , n6449 );
nand ( n23133 , n8923 , n23132 );
buf ( n23134 , n6450 );
buf ( n23135 , n23134 );
and ( n23136 , n23133 , n23135 );
not ( n23137 , n23133 );
not ( n23138 , n23134 );
and ( n23139 , n23137 , n23138 );
nor ( n23140 , n23136 , n23139 );
not ( n23141 , n23140 );
buf ( n23142 , n6451 );
nand ( n23143 , n7921 , n23142 );
buf ( n23144 , n6452 );
not ( n23145 , n23144 );
and ( n23146 , n23143 , n23145 );
not ( n23147 , n23143 );
buf ( n23148 , n23144 );
and ( n23149 , n23147 , n23148 );
nor ( n23150 , n23146 , n23149 );
not ( n23151 , n23150 );
or ( n23152 , n23141 , n23151 );
or ( n23153 , n23140 , n23150 );
nand ( n23154 , n23152 , n23153 );
buf ( n23155 , n6453 );
buf ( n23156 , n23155 );
not ( n23157 , n23156 );
buf ( n23158 , n6454 );
not ( n23159 , n23158 );
not ( n23160 , n23159 );
or ( n23161 , n23157 , n23160 );
not ( n23162 , n23155 );
buf ( n23163 , n23158 );
nand ( n23164 , n23162 , n23163 );
nand ( n23165 , n23161 , n23164 );
buf ( n23166 , n6455 );
not ( n23167 , n23166 );
and ( n23168 , n23165 , n23167 );
not ( n23169 , n23165 );
buf ( n23170 , n23166 );
and ( n23171 , n23169 , n23170 );
nor ( n23172 , n23168 , n23171 );
not ( n23173 , n23172 );
and ( n23174 , n23154 , n23173 );
not ( n23175 , n23154 );
and ( n23176 , n23175 , n23172 );
nor ( n23177 , n23174 , n23176 );
buf ( n23178 , n23177 );
and ( n23179 , n23131 , n23178 );
not ( n23180 , n23131 );
xor ( n23181 , n23172 , n23140 );
xnor ( n23182 , n23181 , n23150 );
buf ( n23183 , n23182 );
and ( n23184 , n23180 , n23183 );
nor ( n23185 , n23179 , n23184 );
not ( n23186 , n23185 );
nand ( n23187 , n23095 , n23186 );
not ( n23188 , n23187 );
or ( n23189 , n23079 , n23188 );
not ( n23190 , n23185 );
nand ( n23191 , n23190 , n23095 );
or ( n23192 , n23191 , n23078 );
nand ( n23193 , n23189 , n23192 );
not ( n23194 , n23193 );
not ( n23195 , n11395 );
not ( n23196 , n14520 );
not ( n23197 , n23196 );
or ( n23198 , n23195 , n23197 );
or ( n23199 , n23196 , n11395 );
nand ( n23200 , n23198 , n23199 );
xor ( n23201 , n18136 , n18132 );
and ( n23202 , n23200 , n23201 );
not ( n23203 , n23200 );
and ( n23204 , n23203 , n18138 );
nor ( n23205 , n23202 , n23204 );
not ( n23206 , n20204 );
xor ( n23207 , n19605 , n19624 );
not ( n23208 , n19614 );
xnor ( n23209 , n23207 , n23208 );
not ( n23210 , n23209 );
or ( n23211 , n23206 , n23210 );
or ( n23212 , n23209 , n20204 );
nand ( n23213 , n23211 , n23212 );
and ( n23214 , n23213 , n19634 );
not ( n23215 , n23213 );
and ( n23216 , n23215 , n19631 );
nor ( n23217 , n23214 , n23216 );
not ( n23218 , n23217 );
nand ( n23219 , n23205 , n23218 );
not ( n23220 , n23219 );
not ( n23221 , n9687 );
not ( n23222 , n6902 );
and ( n23223 , n23221 , n23222 );
not ( n23224 , n11378 );
and ( n23225 , n23224 , n6902 );
nor ( n23226 , n23223 , n23225 );
not ( n23227 , n22508 );
buf ( n23228 , n6456 );
not ( n23229 , n23228 );
not ( n23230 , n23229 );
or ( n23231 , n23227 , n23230 );
not ( n23232 , n22507 );
buf ( n23233 , n23228 );
nand ( n23234 , n23232 , n23233 );
nand ( n23235 , n23231 , n23234 );
buf ( n23236 , n6457 );
buf ( n23237 , n23236 );
and ( n23238 , n23235 , n23237 );
not ( n23239 , n23235 );
not ( n23240 , n23236 );
and ( n23241 , n23239 , n23240 );
nor ( n23242 , n23238 , n23241 );
xor ( n23243 , n23242 , n10213 );
xnor ( n23244 , n23243 , n21118 );
buf ( n23245 , n23244 );
buf ( n23246 , n23245 );
xor ( n23247 , n23226 , n23246 );
buf ( n23248 , n23247 );
not ( n23249 , n23248 );
and ( n23250 , n23220 , n23249 );
and ( n23251 , n23219 , n23248 );
nor ( n23252 , n23250 , n23251 );
not ( n23253 , n23252 );
or ( n23254 , n23194 , n23253 );
or ( n23255 , n23252 , n23193 );
nand ( n23256 , n23254 , n23255 );
buf ( n23257 , n21959 );
not ( n23258 , n23257 );
xor ( n23259 , n12968 , n23258 );
xnor ( n23260 , n23259 , n16446 );
not ( n23261 , n6647 );
not ( n23262 , n18982 );
or ( n23263 , n23261 , n23262 );
not ( n23264 , n6647 );
nand ( n23265 , n23264 , n18981 );
nand ( n23266 , n23263 , n23265 );
not ( n23267 , n12157 );
not ( n23268 , n23267 );
and ( n23269 , n23266 , n23268 );
not ( n23270 , n23266 );
xor ( n23271 , n12137 , n12156 );
xnor ( n23272 , n23271 , n12146 );
and ( n23273 , n23270 , n23272 );
nor ( n23274 , n23269 , n23273 );
not ( n23275 , n23274 );
nand ( n23276 , n23260 , n23275 );
not ( n23277 , n23276 );
not ( n23278 , n20055 );
not ( n23279 , n22614 );
or ( n23280 , n23278 , n23279 );
not ( n23281 , n20055 );
nand ( n23282 , n23281 , n22619 );
nand ( n23283 , n23280 , n23282 );
not ( n23284 , n23283 );
not ( n23285 , n23048 );
and ( n23286 , n23284 , n23285 );
and ( n23287 , n23283 , n23048 );
nor ( n23288 , n23286 , n23287 );
not ( n23289 , n23288 );
not ( n23290 , n23289 );
and ( n23291 , n23277 , n23290 );
and ( n23292 , n23276 , n23289 );
nor ( n23293 , n23291 , n23292 );
and ( n23294 , n23256 , n23293 );
not ( n23295 , n23256 );
not ( n23296 , n23293 );
and ( n23297 , n23295 , n23296 );
nor ( n23298 , n23294 , n23297 );
not ( n23299 , n23298 );
buf ( n23300 , n20783 );
not ( n23301 , n23300 );
buf ( n23302 , n21687 );
not ( n23303 , n23302 );
not ( n23304 , n23303 );
or ( n23305 , n23301 , n23304 );
not ( n23306 , n23300 );
not ( n23307 , n21688 );
nand ( n23308 , n23306 , n23307 );
nand ( n23309 , n23305 , n23308 );
not ( n23310 , n18593 );
not ( n23311 , n23310 );
and ( n23312 , n23309 , n23311 );
not ( n23313 , n23309 );
not ( n23314 , n23311 );
and ( n23315 , n23313 , n23314 );
nor ( n23316 , n23312 , n23315 );
not ( n23317 , n23316 );
not ( n23318 , n11229 );
not ( n23319 , n7855 );
and ( n23320 , n23318 , n23319 );
and ( n23321 , n19691 , n7855 );
nor ( n23322 , n23320 , n23321 );
and ( n23323 , n23322 , n20941 );
not ( n23324 , n23322 );
and ( n23325 , n23324 , n20940 );
nor ( n23326 , n23323 , n23325 );
not ( n23327 , n23326 );
not ( n23328 , n16254 );
not ( n23329 , n13798 );
buf ( n23330 , n23329 );
not ( n23331 , n23330 );
or ( n23332 , n23328 , n23331 );
not ( n23333 , n13799 );
nand ( n23334 , n23333 , n16260 );
nand ( n23335 , n23332 , n23334 );
not ( n23336 , n18511 );
buf ( n23337 , n6458 );
not ( n23338 , n23337 );
not ( n23339 , n23338 );
or ( n23340 , n23336 , n23339 );
not ( n23341 , n18510 );
buf ( n23342 , n23337 );
nand ( n23343 , n23341 , n23342 );
nand ( n23344 , n23340 , n23343 );
buf ( n23345 , n6459 );
not ( n23346 , n23345 );
and ( n23347 , n23344 , n23346 );
not ( n23348 , n23344 );
buf ( n23349 , n23345 );
and ( n23350 , n23348 , n23349 );
nor ( n23351 , n23347 , n23350 );
buf ( n23352 , n6460 );
nand ( n23353 , n7401 , n23352 );
buf ( n23354 , n6461 );
buf ( n23355 , n23354 );
and ( n23356 , n23353 , n23355 );
not ( n23357 , n23353 );
not ( n23358 , n23354 );
and ( n23359 , n23357 , n23358 );
nor ( n23360 , n23356 , n23359 );
not ( n23361 , n23360 );
xor ( n23362 , n23351 , n23361 );
buf ( n23363 , n6462 );
nand ( n23364 , n10204 , n23363 );
buf ( n23365 , n6463 );
not ( n23366 , n23365 );
and ( n23367 , n23364 , n23366 );
not ( n23368 , n23364 );
buf ( n23369 , n23365 );
and ( n23370 , n23368 , n23369 );
nor ( n23371 , n23367 , n23370 );
xnor ( n23372 , n23362 , n23371 );
buf ( n23373 , n23372 );
and ( n23374 , n23335 , n23373 );
not ( n23375 , n23335 );
not ( n23376 , n23360 );
not ( n23377 , n23371 );
or ( n23378 , n23376 , n23377 );
or ( n23379 , n23360 , n23371 );
nand ( n23380 , n23378 , n23379 );
and ( n23381 , n23380 , n23351 );
not ( n23382 , n23380 );
not ( n23383 , n23351 );
and ( n23384 , n23382 , n23383 );
nor ( n23385 , n23381 , n23384 );
buf ( n23386 , n23385 );
buf ( n23387 , n23386 );
and ( n23388 , n23375 , n23387 );
nor ( n23389 , n23374 , n23388 );
nand ( n23390 , n23327 , n23389 );
not ( n23391 , n23390 );
or ( n23392 , n23317 , n23391 );
nand ( n23393 , n23327 , n23389 );
or ( n23394 , n23393 , n23316 );
nand ( n23395 , n23392 , n23394 );
not ( n23396 , n23395 );
buf ( n23397 , n6464 );
buf ( n23398 , n23397 );
buf ( n23399 , n12591 );
xor ( n23400 , n23398 , n23399 );
xor ( n23401 , n23400 , n12531 );
not ( n23402 , n18513 );
buf ( n23403 , n6465 );
buf ( n23404 , n23403 );
not ( n23405 , n23404 );
buf ( n23406 , n6466 );
not ( n23407 , n23406 );
not ( n23408 , n23407 );
or ( n23409 , n23405 , n23408 );
not ( n23410 , n23403 );
buf ( n23411 , n23406 );
nand ( n23412 , n23410 , n23411 );
nand ( n23413 , n23409 , n23412 );
buf ( n23414 , n6467 );
not ( n23415 , n23414 );
and ( n23416 , n23413 , n23415 );
not ( n23417 , n23413 );
buf ( n23418 , n23414 );
and ( n23419 , n23417 , n23418 );
nor ( n23420 , n23416 , n23419 );
buf ( n23421 , n6468 );
nand ( n23422 , n7442 , n23421 );
buf ( n23423 , n6469 );
buf ( n23424 , n23423 );
and ( n23425 , n23422 , n23424 );
not ( n23426 , n23422 );
not ( n23427 , n23423 );
and ( n23428 , n23426 , n23427 );
nor ( n23429 , n23425 , n23428 );
xor ( n23430 , n23420 , n23429 );
buf ( n23431 , n6470 );
nand ( n23432 , n7288 , n23431 );
buf ( n23433 , n6471 );
buf ( n23434 , n23433 );
and ( n23435 , n23432 , n23434 );
not ( n23436 , n23432 );
not ( n23437 , n23433 );
and ( n23438 , n23436 , n23437 );
nor ( n23439 , n23435 , n23438 );
not ( n23440 , n23439 );
xnor ( n23441 , n23430 , n23440 );
not ( n23442 , n23441 );
or ( n23443 , n23402 , n23442 );
buf ( n23444 , n23441 );
or ( n23445 , n23444 , n18513 );
nand ( n23446 , n23443 , n23445 );
buf ( n23447 , n6472 );
buf ( n23448 , n23447 );
not ( n23449 , n23448 );
not ( n23450 , n18303 );
or ( n23451 , n23449 , n23450 );
not ( n23452 , n23447 );
buf ( n23453 , n18302 );
nand ( n23454 , n23452 , n23453 );
nand ( n23455 , n23451 , n23454 );
buf ( n23456 , n6473 );
not ( n23457 , n23456 );
and ( n23458 , n23455 , n23457 );
not ( n23459 , n23455 );
buf ( n23460 , n23456 );
and ( n23461 , n23459 , n23460 );
nor ( n23462 , n23458 , n23461 );
buf ( n23463 , n6474 );
nand ( n23464 , n7865 , n23463 );
buf ( n23465 , n6475 );
buf ( n23466 , n23465 );
and ( n23467 , n23464 , n23466 );
not ( n23468 , n23464 );
not ( n23469 , n23465 );
and ( n23470 , n23468 , n23469 );
nor ( n23471 , n23467 , n23470 );
xor ( n23472 , n23462 , n23471 );
buf ( n23473 , n6476 );
nand ( n23474 , n7477 , n23473 );
buf ( n23475 , n6477 );
buf ( n23476 , n23475 );
and ( n23477 , n23474 , n23476 );
not ( n23478 , n23474 );
not ( n23479 , n23475 );
and ( n23480 , n23478 , n23479 );
nor ( n23481 , n23477 , n23480 );
xnor ( n23482 , n23472 , n23481 );
buf ( n23483 , n23482 );
and ( n23484 , n23446 , n23483 );
not ( n23485 , n23446 );
xor ( n23486 , n23462 , n23481 );
not ( n23487 , n23471 );
xnor ( n23488 , n23486 , n23487 );
not ( n23489 , n23488 );
not ( n23490 , n23489 );
and ( n23491 , n23485 , n23490 );
nor ( n23492 , n23484 , n23491 );
not ( n23493 , n23492 );
nand ( n23494 , n23401 , n23493 );
not ( n23495 , n23494 );
buf ( n23496 , n17026 );
xor ( n23497 , n23496 , n18018 );
xor ( n23498 , n23497 , n9244 );
not ( n23499 , n23498 );
and ( n23500 , n23495 , n23499 );
nand ( n23501 , n23401 , n23493 );
and ( n23502 , n23501 , n23498 );
nor ( n23503 , n23500 , n23502 );
not ( n23504 , n23503 );
or ( n23505 , n23396 , n23504 );
or ( n23506 , n23503 , n23395 );
nand ( n23507 , n23505 , n23506 );
not ( n23508 , n23507 );
and ( n23509 , n23299 , n23508 );
and ( n23510 , n23298 , n23507 );
nor ( n23511 , n23509 , n23510 );
not ( n23512 , n23511 );
not ( n23513 , n23512 );
not ( n23514 , n23513 );
and ( n23515 , n23067 , n23514 );
not ( n23516 , n23067 );
buf ( n23517 , n23511 );
and ( n23518 , n23516 , n23517 );
nor ( n23519 , n23515 , n23518 );
not ( n23520 , n23519 );
nor ( n23521 , n22716 , n23520 );
not ( n23522 , n23521 );
or ( n23523 , n22714 , n23522 );
not ( n23524 , n22712 );
nand ( n23525 , n22689 , n13746 );
nor ( n23526 , n23524 , n23525 );
and ( n23527 , n23526 , n23520 );
buf ( n23528 , n13766 );
and ( n23529 , n8828 , n23528 );
nor ( n23530 , n23527 , n23529 );
nand ( n23531 , n23523 , n23530 );
buf ( n23532 , n23531 );
buf ( n23533 , n23532 );
nand ( n23534 , n11273 , n17300 );
not ( n23535 , n23534 );
not ( n23536 , n11191 );
not ( n23537 , n23536 );
or ( n23538 , n23535 , n23537 );
or ( n23539 , n23536 , n23534 );
nand ( n23540 , n23538 , n23539 );
not ( n23541 , n23540 );
not ( n23542 , n23541 );
not ( n23543 , n11750 );
or ( n23544 , n23542 , n23543 );
not ( n23545 , n23541 );
nand ( n23546 , n23545 , n11739 );
nand ( n23547 , n23544 , n23546 );
xor ( n23548 , n13328 , n13337 );
xnor ( n23549 , n23548 , n13341 );
xor ( n23550 , n17108 , n23549 );
xnor ( n23551 , n23550 , n21576 );
not ( n23552 , n11473 );
buf ( n23553 , n13481 );
not ( n23554 , n23553 );
not ( n23555 , n21832 );
or ( n23556 , n23554 , n23555 );
or ( n23557 , n21832 , n23553 );
nand ( n23558 , n23556 , n23557 );
not ( n23559 , n23558 );
or ( n23560 , n23552 , n23559 );
buf ( n23561 , n11468 );
or ( n23562 , n23558 , n23561 );
nand ( n23563 , n23560 , n23562 );
nand ( n23564 , n23551 , n23563 );
not ( n23565 , n23564 );
not ( n23566 , n16567 );
not ( n23567 , n17208 );
or ( n23568 , n23566 , n23567 );
not ( n23569 , n16567 );
nand ( n23570 , n23569 , n7105 );
nand ( n23571 , n23568 , n23570 );
buf ( n23572 , n7144 );
and ( n23573 , n23571 , n23572 );
not ( n23574 , n23571 );
not ( n23575 , n23572 );
and ( n23576 , n23574 , n23575 );
nor ( n23577 , n23573 , n23576 );
not ( n23578 , n23577 );
not ( n23579 , n23578 );
and ( n23580 , n23565 , n23579 );
and ( n23581 , n23564 , n23578 );
nor ( n23582 , n23580 , n23581 );
not ( n23583 , n12076 );
not ( n23584 , n17774 );
and ( n23585 , n23583 , n23584 );
and ( n23586 , n12076 , n17774 );
nor ( n23587 , n23585 , n23586 );
and ( n23588 , n23587 , n12019 );
not ( n23589 , n23587 );
and ( n23590 , n23589 , n12089 );
nor ( n23591 , n23588 , n23590 );
not ( n23592 , n7953 );
not ( n23593 , n21918 );
or ( n23594 , n23592 , n23593 );
or ( n23595 , n21918 , n7953 );
nand ( n23596 , n23594 , n23595 );
and ( n23597 , n23596 , n23069 );
not ( n23598 , n23596 );
not ( n23599 , n23069 );
and ( n23600 , n23598 , n23599 );
nor ( n23601 , n23597 , n23600 );
nor ( n23602 , n23591 , n23601 );
not ( n23603 , n23602 );
not ( n23604 , n15793 );
not ( n23605 , n9320 );
not ( n23606 , n19026 );
or ( n23607 , n23605 , n23606 );
or ( n23608 , n19026 , n9320 );
nand ( n23609 , n23607 , n23608 );
not ( n23610 , n23609 );
and ( n23611 , n23604 , n23610 );
and ( n23612 , n15793 , n23609 );
nor ( n23613 , n23611 , n23612 );
not ( n23614 , n23613 );
or ( n23615 , n23603 , n23614 );
not ( n23616 , n23602 );
not ( n23617 , n23613 );
nand ( n23618 , n23616 , n23617 );
nand ( n23619 , n23615 , n23618 );
xor ( n23620 , n23582 , n23619 );
not ( n23621 , n10845 );
buf ( n23622 , n6478 );
nand ( n23623 , n8934 , n23622 );
buf ( n23624 , n6479 );
not ( n23625 , n23624 );
and ( n23626 , n23623 , n23625 );
not ( n23627 , n23623 );
buf ( n23628 , n23624 );
and ( n23629 , n23627 , n23628 );
nor ( n23630 , n23626 , n23629 );
buf ( n23631 , n23630 );
not ( n23632 , n23631 );
not ( n23633 , n14756 );
or ( n23634 , n23632 , n23633 );
not ( n23635 , n23631 );
nand ( n23636 , n23635 , n10809 );
nand ( n23637 , n23634 , n23636 );
not ( n23638 , n23637 );
and ( n23639 , n23621 , n23638 );
not ( n23640 , n10844 );
and ( n23641 , n23640 , n23637 );
nor ( n23642 , n23639 , n23641 );
not ( n23643 , n23642 );
buf ( n23644 , n8232 );
not ( n23645 , n23644 );
not ( n23646 , n6960 );
or ( n23647 , n23645 , n23646 );
not ( n23648 , n23644 );
nand ( n23649 , n23648 , n6956 );
nand ( n23650 , n23647 , n23649 );
and ( n23651 , n23650 , n19174 );
not ( n23652 , n23650 );
and ( n23653 , n23652 , n19187 );
nor ( n23654 , n23651 , n23653 );
nand ( n23655 , n23643 , n23654 );
not ( n23656 , n23655 );
not ( n23657 , n10516 );
not ( n23658 , n16309 );
or ( n23659 , n23657 , n23658 );
nand ( n23660 , n14056 , n10513 );
nand ( n23661 , n23659 , n23660 );
and ( n23662 , n23661 , n16357 );
not ( n23663 , n23661 );
and ( n23664 , n23663 , n16363 );
nor ( n23665 , n23662 , n23664 );
not ( n23666 , n23665 );
and ( n23667 , n23656 , n23666 );
and ( n23668 , n23655 , n23665 );
nor ( n23669 , n23667 , n23668 );
xor ( n23670 , n23620 , n23669 );
not ( n23671 , n21570 );
nor ( n23672 , n23671 , n11260 );
not ( n23673 , n23672 );
not ( n23674 , n21570 );
nand ( n23675 , n23674 , n11260 );
nand ( n23676 , n23673 , n23675 );
and ( n23677 , n23676 , n19690 );
not ( n23678 , n23676 );
and ( n23679 , n23678 , n19691 );
nor ( n23680 , n23677 , n23679 );
not ( n23681 , n23680 );
not ( n23682 , n20363 );
not ( n23683 , n14641 );
or ( n23684 , n23682 , n23683 );
not ( n23685 , n20363 );
nand ( n23686 , n23685 , n14642 );
nand ( n23687 , n23684 , n23686 );
and ( n23688 , n23687 , n10995 );
not ( n23689 , n23687 );
and ( n23690 , n23689 , n11009 );
nor ( n23691 , n23688 , n23690 );
not ( n23692 , n23691 );
nand ( n23693 , n23681 , n23692 );
buf ( n23694 , n21960 );
xor ( n23695 , n12979 , n23694 );
xor ( n23696 , n23695 , n16446 );
not ( n23697 , n23696 );
and ( n23698 , n23693 , n23697 );
not ( n23699 , n23693 );
and ( n23700 , n23699 , n23696 );
nor ( n23701 , n23698 , n23700 );
not ( n23702 , n23701 );
not ( n23703 , n23702 );
buf ( n23704 , n18186 );
not ( n23705 , n6828 );
xor ( n23706 , n23704 , n23705 );
buf ( n23707 , n8328 );
not ( n23708 , n23707 );
xnor ( n23709 , n23706 , n23708 );
xor ( n23710 , n19437 , n17495 );
not ( n23711 , n19447 );
xnor ( n23712 , n23710 , n23711 );
not ( n23713 , n23712 );
buf ( n23714 , n10728 );
nor ( n23715 , n23713 , n23714 );
not ( n23716 , n23715 );
nand ( n23717 , n23714 , n22233 );
nand ( n23718 , n23716 , n23717 );
and ( n23719 , n23718 , n19493 );
not ( n23720 , n23718 );
not ( n23721 , n19490 );
not ( n23722 , n23721 );
and ( n23723 , n23720 , n23722 );
nor ( n23724 , n23719 , n23723 );
not ( n23725 , n23724 );
nand ( n23726 , n23709 , n23725 );
buf ( n23727 , n6480 );
buf ( n23728 , n23727 );
not ( n23729 , n23728 );
not ( n23730 , n23398 );
buf ( n23731 , n6481 );
not ( n23732 , n23731 );
not ( n23733 , n23732 );
or ( n23734 , n23730 , n23733 );
not ( n23735 , n23397 );
buf ( n23736 , n23731 );
nand ( n23737 , n23735 , n23736 );
nand ( n23738 , n23734 , n23737 );
and ( n23739 , n23738 , n8627 );
not ( n23740 , n23738 );
not ( n23741 , n8626 );
and ( n23742 , n23740 , n23741 );
nor ( n23743 , n23739 , n23742 );
buf ( n23744 , n6482 );
nand ( n23745 , n7865 , n23744 );
buf ( n23746 , n6483 );
not ( n23747 , n23746 );
and ( n23748 , n23745 , n23747 );
not ( n23749 , n23745 );
buf ( n23750 , n23746 );
and ( n23751 , n23749 , n23750 );
nor ( n23752 , n23748 , n23751 );
xor ( n23753 , n23743 , n23752 );
buf ( n23754 , n6484 );
nand ( n23755 , n8785 , n23754 );
buf ( n23756 , n6485 );
not ( n23757 , n23756 );
and ( n23758 , n23755 , n23757 );
not ( n23759 , n23755 );
buf ( n23760 , n23756 );
and ( n23761 , n23759 , n23760 );
nor ( n23762 , n23758 , n23761 );
xnor ( n23763 , n23753 , n23762 );
not ( n23764 , n23763 );
not ( n23765 , n23764 );
not ( n23766 , n23765 );
or ( n23767 , n23729 , n23766 );
not ( n23768 , n23763 );
not ( n23769 , n23768 );
or ( n23770 , n23769 , n23728 );
nand ( n23771 , n23767 , n23770 );
buf ( n23772 , n6486 );
buf ( n23773 , n6487 );
buf ( n23774 , n23773 );
not ( n23775 , n23774 );
buf ( n23776 , n6488 );
not ( n23777 , n23776 );
not ( n23778 , n23777 );
or ( n23779 , n23775 , n23778 );
not ( n23780 , n23773 );
buf ( n23781 , n23776 );
nand ( n23782 , n23780 , n23781 );
nand ( n23783 , n23779 , n23782 );
xor ( n23784 , n23772 , n23783 );
buf ( n23785 , n6489 );
xor ( n23786 , n12589 , n23785 );
buf ( n23787 , n6490 );
nand ( n23788 , n6985 , n23787 );
xnor ( n23789 , n23786 , n23788 );
xnor ( n23790 , n23784 , n23789 );
not ( n23791 , n23790 );
not ( n23792 , n23791 );
and ( n23793 , n23771 , n23792 );
not ( n23794 , n23771 );
and ( n23795 , n23794 , n23791 );
nor ( n23796 , n23793 , n23795 );
and ( n23797 , n23726 , n23796 );
not ( n23798 , n23726 );
not ( n23799 , n23796 );
and ( n23800 , n23798 , n23799 );
nor ( n23801 , n23797 , n23800 );
not ( n23802 , n23801 );
not ( n23803 , n23802 );
or ( n23804 , n23703 , n23803 );
nand ( n23805 , n23801 , n23701 );
nand ( n23806 , n23804 , n23805 );
and ( n23807 , n23670 , n23806 );
not ( n23808 , n23670 );
not ( n23809 , n23806 );
and ( n23810 , n23808 , n23809 );
nor ( n23811 , n23807 , n23810 );
not ( n23812 , n23811 );
buf ( n23813 , n23812 );
and ( n23814 , n23547 , n23813 );
not ( n23815 , n23547 );
not ( n23816 , n23813 );
and ( n23817 , n23815 , n23816 );
nor ( n23818 , n23814 , n23817 );
not ( n23819 , n23818 );
not ( n23820 , n21004 );
not ( n23821 , n16801 );
or ( n23822 , n23820 , n23821 );
buf ( n23823 , n15053 );
nand ( n23824 , n23823 , n21000 );
nand ( n23825 , n23822 , n23824 );
not ( n23826 , n13946 );
and ( n23827 , n23825 , n23826 );
not ( n23828 , n23825 );
buf ( n23829 , n13946 );
and ( n23830 , n23828 , n23829 );
nor ( n23831 , n23827 , n23830 );
not ( n23832 , n23831 );
not ( n23833 , n7076 );
not ( n23834 , n21193 );
or ( n23835 , n23833 , n23834 );
nand ( n23836 , n21178 , n7079 );
nand ( n23837 , n23835 , n23836 );
and ( n23838 , n23837 , n13158 );
not ( n23839 , n23837 );
and ( n23840 , n23839 , n13165 );
nor ( n23841 , n23838 , n23840 );
not ( n23842 , n21061 );
not ( n23843 , n8293 );
or ( n23844 , n23842 , n23843 );
or ( n23845 , n8293 , n21061 );
nand ( n23846 , n23844 , n23845 );
not ( n23847 , n6877 );
and ( n23848 , n23846 , n23847 );
not ( n23849 , n23846 );
and ( n23850 , n23849 , n6877 );
nor ( n23851 , n23848 , n23850 );
nand ( n23852 , n23841 , n23851 );
not ( n23853 , n23852 );
or ( n23854 , n23832 , n23853 );
or ( n23855 , n23852 , n23831 );
nand ( n23856 , n23854 , n23855 );
not ( n23857 , n23856 );
not ( n23858 , n10527 );
not ( n23859 , n14055 );
or ( n23860 , n23858 , n23859 );
not ( n23861 , n10527 );
nand ( n23862 , n23861 , n22406 );
nand ( n23863 , n23860 , n23862 );
and ( n23864 , n23863 , n16363 );
not ( n23865 , n23863 );
and ( n23866 , n23865 , n16357 );
nor ( n23867 , n23864 , n23866 );
not ( n23868 , n23867 );
not ( n23869 , n23868 );
not ( n23870 , n23196 );
not ( n23871 , n11687 );
not ( n23872 , n10375 );
or ( n23873 , n23871 , n23872 );
nand ( n23874 , n10374 , n11683 );
nand ( n23875 , n23873 , n23874 );
not ( n23876 , n23875 );
and ( n23877 , n23870 , n23876 );
and ( n23878 , n14522 , n23875 );
nor ( n23879 , n23877 , n23878 );
not ( n23880 , n23879 );
not ( n23881 , n12555 );
not ( n23882 , n21571 );
or ( n23883 , n23881 , n23882 );
or ( n23884 , n21571 , n12555 );
nand ( n23885 , n23883 , n23884 );
not ( n23886 , n23885 );
not ( n23887 , n7886 );
or ( n23888 , n23886 , n23887 );
or ( n23889 , n7886 , n23885 );
nand ( n23890 , n23888 , n23889 );
not ( n23891 , n23890 );
nand ( n23892 , n23880 , n23891 );
not ( n23893 , n23892 );
or ( n23894 , n23869 , n23893 );
or ( n23895 , n23892 , n23868 );
nand ( n23896 , n23894 , n23895 );
not ( n23897 , n23896 );
buf ( n23898 , n6491 );
buf ( n23899 , n23898 );
not ( n23900 , n23899 );
not ( n23901 , n11129 );
or ( n23902 , n23900 , n23901 );
not ( n23903 , n23899 );
nand ( n23904 , n23903 , n20391 );
nand ( n23905 , n23902 , n23904 );
and ( n23906 , n23905 , n20437 );
not ( n23907 , n23905 );
and ( n23908 , n23907 , n20431 );
nor ( n23909 , n23906 , n23908 );
not ( n23910 , n23909 );
not ( n23911 , n22846 );
not ( n23912 , n23911 );
not ( n23913 , n23912 );
not ( n23914 , n11325 );
xor ( n23915 , n7823 , n7842 );
xnor ( n23916 , n23915 , n7832 );
not ( n23917 , n23916 );
or ( n23918 , n23914 , n23917 );
or ( n23919 , n23916 , n11325 );
nand ( n23920 , n23918 , n23919 );
not ( n23921 , n23920 );
or ( n23922 , n23913 , n23921 );
not ( n23923 , n23911 );
or ( n23924 , n23920 , n23923 );
nand ( n23925 , n23922 , n23924 );
nand ( n23926 , n23910 , n23925 );
not ( n23927 , n23926 );
not ( n23928 , n19959 );
not ( n23929 , n10462 );
or ( n23930 , n23928 , n23929 );
or ( n23931 , n10462 , n19959 );
nand ( n23932 , n23930 , n23931 );
and ( n23933 , n23932 , n21528 );
not ( n23934 , n23932 );
not ( n23935 , n21528 );
and ( n23936 , n23934 , n23935 );
nor ( n23937 , n23933 , n23936 );
not ( n23938 , n23937 );
not ( n23939 , n23938 );
and ( n23940 , n23927 , n23939 );
and ( n23941 , n23926 , n23938 );
nor ( n23942 , n23940 , n23941 );
not ( n23943 , n23942 );
or ( n23944 , n23897 , n23943 );
or ( n23945 , n23942 , n23896 );
nand ( n23946 , n23944 , n23945 );
xor ( n23947 , n9739 , n17582 );
buf ( n23948 , n23090 );
xnor ( n23949 , n23947 , n23948 );
not ( n23950 , n23949 );
not ( n23951 , n6895 );
not ( n23952 , n11379 );
not ( n23953 , n23952 );
or ( n23954 , n23951 , n23953 );
not ( n23955 , n23224 );
nand ( n23956 , n23955 , n6898 );
nand ( n23957 , n23954 , n23956 );
not ( n23958 , n23246 );
not ( n23959 , n23958 );
and ( n23960 , n23957 , n23959 );
not ( n23961 , n23957 );
not ( n23962 , n23246 );
and ( n23963 , n23961 , n23962 );
nor ( n23964 , n23960 , n23963 );
nand ( n23965 , n23950 , n23964 );
buf ( n23966 , n11618 );
nor ( n23967 , n22550 , n23966 );
not ( n23968 , n23967 );
nand ( n23969 , n23966 , n22550 );
nand ( n23970 , n23968 , n23969 );
xnor ( n23971 , n23970 , n22557 );
not ( n23972 , n23971 );
and ( n23973 , n23965 , n23972 );
not ( n23974 , n23965 );
and ( n23975 , n23974 , n23971 );
nor ( n23976 , n23973 , n23975 );
and ( n23977 , n23946 , n23976 );
not ( n23978 , n23946 );
not ( n23979 , n23976 );
and ( n23980 , n23978 , n23979 );
nor ( n23981 , n23977 , n23980 );
not ( n23982 , n23831 );
not ( n23983 , n23851 );
nand ( n23984 , n23982 , n23983 );
not ( n23985 , n23984 );
buf ( n23986 , n12624 );
not ( n23987 , n23986 );
buf ( n23988 , n16137 );
not ( n23989 , n23988 );
or ( n23990 , n23987 , n23989 );
or ( n23991 , n23988 , n23986 );
nand ( n23992 , n23990 , n23991 );
and ( n23993 , n23992 , n16184 );
not ( n23994 , n23992 );
and ( n23995 , n23994 , n16183 );
nor ( n23996 , n23993 , n23995 );
not ( n23997 , n23996 );
not ( n23998 , n23997 );
and ( n23999 , n23985 , n23998 );
and ( n24000 , n23984 , n23997 );
nor ( n24001 , n23999 , n24000 );
not ( n24002 , n24001 );
not ( n24003 , n20794 );
buf ( n24004 , n24003 );
and ( n24005 , n17637 , n24004 );
not ( n24006 , n17637 );
buf ( n24007 , n20795 );
not ( n24008 , n24007 );
and ( n24009 , n24006 , n24008 );
nor ( n24010 , n24005 , n24009 );
not ( n24011 , n24010 );
not ( n24012 , n24011 );
buf ( n24013 , n20809 );
not ( n24014 , n24013 );
not ( n24015 , n24014 );
or ( n24016 , n24012 , n24015 );
nand ( n24017 , n24013 , n24010 );
nand ( n24018 , n24016 , n24017 );
not ( n24019 , n24018 );
not ( n24020 , n7735 );
not ( n24021 , n15743 );
or ( n24022 , n24020 , n24021 );
or ( n24023 , n15743 , n7735 );
nand ( n24024 , n24022 , n24023 );
not ( n24025 , n24024 );
not ( n24026 , n21273 );
not ( n24027 , n24026 );
and ( n24028 , n24025 , n24027 );
and ( n24029 , n24024 , n15697 );
nor ( n24030 , n24028 , n24029 );
not ( n24031 , n24030 );
nand ( n24032 , n24019 , n24031 );
not ( n24033 , n12039 );
not ( n24034 , n24033 );
not ( n24035 , n15988 );
not ( n24036 , n24035 );
or ( n24037 , n24034 , n24036 );
not ( n24038 , n24035 );
nand ( n24039 , n24038 , n12039 );
nand ( n24040 , n24037 , n24039 );
and ( n24041 , n24040 , n22634 );
not ( n24042 , n24040 );
not ( n24043 , n22634 );
and ( n24044 , n24042 , n24043 );
nor ( n24045 , n24041 , n24044 );
buf ( n24046 , n24045 );
xor ( n24047 , n24032 , n24046 );
not ( n24048 , n24047 );
or ( n24049 , n24002 , n24048 );
or ( n24050 , n24047 , n24001 );
nand ( n24051 , n24049 , n24050 );
not ( n24052 , n24051 );
and ( n24053 , n23981 , n24052 );
not ( n24054 , n23981 );
and ( n24055 , n24054 , n24051 );
nor ( n24056 , n24053 , n24055 );
buf ( n24057 , n24056 );
not ( n24058 , n24057 );
or ( n24059 , n23857 , n24058 );
not ( n24060 , n23856 );
not ( n24061 , n24056 );
nand ( n24062 , n24060 , n24061 );
nand ( n24063 , n24059 , n24062 );
not ( n24064 , n24063 );
buf ( n24065 , n9063 );
not ( n24066 , n24065 );
not ( n24067 , n22088 );
or ( n24068 , n24066 , n24067 );
or ( n24069 , n22088 , n24065 );
nand ( n24070 , n24068 , n24069 );
not ( n24071 , n24070 );
not ( n24072 , n18780 );
or ( n24073 , n24071 , n24072 );
or ( n24074 , n18780 , n24070 );
nand ( n24075 , n24073 , n24074 );
not ( n24076 , n17730 );
not ( n24077 , n22570 );
or ( n24078 , n24076 , n24077 );
not ( n24079 , n17730 );
nand ( n24080 , n24079 , n9532 );
nand ( n24081 , n24078 , n24080 );
and ( n24082 , n24081 , n9538 );
not ( n24083 , n24081 );
not ( n24084 , n9543 );
not ( n24085 , n24084 );
and ( n24086 , n24083 , n24085 );
nor ( n24087 , n24082 , n24086 );
not ( n24088 , n24087 );
nand ( n24089 , n24075 , n24088 );
not ( n24090 , n24089 );
not ( n24091 , n12428 );
not ( n24092 , n19411 );
or ( n24093 , n24091 , n24092 );
not ( n24094 , n12428 );
nand ( n24095 , n24094 , n15369 );
nand ( n24096 , n24093 , n24095 );
and ( n24097 , n24096 , n15395 );
not ( n24098 , n24096 );
not ( n24099 , n15395 );
and ( n24100 , n24098 , n24099 );
nor ( n24101 , n24097 , n24100 );
not ( n24102 , n24101 );
not ( n24103 , n24102 );
not ( n24104 , n24103 );
and ( n24105 , n24090 , n24104 );
and ( n24106 , n24089 , n24103 );
nor ( n24107 , n24105 , n24106 );
not ( n24108 , n24107 );
not ( n24109 , n24108 );
xor ( n24110 , n11517 , n23178 );
not ( n24111 , n23126 );
not ( n24112 , n23108 );
and ( n24113 , n24111 , n24112 );
and ( n24114 , n23126 , n23108 );
nor ( n24115 , n24113 , n24114 );
not ( n24116 , n24115 );
xnor ( n24117 , n24110 , n24116 );
not ( n24118 , n12323 );
not ( n24119 , n24118 );
not ( n24120 , n8950 );
or ( n24121 , n24119 , n24120 );
nand ( n24122 , n8945 , n12323 );
nand ( n24123 , n24121 , n24122 );
not ( n24124 , n24123 );
not ( n24125 , n8977 );
and ( n24126 , n24124 , n24125 );
and ( n24127 , n8977 , n24123 );
nor ( n24128 , n24126 , n24127 );
not ( n24129 , n24128 );
nand ( n24130 , n24117 , n24129 );
not ( n24131 , n9816 );
not ( n24132 , n7671 );
or ( n24133 , n24131 , n24132 );
or ( n24134 , n7671 , n9816 );
nand ( n24135 , n24133 , n24134 );
and ( n24136 , n24135 , n7716 );
not ( n24137 , n24135 );
not ( n24138 , n21251 );
and ( n24139 , n24137 , n24138 );
nor ( n24140 , n24136 , n24139 );
and ( n24141 , n24130 , n24140 );
not ( n24142 , n24130 );
not ( n24143 , n24140 );
and ( n24144 , n24142 , n24143 );
nor ( n24145 , n24141 , n24144 );
not ( n24146 , n24145 );
not ( n24147 , n24146 );
or ( n24148 , n24109 , n24147 );
nand ( n24149 , n24145 , n24107 );
nand ( n24150 , n24148 , n24149 );
xor ( n24151 , n22780 , n9032 );
xnor ( n24152 , n24151 , n19924 );
buf ( n24153 , n15215 );
not ( n24154 , n24153 );
buf ( n24155 , n6492 );
buf ( n24156 , n24155 );
not ( n24157 , n24156 );
not ( n24158 , n23898 );
not ( n24159 , n24158 );
or ( n24160 , n24157 , n24159 );
not ( n24161 , n24155 );
nand ( n24162 , n24161 , n23899 );
nand ( n24163 , n24160 , n24162 );
buf ( n24164 , n6493 );
not ( n24165 , n24164 );
and ( n24166 , n24163 , n24165 );
not ( n24167 , n24163 );
buf ( n24168 , n24164 );
and ( n24169 , n24167 , n24168 );
nor ( n24170 , n24166 , n24169 );
buf ( n24171 , n6494 );
nand ( n24172 , n7093 , n24171 );
buf ( n24173 , n6495 );
buf ( n24174 , n24173 );
and ( n24175 , n24172 , n24174 );
not ( n24176 , n24172 );
not ( n24177 , n24173 );
and ( n24178 , n24176 , n24177 );
nor ( n24179 , n24175 , n24178 );
xor ( n24180 , n24170 , n24179 );
xnor ( n24181 , n24180 , n20384 );
not ( n24182 , n24181 );
not ( n24183 , n24182 );
not ( n24184 , n24183 );
or ( n24185 , n24154 , n24184 );
buf ( n24186 , n24181 );
not ( n24187 , n24186 );
nand ( n24188 , n24187 , n15216 );
nand ( n24189 , n24185 , n24188 );
buf ( n24190 , n10696 );
and ( n24191 , n24189 , n24190 );
not ( n24192 , n24189 );
not ( n24193 , n24190 );
and ( n24194 , n24192 , n24193 );
nor ( n24195 , n24191 , n24194 );
nand ( n24196 , n24152 , n24195 );
not ( n24197 , n24196 );
not ( n24198 , n17073 );
not ( n24199 , n13343 );
or ( n24200 , n24198 , n24199 );
or ( n24201 , n13343 , n17073 );
nand ( n24202 , n24200 , n24201 );
not ( n24203 , n21572 );
xor ( n24204 , n24202 , n24203 );
not ( n24205 , n24204 );
and ( n24206 , n24197 , n24205 );
and ( n24207 , n24196 , n24204 );
nor ( n24208 , n24206 , n24207 );
and ( n24209 , n24150 , n24208 );
not ( n24210 , n24150 );
not ( n24211 , n24208 );
and ( n24212 , n24210 , n24211 );
nor ( n24213 , n24209 , n24212 );
not ( n24214 , n24213 );
buf ( n24215 , n18234 );
not ( n24216 , n24215 );
not ( n24217 , n14208 );
or ( n24218 , n24216 , n24217 );
nand ( n24219 , n14213 , n18235 );
nand ( n24220 , n24218 , n24219 );
and ( n24221 , n24220 , n23823 );
not ( n24222 , n24220 );
and ( n24223 , n24222 , n16801 );
nor ( n24224 , n24221 , n24223 );
not ( n24225 , n24224 );
not ( n24226 , n13072 );
not ( n24227 , n24226 );
xor ( n24228 , n22161 , n24227 );
not ( n24229 , n19205 );
xnor ( n24230 , n24228 , n24229 );
not ( n24231 , n24230 );
buf ( n24232 , n18761 );
not ( n24233 , n24232 );
not ( n24234 , n21399 );
or ( n24235 , n24233 , n24234 );
or ( n24236 , n21399 , n24232 );
nand ( n24237 , n24235 , n24236 );
not ( n24238 , n21648 );
not ( n24239 , n24238 );
and ( n24240 , n24237 , n24239 );
not ( n24241 , n24237 );
xor ( n24242 , n21636 , n21645 );
xnor ( n24243 , n24242 , n19509 );
not ( n24244 , n24243 );
not ( n24245 , n24244 );
and ( n24246 , n24241 , n24245 );
nor ( n24247 , n24240 , n24246 );
not ( n24248 , n24247 );
nand ( n24249 , n24231 , n24248 );
not ( n24250 , n24249 );
or ( n24251 , n24225 , n24250 );
not ( n24252 , n24247 );
nand ( n24253 , n24252 , n24231 );
or ( n24254 , n24253 , n24224 );
nand ( n24255 , n24251 , n24254 );
not ( n24256 , n24255 );
not ( n24257 , n7512 );
and ( n24258 , n7518 , n24257 );
not ( n24259 , n7518 );
and ( n24260 , n24259 , n7513 );
nor ( n24261 , n24258 , n24260 );
xor ( n24262 , n24261 , n23444 );
buf ( n24263 , n14970 );
xnor ( n24264 , n24262 , n24263 );
not ( n24265 , n24264 );
not ( n24266 , n21977 );
not ( n24267 , n10872 );
and ( n24268 , n24266 , n24267 );
and ( n24269 , n21977 , n10872 );
nor ( n24270 , n24268 , n24269 );
not ( n24271 , n24270 );
not ( n24272 , n6682 );
or ( n24273 , n24271 , n24272 );
or ( n24274 , n6682 , n24270 );
nand ( n24275 , n24273 , n24274 );
not ( n24276 , n24275 );
nand ( n24277 , n24265 , n24276 );
not ( n24278 , n24277 );
not ( n24279 , n16496 );
not ( n24280 , n12271 );
or ( n24281 , n24279 , n24280 );
or ( n24282 , n12271 , n16496 );
nand ( n24283 , n24281 , n24282 );
and ( n24284 , n24283 , n22895 );
not ( n24285 , n24283 );
not ( n24286 , n22895 );
and ( n24287 , n24285 , n24286 );
nor ( n24288 , n24284 , n24287 );
not ( n24289 , n24288 );
not ( n24290 , n24289 );
and ( n24291 , n24278 , n24290 );
and ( n24292 , n24277 , n24289 );
nor ( n24293 , n24291 , n24292 );
not ( n24294 , n24293 );
or ( n24295 , n24256 , n24294 );
or ( n24296 , n24255 , n24293 );
nand ( n24297 , n24295 , n24296 );
not ( n24298 , n24297 );
and ( n24299 , n24214 , n24298 );
and ( n24300 , n24213 , n24297 );
nor ( n24301 , n24299 , n24300 );
buf ( n24302 , n24301 );
not ( n24303 , n24302 );
and ( n24304 , n24064 , n24303 );
and ( n24305 , n24063 , n24302 );
nor ( n24306 , n24304 , n24305 );
nand ( n24307 , n23819 , n24306 );
not ( n24308 , n10244 );
not ( n24309 , n9776 );
or ( n24310 , n24308 , n24309 );
or ( n24311 , n9776 , n10244 );
nand ( n24312 , n24310 , n24311 );
not ( n24313 , n24312 );
not ( n24314 , n9725 );
or ( n24315 , n24313 , n24314 );
or ( n24316 , n9725 , n24312 );
nand ( n24317 , n24315 , n24316 );
not ( n24318 , n24317 );
not ( n24319 , n6595 );
not ( n24320 , n18930 );
xor ( n24321 , n24320 , n18949 );
not ( n24322 , n18939 );
xnor ( n24323 , n24321 , n24322 );
not ( n24324 , n24323 );
or ( n24325 , n24319 , n24324 );
nand ( n24326 , n18951 , n6598 );
nand ( n24327 , n24325 , n24326 );
not ( n24328 , n24327 );
buf ( n24329 , n18981 );
not ( n24330 , n24329 );
and ( n24331 , n24328 , n24330 );
and ( n24332 , n24327 , n24329 );
nor ( n24333 , n24331 , n24332 );
not ( n24334 , n24333 );
nand ( n24335 , n24318 , n24334 );
and ( n24336 , n19032 , n11503 );
not ( n24337 , n19032 );
and ( n24338 , n24337 , n11502 );
nor ( n24339 , n24336 , n24338 );
and ( n24340 , n24339 , n20218 );
not ( n24341 , n24339 );
not ( n24342 , n20218 );
and ( n24343 , n24341 , n24342 );
nor ( n24344 , n24340 , n24343 );
not ( n24345 , n24344 );
and ( n24346 , n24335 , n24345 );
not ( n24347 , n24335 );
and ( n24348 , n24347 , n24344 );
nor ( n24349 , n24346 , n24348 );
not ( n24350 , n24349 );
not ( n24351 , n24350 );
buf ( n24352 , n21417 );
not ( n24353 , n24352 );
not ( n24354 , n20056 );
or ( n24355 , n24353 , n24354 );
not ( n24356 , n24352 );
nand ( n24357 , n24356 , n20062 );
nand ( n24358 , n24355 , n24357 );
not ( n24359 , n24358 );
not ( n24360 , n16750 );
buf ( n24361 , n6496 );
not ( n24362 , n24361 );
not ( n24363 , n24362 );
or ( n24364 , n24360 , n24363 );
not ( n24365 , n16749 );
buf ( n24366 , n24361 );
nand ( n24367 , n24365 , n24366 );
nand ( n24368 , n24364 , n24367 );
buf ( n24369 , n6497 );
not ( n24370 , n24369 );
and ( n24371 , n24368 , n24370 );
not ( n24372 , n24368 );
buf ( n24373 , n24369 );
and ( n24374 , n24372 , n24373 );
nor ( n24375 , n24371 , n24374 );
buf ( n24376 , n6498 );
nand ( n24377 , n7412 , n24376 );
buf ( n24378 , n6499 );
xor ( n24379 , n24377 , n24378 );
xor ( n24380 , n24375 , n24379 );
buf ( n24381 , n6500 );
nand ( n24382 , n13379 , n24381 );
buf ( n24383 , n6501 );
not ( n24384 , n24383 );
and ( n24385 , n24382 , n24384 );
not ( n24386 , n24382 );
buf ( n24387 , n24383 );
and ( n24388 , n24386 , n24387 );
nor ( n24389 , n24385 , n24388 );
xnor ( n24390 , n24380 , n24389 );
not ( n24391 , n24390 );
not ( n24392 , n24391 );
not ( n24393 , n24392 );
and ( n24394 , n24359 , n24393 );
and ( n24395 , n24358 , n24392 );
nor ( n24396 , n24394 , n24395 );
not ( n24397 , n24396 );
not ( n24398 , n7250 );
not ( n24399 , n19305 );
and ( n24400 , n24398 , n24399 );
and ( n24401 , n7250 , n19305 );
nor ( n24402 , n24400 , n24401 );
not ( n24403 , n24402 );
not ( n24404 , n11176 );
not ( n24405 , n24404 );
or ( n24406 , n24403 , n24405 );
not ( n24407 , n11176 );
or ( n24408 , n24407 , n24402 );
nand ( n24409 , n24406 , n24408 );
not ( n24410 , n24409 );
nand ( n24411 , n24397 , n24410 );
not ( n24412 , n24411 );
not ( n24413 , n15793 );
not ( n24414 , n9313 );
not ( n24415 , n19026 );
or ( n24416 , n24414 , n24415 );
nand ( n24417 , n15830 , n9309 );
nand ( n24418 , n24416 , n24417 );
not ( n24419 , n24418 );
and ( n24420 , n24413 , n24419 );
and ( n24421 , n15793 , n24418 );
nor ( n24422 , n24420 , n24421 );
not ( n24423 , n24422 );
not ( n24424 , n24423 );
and ( n24425 , n24412 , n24424 );
and ( n24426 , n24411 , n24423 );
nor ( n24427 , n24425 , n24426 );
not ( n24428 , n24427 );
not ( n24429 , n24428 );
or ( n24430 , n24351 , n24429 );
nand ( n24431 , n24349 , n24427 );
nand ( n24432 , n24430 , n24431 );
buf ( n24433 , n24432 );
xor ( n24434 , n13093 , n8441 );
xnor ( n24435 , n24434 , n21521 );
not ( n24436 , n23115 );
buf ( n24437 , n17480 );
not ( n24438 , n24437 );
or ( n24439 , n24436 , n24438 );
not ( n24440 , n24437 );
not ( n24441 , n23114 );
nand ( n24442 , n24440 , n24441 );
nand ( n24443 , n24439 , n24442 );
not ( n24444 , n22783 );
and ( n24445 , n24443 , n24444 );
not ( n24446 , n24443 );
not ( n24447 , n22784 );
not ( n24448 , n24447 );
and ( n24449 , n24446 , n24448 );
nor ( n24450 , n24445 , n24449 );
nand ( n24451 , n24435 , n24450 );
not ( n24452 , n24451 );
not ( n24453 , n23781 );
not ( n24454 , n12592 );
or ( n24455 , n24453 , n24454 );
or ( n24456 , n12592 , n23781 );
nand ( n24457 , n24455 , n24456 );
not ( n24458 , n24457 );
not ( n24459 , n12641 );
and ( n24460 , n24458 , n24459 );
and ( n24461 , n24457 , n12641 );
nor ( n24462 , n24460 , n24461 );
not ( n24463 , n24462 );
not ( n24464 , n24463 );
and ( n24465 , n24452 , n24464 );
and ( n24466 , n24451 , n24463 );
nor ( n24467 , n24465 , n24466 );
buf ( n24468 , n24467 );
not ( n24469 , n24468 );
and ( n24470 , n24433 , n24469 );
not ( n24471 , n24433 );
and ( n24472 , n24471 , n24468 );
nor ( n24473 , n24470 , n24472 );
not ( n24474 , n19889 );
not ( n24475 , n13908 );
buf ( n24476 , n6502 );
buf ( n24477 , n24476 );
not ( n24478 , n24477 );
buf ( n24479 , n6503 );
not ( n24480 , n24479 );
not ( n24481 , n24480 );
or ( n24482 , n24478 , n24481 );
not ( n24483 , n24476 );
buf ( n24484 , n24479 );
nand ( n24485 , n24483 , n24484 );
nand ( n24486 , n24482 , n24485 );
buf ( n24487 , n6504 );
buf ( n24488 , n24487 );
and ( n24489 , n24486 , n24488 );
not ( n24490 , n24486 );
not ( n24491 , n24487 );
and ( n24492 , n24490 , n24491 );
nor ( n24493 , n24489 , n24492 );
buf ( n24494 , n6505 );
nand ( n24495 , n8740 , n24494 );
buf ( n24496 , n6506 );
buf ( n24497 , n24496 );
and ( n24498 , n24495 , n24497 );
not ( n24499 , n24495 );
not ( n24500 , n24496 );
and ( n24501 , n24499 , n24500 );
nor ( n24502 , n24498 , n24501 );
xor ( n24503 , n24493 , n24502 );
buf ( n24504 , n6507 );
nand ( n24505 , n7617 , n24504 );
buf ( n24506 , n6508 );
buf ( n24507 , n24506 );
and ( n24508 , n24505 , n24507 );
not ( n24509 , n24505 );
not ( n24510 , n24506 );
and ( n24511 , n24509 , n24510 );
nor ( n24512 , n24508 , n24511 );
xnor ( n24513 , n24503 , n24512 );
buf ( n24514 , n24513 );
not ( n24515 , n24514 );
or ( n24516 , n24475 , n24515 );
buf ( n24517 , n24514 );
or ( n24518 , n24517 , n13908 );
nand ( n24519 , n24516 , n24518 );
not ( n24520 , n24519 );
and ( n24521 , n24474 , n24520 );
not ( n24522 , n19888 );
and ( n24523 , n24522 , n24519 );
nor ( n24524 , n24521 , n24523 );
not ( n24525 , n7603 );
not ( n24526 , n18000 );
or ( n24527 , n24525 , n24526 );
nand ( n24528 , n10942 , n7600 );
nand ( n24529 , n24527 , n24528 );
and ( n24530 , n24529 , n19393 );
not ( n24531 , n24529 );
and ( n24532 , n24531 , n19392 );
nor ( n24533 , n24530 , n24532 );
nand ( n24534 , n24524 , n24533 );
not ( n24535 , n15958 );
not ( n24536 , n19492 );
or ( n24537 , n24535 , n24536 );
nand ( n24538 , n23721 , n15954 );
nand ( n24539 , n24537 , n24538 );
and ( n24540 , n24539 , n13256 );
not ( n24541 , n24539 );
and ( n24542 , n24541 , n12804 );
nor ( n24543 , n24540 , n24542 );
not ( n24544 , n24543 );
and ( n24545 , n24534 , n24544 );
not ( n24546 , n24534 );
and ( n24547 , n24546 , n24543 );
nor ( n24548 , n24545 , n24547 );
not ( n24549 , n24548 );
xor ( n24550 , n18161 , n23705 );
buf ( n24551 , n8329 );
xnor ( n24552 , n24550 , n24551 );
buf ( n24553 , n18072 );
not ( n24554 , n24553 );
not ( n24555 , n17390 );
or ( n24556 , n24554 , n24555 );
or ( n24557 , n17390 , n24553 );
nand ( n24558 , n24556 , n24557 );
and ( n24559 , n24558 , n17396 );
not ( n24560 , n24558 );
and ( n24561 , n24560 , n17397 );
nor ( n24562 , n24559 , n24561 );
nand ( n24563 , n24552 , n24562 );
not ( n24564 , n24563 );
not ( n24565 , n11680 );
not ( n24566 , n10376 );
or ( n24567 , n24565 , n24566 );
or ( n24568 , n14494 , n11680 );
nand ( n24569 , n24567 , n24568 );
and ( n24570 , n24569 , n14521 );
not ( n24571 , n24569 );
and ( n24572 , n24571 , n14522 );
nor ( n24573 , n24570 , n24572 );
not ( n24574 , n24573 );
and ( n24575 , n24564 , n24574 );
nand ( n24576 , n24562 , n24552 );
and ( n24577 , n24576 , n24573 );
nor ( n24578 , n24575 , n24577 );
not ( n24579 , n24578 );
or ( n24580 , n24549 , n24579 );
or ( n24581 , n24578 , n24548 );
nand ( n24582 , n24580 , n24581 );
buf ( n24583 , n24582 );
not ( n24584 , n24583 );
and ( n24585 , n24473 , n24584 );
not ( n24586 , n24473 );
and ( n24587 , n24586 , n24583 );
nor ( n24588 , n24585 , n24587 );
buf ( n24589 , n24588 );
not ( n24590 , n24589 );
not ( n24591 , n10425 );
not ( n24592 , n22984 );
or ( n24593 , n24591 , n24592 );
or ( n24594 , n22984 , n10425 );
nand ( n24595 , n24593 , n24594 );
not ( n24596 , n20564 );
and ( n24597 , n24595 , n24596 );
not ( n24598 , n24595 );
and ( n24599 , n24598 , n20564 );
nor ( n24600 , n24597 , n24599 );
not ( n24601 , n11122 );
not ( n24602 , n18737 );
or ( n24603 , n24601 , n24602 );
buf ( n24604 , n10117 );
nand ( n24605 , n24604 , n11117 );
nand ( n24606 , n24603 , n24605 );
and ( n24607 , n24606 , n10170 );
not ( n24608 , n24606 );
and ( n24609 , n24608 , n20136 );
nor ( n24610 , n24607 , n24609 );
not ( n24611 , n24610 );
nand ( n24612 , n24600 , n24611 );
not ( n24613 , n24612 );
buf ( n24614 , n8759 );
xor ( n24615 , n24614 , n19282 );
xor ( n24616 , n20479 , n20498 );
not ( n24617 , n20488 );
xnor ( n24618 , n24616 , n24617 );
not ( n24619 , n24618 );
not ( n24620 , n24619 );
xor ( n24621 , n24615 , n24620 );
not ( n24622 , n24621 );
not ( n24623 , n24622 );
not ( n24624 , n24623 );
and ( n24625 , n24613 , n24624 );
and ( n24626 , n24612 , n24623 );
nor ( n24627 , n24625 , n24626 );
not ( n24628 , n24627 );
buf ( n24629 , n11047 );
not ( n24630 , n24629 );
not ( n24631 , n18906 );
or ( n24632 , n24630 , n24631 );
or ( n24633 , n18906 , n24629 );
nand ( n24634 , n24632 , n24633 );
not ( n24635 , n24634 );
not ( n24636 , n13015 );
and ( n24637 , n24635 , n24636 );
buf ( n24638 , n7933 );
and ( n24639 , n24634 , n24638 );
nor ( n24640 , n24637 , n24639 );
not ( n24641 , n24640 );
not ( n24642 , n24641 );
not ( n24643 , n24600 );
nand ( n24644 , n24622 , n24643 );
not ( n24645 , n24644 );
or ( n24646 , n24642 , n24645 );
or ( n24647 , n24644 , n24641 );
nand ( n24648 , n24646 , n24647 );
not ( n24649 , n24648 );
not ( n24650 , n24649 );
not ( n24651 , n18415 );
buf ( n24652 , n6509 );
not ( n24653 , n24652 );
not ( n24654 , n24653 );
or ( n24655 , n24651 , n24654 );
not ( n24656 , n18414 );
buf ( n24657 , n24652 );
nand ( n24658 , n24656 , n24657 );
nand ( n24659 , n24655 , n24658 );
not ( n24660 , n14759 );
and ( n24661 , n24659 , n24660 );
not ( n24662 , n24659 );
and ( n24663 , n24662 , n14760 );
nor ( n24664 , n24661 , n24663 );
buf ( n24665 , n6510 );
nand ( n24666 , n7133 , n24665 );
buf ( n24667 , n6511 );
buf ( n24668 , n24667 );
and ( n24669 , n24666 , n24668 );
not ( n24670 , n24666 );
not ( n24671 , n24667 );
and ( n24672 , n24670 , n24671 );
nor ( n24673 , n24669 , n24672 );
xor ( n24674 , n24664 , n24673 );
buf ( n24675 , n6512 );
nand ( n24676 , n6608 , n24675 );
buf ( n24677 , n6513 );
not ( n24678 , n24677 );
and ( n24679 , n24676 , n24678 );
not ( n24680 , n24676 );
buf ( n24681 , n24677 );
and ( n24682 , n24680 , n24681 );
nor ( n24683 , n24679 , n24682 );
xor ( n24684 , n24674 , n24683 );
not ( n24685 , n24684 );
not ( n24686 , n24685 );
buf ( n24687 , n24686 );
xor ( n24688 , n14335 , n24687 );
buf ( n24689 , n6514 );
buf ( n24690 , n6515 );
buf ( n24691 , n24690 );
not ( n24692 , n24691 );
buf ( n24693 , n6516 );
not ( n24694 , n24693 );
not ( n24695 , n24694 );
or ( n24696 , n24692 , n24695 );
not ( n24697 , n24690 );
buf ( n24698 , n24693 );
nand ( n24699 , n24697 , n24698 );
nand ( n24700 , n24696 , n24699 );
xor ( n24701 , n24689 , n24700 );
buf ( n24702 , n6517 );
buf ( n24703 , n6518 );
not ( n24704 , n24703 );
xor ( n24705 , n24702 , n24704 );
buf ( n24706 , n6519 );
nand ( n24707 , n6608 , n24706 );
xnor ( n24708 , n24705 , n24707 );
xnor ( n24709 , n24701 , n24708 );
buf ( n24710 , n24709 );
not ( n24711 , n24710 );
xnor ( n24712 , n24688 , n24711 );
not ( n24713 , n24712 );
not ( n24714 , n18038 );
not ( n24715 , n14430 );
or ( n24716 , n24714 , n24715 );
or ( n24717 , n14430 , n18038 );
nand ( n24718 , n24716 , n24717 );
and ( n24719 , n24718 , n21227 );
not ( n24720 , n24718 );
and ( n24721 , n24720 , n20518 );
nor ( n24722 , n24719 , n24721 );
nand ( n24723 , n24713 , n24722 );
not ( n24724 , n24723 );
buf ( n24725 , n14514 );
and ( n24726 , n14518 , n24725 );
not ( n24727 , n14518 );
and ( n24728 , n24727 , n14515 );
nor ( n24729 , n24726 , n24728 );
xor ( n24730 , n24729 , n12465 );
not ( n24731 , n24730 );
buf ( n24732 , n21795 );
not ( n24733 , n24732 );
buf ( n24734 , n6520 );
not ( n24735 , n24734 );
not ( n24736 , n24735 );
or ( n24737 , n24733 , n24736 );
buf ( n24738 , n24734 );
nand ( n24739 , n21796 , n24738 );
nand ( n24740 , n24737 , n24739 );
buf ( n24741 , n6521 );
buf ( n24742 , n24741 );
and ( n24743 , n24740 , n24742 );
not ( n24744 , n24740 );
not ( n24745 , n24741 );
and ( n24746 , n24744 , n24745 );
nor ( n24747 , n24743 , n24746 );
xor ( n24748 , n24747 , n18678 );
buf ( n24749 , n6522 );
nand ( n24750 , n7617 , n24749 );
buf ( n24751 , n6523 );
not ( n24752 , n24751 );
and ( n24753 , n24750 , n24752 );
not ( n24754 , n24750 );
buf ( n24755 , n24751 );
and ( n24756 , n24754 , n24755 );
nor ( n24757 , n24753 , n24756 );
xnor ( n24758 , n24748 , n24757 );
not ( n24759 , n24758 );
not ( n24760 , n24759 );
and ( n24761 , n24731 , n24760 );
not ( n24762 , n24759 );
not ( n24763 , n24762 );
and ( n24764 , n24730 , n24763 );
nor ( n24765 , n24761 , n24764 );
not ( n24766 , n24765 );
not ( n24767 , n24766 );
and ( n24768 , n24724 , n24767 );
and ( n24769 , n24723 , n24766 );
nor ( n24770 , n24768 , n24769 );
not ( n24771 , n24770 );
not ( n24772 , n24771 );
or ( n24773 , n24650 , n24772 );
nand ( n24774 , n24770 , n24648 );
nand ( n24775 , n24773 , n24774 );
not ( n24776 , n24775 );
not ( n24777 , n24776 );
not ( n24778 , n11778 );
not ( n24779 , n14113 );
not ( n24780 , n6715 );
and ( n24781 , n24779 , n24780 );
not ( n24782 , n14920 );
and ( n24783 , n14113 , n24782 );
nor ( n24784 , n24781 , n24783 );
not ( n24785 , n24784 );
or ( n24786 , n24778 , n24785 );
or ( n24787 , n24784 , n11778 );
nand ( n24788 , n24786 , n24787 );
not ( n24789 , n24788 );
buf ( n24790 , n6524 );
buf ( n24791 , n24790 );
not ( n24792 , n24791 );
buf ( n24793 , n6525 );
not ( n24794 , n24793 );
not ( n24795 , n24794 );
or ( n24796 , n24792 , n24795 );
not ( n24797 , n24790 );
buf ( n24798 , n24793 );
nand ( n24799 , n24797 , n24798 );
nand ( n24800 , n24796 , n24799 );
not ( n24801 , n23727 );
and ( n24802 , n24800 , n24801 );
not ( n24803 , n24800 );
and ( n24804 , n24803 , n23728 );
nor ( n24805 , n24802 , n24804 );
buf ( n24806 , n6526 );
nand ( n24807 , n6706 , n24806 );
buf ( n24808 , n6527 );
buf ( n24809 , n24808 );
and ( n24810 , n24807 , n24809 );
not ( n24811 , n24807 );
not ( n24812 , n24808 );
and ( n24813 , n24811 , n24812 );
nor ( n24814 , n24810 , n24813 );
xor ( n24815 , n24805 , n24814 );
buf ( n24816 , n6528 );
nand ( n24817 , n6863 , n24816 );
buf ( n24818 , n6529 );
buf ( n24819 , n24818 );
and ( n24820 , n24817 , n24819 );
not ( n24821 , n24817 );
not ( n24822 , n24818 );
and ( n24823 , n24821 , n24822 );
nor ( n24824 , n24820 , n24823 );
not ( n24825 , n24824 );
xor ( n24826 , n24815 , n24825 );
not ( n24827 , n24826 );
not ( n24828 , n24827 );
not ( n24829 , n10825 );
and ( n24830 , n24828 , n24829 );
xor ( n24831 , n24805 , n24824 );
not ( n24832 , n24814 );
xor ( n24833 , n24831 , n24832 );
not ( n24834 , n24833 );
and ( n24835 , n24834 , n10825 );
nor ( n24836 , n24830 , n24835 );
buf ( n24837 , n6530 );
buf ( n24838 , n24837 );
not ( n24839 , n24838 );
buf ( n24840 , n6531 );
not ( n24841 , n24840 );
not ( n24842 , n24841 );
or ( n24843 , n24839 , n24842 );
not ( n24844 , n24837 );
buf ( n24845 , n24840 );
nand ( n24846 , n24844 , n24845 );
nand ( n24847 , n24843 , n24846 );
buf ( n24848 , n6532 );
not ( n24849 , n24848 );
and ( n24850 , n24847 , n24849 );
not ( n24851 , n24847 );
buf ( n24852 , n24848 );
and ( n24853 , n24851 , n24852 );
nor ( n24854 , n24850 , n24853 );
buf ( n24855 , n6533 );
nand ( n24856 , n6660 , n24855 );
buf ( n24857 , n6534 );
buf ( n24858 , n24857 );
and ( n24859 , n24856 , n24858 );
not ( n24860 , n24856 );
not ( n24861 , n24857 );
and ( n24862 , n24860 , n24861 );
nor ( n24863 , n24859 , n24862 );
xor ( n24864 , n24854 , n24863 );
buf ( n24865 , n6535 );
nand ( n24866 , n6608 , n24865 );
buf ( n24867 , n6536 );
buf ( n24868 , n24867 );
and ( n24869 , n24866 , n24868 );
not ( n24870 , n24866 );
not ( n24871 , n24867 );
and ( n24872 , n24870 , n24871 );
nor ( n24873 , n24869 , n24872 );
xnor ( n24874 , n24864 , n24873 );
buf ( n24875 , n24874 );
not ( n24876 , n24875 );
and ( n24877 , n24836 , n24876 );
not ( n24878 , n24836 );
not ( n24879 , n24875 );
not ( n24880 , n24879 );
buf ( n24881 , n24880 );
and ( n24882 , n24878 , n24881 );
nor ( n24883 , n24877 , n24882 );
nand ( n24884 , n24789 , n24883 );
not ( n24885 , n24884 );
not ( n24886 , n6632 );
not ( n24887 , n18951 );
or ( n24888 , n24886 , n24887 );
or ( n24889 , n18951 , n6632 );
nand ( n24890 , n24888 , n24889 );
xor ( n24891 , n24890 , n24329 );
not ( n24892 , n24891 );
not ( n24893 , n24892 );
and ( n24894 , n24885 , n24893 );
and ( n24895 , n24884 , n24892 );
nor ( n24896 , n24894 , n24895 );
not ( n24897 , n24896 );
not ( n24898 , n8287 );
not ( n24899 , n24898 );
not ( n24900 , n19025 );
not ( n24901 , n24900 );
not ( n24902 , n14533 );
or ( n24903 , n24901 , n24902 );
or ( n24904 , n14533 , n24900 );
nand ( n24905 , n24903 , n24904 );
not ( n24906 , n24905 );
and ( n24907 , n24899 , n24906 );
and ( n24908 , n8238 , n24905 );
nor ( n24909 , n24907 , n24908 );
not ( n24910 , n21853 );
not ( n24911 , n8440 );
or ( n24912 , n24910 , n24911 );
nand ( n24913 , n8433 , n21849 );
nand ( n24914 , n24912 , n24913 );
not ( n24915 , n24914 );
not ( n24916 , n9689 );
and ( n24917 , n24915 , n24916 );
and ( n24918 , n24914 , n9689 );
nor ( n24919 , n24917 , n24918 );
not ( n24920 , n24919 );
nand ( n24921 , n24909 , n24920 );
buf ( n24922 , n12146 );
and ( n24923 , n24922 , n11058 );
not ( n24924 , n24922 );
and ( n24925 , n24924 , n21201 );
nor ( n24926 , n24923 , n24925 );
not ( n24927 , n24926 );
not ( n24928 , n24927 );
not ( n24929 , n11061 );
or ( n24930 , n24928 , n24929 );
nand ( n24931 , n8612 , n24926 );
nand ( n24932 , n24930 , n24931 );
not ( n24933 , n24932 );
and ( n24934 , n24921 , n24933 );
not ( n24935 , n24921 );
and ( n24936 , n24935 , n24932 );
nor ( n24937 , n24934 , n24936 );
not ( n24938 , n24937 );
or ( n24939 , n24897 , n24938 );
or ( n24940 , n24937 , n24896 );
nand ( n24941 , n24939 , n24940 );
not ( n24942 , n19931 );
and ( n24943 , n17451 , n7969 );
not ( n24944 , n17451 );
and ( n24945 , n24944 , n7976 );
nor ( n24946 , n24943 , n24945 );
not ( n24947 , n24946 );
not ( n24948 , n24947 );
or ( n24949 , n24942 , n24948 );
nand ( n24950 , n24946 , n19923 );
nand ( n24951 , n24949 , n24950 );
not ( n24952 , n9544 );
not ( n24953 , n12230 );
not ( n24954 , n9532 );
or ( n24955 , n24953 , n24954 );
or ( n24956 , n9532 , n12230 );
nand ( n24957 , n24955 , n24956 );
not ( n24958 , n24957 );
or ( n24959 , n24952 , n24958 );
or ( n24960 , n24957 , n24085 );
nand ( n24961 , n24959 , n24960 );
not ( n24962 , n24961 );
nand ( n24963 , n24951 , n24962 );
buf ( n24964 , n13444 );
not ( n24965 , n24964 );
xor ( n24966 , n11447 , n11466 );
not ( n24967 , n11456 );
xnor ( n24968 , n24966 , n24967 );
not ( n24969 , n24968 );
or ( n24970 , n24965 , n24969 );
or ( n24971 , n24968 , n24964 );
nand ( n24972 , n24970 , n24971 );
xnor ( n24973 , n24972 , n22215 );
not ( n24974 , n24973 );
xor ( n24975 , n24963 , n24974 );
not ( n24976 , n24975 );
and ( n24977 , n24941 , n24976 );
not ( n24978 , n24941 );
and ( n24979 , n24978 , n24975 );
nor ( n24980 , n24977 , n24979 );
not ( n24981 , n24980 );
not ( n24982 , n24981 );
or ( n24983 , n24777 , n24982 );
nand ( n24984 , n24980 , n24775 );
nand ( n24985 , n24983 , n24984 );
not ( n24986 , n24985 );
or ( n24987 , n24628 , n24986 );
and ( n24988 , n24980 , n24775 );
not ( n24989 , n24980 );
and ( n24990 , n24989 , n24776 );
nor ( n24991 , n24988 , n24990 );
not ( n24992 , n24627 );
nand ( n24993 , n24991 , n24992 );
nand ( n24994 , n24987 , n24993 );
not ( n24995 , n24994 );
and ( n24996 , n24590 , n24995 );
and ( n24997 , n24589 , n24994 );
nor ( n24998 , n24996 , n24997 );
not ( n24999 , n24998 );
buf ( n25000 , n13743 );
buf ( n25001 , n25000 );
nor ( n25002 , n24999 , n25001 );
not ( n25003 , n25002 );
or ( n25004 , n24307 , n25003 );
nor ( n25005 , n24998 , n25001 );
nand ( n25006 , n24307 , n25005 );
buf ( n25007 , n13766 );
nand ( n25008 , n25007 , n16293 );
nand ( n25009 , n25004 , n25006 , n25008 );
buf ( n25010 , n25009 );
buf ( n25011 , n25010 );
buf ( n25012 , n19764 );
not ( n25013 , n25012 );
not ( n25014 , n25013 );
not ( n25015 , n11284 );
or ( n25016 , n25014 , n25015 );
nand ( n25017 , n11287 , n25012 );
nand ( n25018 , n25016 , n25017 );
buf ( n25019 , n7053 );
not ( n25020 , n25019 );
and ( n25021 , n25018 , n25020 );
not ( n25022 , n25018 );
and ( n25023 , n25022 , n25019 );
nor ( n25024 , n25021 , n25023 );
not ( n25025 , n25024 );
nand ( n25026 , n13502 , n25025 );
not ( n25027 , n25026 );
not ( n25028 , n15875 );
not ( n25029 , n10844 );
or ( n25030 , n25028 , n25029 );
not ( n25031 , n15875 );
nand ( n25032 , n25031 , n23640 );
nand ( n25033 , n25030 , n25032 );
buf ( n25034 , n8150 );
and ( n25035 , n25033 , n25034 );
not ( n25036 , n25033 );
and ( n25037 , n25036 , n22289 );
nor ( n25038 , n25035 , n25037 );
not ( n25039 , n25038 );
not ( n25040 , n25039 );
not ( n25041 , n25040 );
and ( n25042 , n25027 , n25041 );
and ( n25043 , n25026 , n25040 );
nor ( n25044 , n25042 , n25043 );
buf ( n25045 , n25044 );
not ( n25046 , n25045 );
not ( n25047 , n9542 );
not ( n25048 , n25047 );
buf ( n25049 , n19777 );
xor ( n25050 , n25049 , n19787 );
xnor ( n25051 , n25050 , n19803 );
not ( n25052 , n25051 );
not ( n25053 , n25052 );
or ( n25054 , n25048 , n25053 );
not ( n25055 , n25047 );
nand ( n25056 , n25055 , n25051 );
nand ( n25057 , n25054 , n25056 );
xor ( n25058 , n19760 , n19764 );
xor ( n25059 , n25058 , n19774 );
not ( n25060 , n25059 );
and ( n25061 , n25057 , n25060 );
not ( n25062 , n25057 );
buf ( n25063 , n25059 );
and ( n25064 , n25062 , n25063 );
nor ( n25065 , n25061 , n25064 );
not ( n25066 , n8954 );
xor ( n25067 , n20611 , n20620 );
xnor ( n25068 , n25067 , n20630 );
not ( n25069 , n25068 );
or ( n25070 , n25066 , n25069 );
or ( n25071 , n25068 , n8954 );
nand ( n25072 , n25070 , n25071 );
xnor ( n25073 , n25072 , n14342 );
nand ( n25074 , n25065 , n25073 );
not ( n25075 , n25074 );
buf ( n25076 , n12963 );
not ( n25077 , n25076 );
and ( n25078 , n25075 , n25077 );
and ( n25079 , n25074 , n25076 );
nor ( n25080 , n25078 , n25079 );
not ( n25081 , n25080 );
buf ( n25082 , n7868 );
xor ( n25083 , n25082 , n11228 );
and ( n25084 , n25083 , n20940 );
not ( n25085 , n25083 );
and ( n25086 , n25085 , n20941 );
nor ( n25087 , n25084 , n25086 );
not ( n25088 , n11948 );
buf ( n25089 , n6537 );
buf ( n25090 , n25089 );
not ( n25091 , n25090 );
and ( n25092 , n25088 , n25091 );
and ( n25093 , n11948 , n25090 );
nor ( n25094 , n25092 , n25093 );
and ( n25095 , n25094 , n16737 );
not ( n25096 , n25094 );
buf ( n25097 , n11996 );
and ( n25098 , n25096 , n25097 );
nor ( n25099 , n25095 , n25098 );
not ( n25100 , n25099 );
nand ( n25101 , n25087 , n25100 );
buf ( n25102 , n13033 );
xor ( n25103 , n25101 , n25102 );
not ( n25104 , n25103 );
or ( n25105 , n25081 , n25104 );
or ( n25106 , n25080 , n25103 );
nand ( n25107 , n25105 , n25106 );
not ( n25108 , n8847 );
not ( n25109 , n9441 );
and ( n25110 , n25108 , n25109 );
not ( n25111 , n19353 );
and ( n25112 , n25111 , n9441 );
nor ( n25113 , n25110 , n25112 );
not ( n25114 , n8889 );
and ( n25115 , n25113 , n25114 );
not ( n25116 , n25113 );
and ( n25117 , n25116 , n8888 );
nor ( n25118 , n25115 , n25117 );
not ( n25119 , n25118 );
not ( n25120 , n15547 );
not ( n25121 , n7310 );
not ( n25122 , n25121 );
or ( n25123 , n25120 , n25122 );
not ( n25124 , n15547 );
nand ( n25125 , n25124 , n7310 );
nand ( n25126 , n25123 , n25125 );
not ( n25127 , n9532 );
not ( n25128 , n25127 );
xor ( n25129 , n25126 , n25128 );
not ( n25130 , n25129 );
nand ( n25131 , n25119 , n25130 );
not ( n25132 , n13225 );
and ( n25133 , n25131 , n25132 );
not ( n25134 , n25131 );
and ( n25135 , n25134 , n13225 );
nor ( n25136 , n25133 , n25135 );
and ( n25137 , n25107 , n25136 );
not ( n25138 , n25107 );
not ( n25139 , n25136 );
and ( n25140 , n25138 , n25139 );
nor ( n25141 , n25137 , n25140 );
not ( n25142 , n13713 );
not ( n25143 , n25142 );
not ( n25144 , n15712 );
not ( n25145 , n18286 );
or ( n25146 , n25144 , n25145 );
or ( n25147 , n19523 , n15712 );
nand ( n25148 , n25146 , n25147 );
nor ( n25149 , n25148 , n18299 );
not ( n25150 , n25149 );
nand ( n25151 , n25148 , n18299 );
nand ( n25152 , n25150 , n25151 );
not ( n25153 , n25152 );
not ( n25154 , n10492 );
not ( n25155 , n10489 );
and ( n25156 , n25154 , n25155 );
and ( n25157 , n10492 , n10489 );
nor ( n25158 , n25156 , n25157 );
xor ( n25159 , n25158 , n14056 );
xnor ( n25160 , n25159 , n8074 );
not ( n25161 , n25160 );
nand ( n25162 , n25153 , n25161 );
not ( n25163 , n25162 );
or ( n25164 , n25143 , n25163 );
not ( n25165 , n25152 );
nand ( n25166 , n25165 , n25161 );
or ( n25167 , n25166 , n25142 );
nand ( n25168 , n25164 , n25167 );
not ( n25169 , n25168 );
nand ( n25170 , n25039 , n25024 );
not ( n25171 , n25170 );
buf ( n25172 , n13406 );
not ( n25173 , n25172 );
and ( n25174 , n25171 , n25173 );
and ( n25175 , n25170 , n25172 );
nor ( n25176 , n25174 , n25175 );
not ( n25177 , n25176 );
and ( n25178 , n25169 , n25177 );
and ( n25179 , n25168 , n25176 );
nor ( n25180 , n25178 , n25179 );
and ( n25181 , n25141 , n25180 );
not ( n25182 , n25141 );
not ( n25183 , n25180 );
and ( n25184 , n25182 , n25183 );
or ( n25185 , n25181 , n25184 );
not ( n25186 , n25185 );
or ( n25187 , n25046 , n25186 );
and ( n25188 , n25141 , n25180 );
not ( n25189 , n25141 );
and ( n25190 , n25189 , n25183 );
nor ( n25191 , n25188 , n25190 );
not ( n25192 , n25191 );
or ( n25193 , n25192 , n25045 );
nand ( n25194 , n25187 , n25193 );
not ( n25195 , n25194 );
buf ( n25196 , n11316 );
not ( n25197 , n25196 );
not ( n25198 , n11313 );
and ( n25199 , n25197 , n25198 );
and ( n25200 , n25196 , n11313 );
nor ( n25201 , n25199 , n25200 );
buf ( n25202 , n23916 );
xor ( n25203 , n25201 , n25202 );
xnor ( n25204 , n25203 , n7886 );
buf ( n25205 , n25204 );
not ( n25206 , n25205 );
buf ( n25207 , n6538 );
nand ( n25208 , n7288 , n25207 );
buf ( n25209 , n6539 );
not ( n25210 , n25209 );
and ( n25211 , n25208 , n25210 );
not ( n25212 , n25208 );
buf ( n25213 , n25209 );
and ( n25214 , n25212 , n25213 );
nor ( n25215 , n25211 , n25214 );
buf ( n25216 , n6540 );
buf ( n25217 , n25216 );
not ( n25218 , n25217 );
buf ( n25219 , n6541 );
not ( n25220 , n25219 );
not ( n25221 , n25220 );
or ( n25222 , n25218 , n25221 );
not ( n25223 , n25216 );
buf ( n25224 , n25219 );
nand ( n25225 , n25223 , n25224 );
nand ( n25226 , n25222 , n25225 );
buf ( n25227 , n6542 );
buf ( n25228 , n25227 );
and ( n25229 , n25226 , n25228 );
not ( n25230 , n25226 );
not ( n25231 , n25227 );
and ( n25232 , n25230 , n25231 );
nor ( n25233 , n25229 , n25232 );
buf ( n25234 , n6543 );
nand ( n25235 , n7981 , n25234 );
buf ( n25236 , n6544 );
buf ( n25237 , n25236 );
and ( n25238 , n25235 , n25237 );
not ( n25239 , n25235 );
not ( n25240 , n25236 );
and ( n25241 , n25239 , n25240 );
nor ( n25242 , n25238 , n25241 );
xor ( n25243 , n25233 , n25242 );
buf ( n25244 , n6545 );
nand ( n25245 , n8740 , n25244 );
buf ( n25246 , n6546 );
not ( n25247 , n25246 );
and ( n25248 , n25245 , n25247 );
not ( n25249 , n25245 );
buf ( n25250 , n25246 );
and ( n25251 , n25249 , n25250 );
nor ( n25252 , n25248 , n25251 );
xor ( n25253 , n25243 , n25252 );
not ( n25254 , n25253 );
buf ( n25255 , n25254 );
xor ( n25256 , n25215 , n25255 );
xnor ( n25257 , n25256 , n19392 );
not ( n25258 , n25257 );
not ( n25259 , n20095 );
not ( n25260 , n14981 );
not ( n25261 , n18645 );
or ( n25262 , n25260 , n25261 );
or ( n25263 , n18645 , n14981 );
nand ( n25264 , n25262 , n25263 );
not ( n25265 , n25264 );
and ( n25266 , n25259 , n25265 );
and ( n25267 , n20095 , n25264 );
nor ( n25268 , n25266 , n25267 );
not ( n25269 , n25268 );
nand ( n25270 , n25258 , n25269 );
not ( n25271 , n25270 );
or ( n25272 , n25206 , n25271 );
or ( n25273 , n25270 , n25205 );
nand ( n25274 , n25272 , n25273 );
not ( n25275 , n25274 );
xor ( n25276 , n11467 , n13391 );
xnor ( n25277 , n25276 , n18138 );
not ( n25278 , n25277 );
xor ( n25279 , n11893 , n10498 );
xnor ( n25280 , n25279 , n9725 );
not ( n25281 , n25280 );
nand ( n25282 , n25278 , n25281 );
not ( n25283 , n25282 );
buf ( n25284 , n9466 );
not ( n25285 , n25284 );
not ( n25286 , n19353 );
or ( n25287 , n25285 , n25286 );
or ( n25288 , n19353 , n25284 );
nand ( n25289 , n25287 , n25288 );
and ( n25290 , n25289 , n8889 );
not ( n25291 , n25289 );
and ( n25292 , n25291 , n19943 );
nor ( n25293 , n25290 , n25292 );
not ( n25294 , n25293 );
and ( n25295 , n25283 , n25294 );
and ( n25296 , n25282 , n25293 );
nor ( n25297 , n25295 , n25296 );
not ( n25298 , n25297 );
or ( n25299 , n25275 , n25298 );
not ( n25300 , n25274 );
not ( n25301 , n25297 );
nand ( n25302 , n25300 , n25301 );
nand ( n25303 , n25299 , n25302 );
not ( n25304 , n15736 );
not ( n25305 , n18286 );
or ( n25306 , n25304 , n25305 );
not ( n25307 , n15736 );
nand ( n25308 , n25307 , n18293 );
nand ( n25309 , n25306 , n25308 );
not ( n25310 , n25309 );
not ( n25311 , n18299 );
and ( n25312 , n25310 , n25311 );
buf ( n25313 , n18247 );
and ( n25314 , n25313 , n25309 );
nor ( n25315 , n25312 , n25314 );
not ( n25316 , n23572 );
nor ( n25317 , n17208 , n16576 );
not ( n25318 , n25317 );
nand ( n25319 , n17208 , n16576 );
nand ( n25320 , n25318 , n25319 );
not ( n25321 , n25320 );
or ( n25322 , n25316 , n25321 );
or ( n25323 , n25320 , n23572 );
nand ( n25324 , n25322 , n25323 );
nand ( n25325 , n25315 , n25324 );
not ( n25326 , n21095 );
not ( n25327 , n6828 );
or ( n25328 , n25326 , n25327 );
not ( n25329 , n21095 );
nand ( n25330 , n25329 , n23705 );
nand ( n25331 , n25328 , n25330 );
and ( n25332 , n25331 , n23847 );
not ( n25333 , n25331 );
and ( n25334 , n25333 , n6877 );
nor ( n25335 , n25332 , n25334 );
and ( n25336 , n25325 , n25335 );
not ( n25337 , n25325 );
not ( n25338 , n25335 );
and ( n25339 , n25337 , n25338 );
nor ( n25340 , n25336 , n25339 );
not ( n25341 , n25340 );
not ( n25342 , n25341 );
buf ( n25343 , n21954 );
not ( n25344 , n25343 );
not ( n25345 , n13030 );
or ( n25346 , n25344 , n25345 );
or ( n25347 , n10640 , n25343 );
nand ( n25348 , n25346 , n25347 );
and ( n25349 , n25348 , n18793 );
not ( n25350 , n25348 );
not ( n25351 , n18793 );
and ( n25352 , n25350 , n25351 );
nor ( n25353 , n25349 , n25352 );
not ( n25354 , n25353 );
not ( n25355 , n12163 );
not ( n25356 , n21201 );
or ( n25357 , n25355 , n25356 );
or ( n25358 , n21201 , n12163 );
nand ( n25359 , n25357 , n25358 );
not ( n25360 , n25359 );
not ( n25361 , n19645 );
and ( n25362 , n25360 , n25361 );
and ( n25363 , n25359 , n19645 );
nor ( n25364 , n25362 , n25363 );
not ( n25365 , n25364 );
nand ( n25366 , n25354 , n25365 );
not ( n25367 , n25366 );
not ( n25368 , n7010 );
not ( n25369 , n9480 );
xor ( n25370 , n20442 , n25369 );
xnor ( n25371 , n25370 , n9487 );
not ( n25372 , n25371 );
or ( n25373 , n25368 , n25372 );
or ( n25374 , n25371 , n7010 );
nand ( n25375 , n25373 , n25374 );
and ( n25376 , n25375 , n21214 );
not ( n25377 , n25375 );
and ( n25378 , n25377 , n9468 );
nor ( n25379 , n25376 , n25378 );
not ( n25380 , n25379 );
not ( n25381 , n25380 );
and ( n25382 , n25367 , n25381 );
not ( n25383 , n25353 );
nand ( n25384 , n25383 , n25365 );
and ( n25385 , n25384 , n25380 );
nor ( n25386 , n25382 , n25385 );
not ( n25387 , n25386 );
not ( n25388 , n25387 );
or ( n25389 , n25342 , n25388 );
nand ( n25390 , n25386 , n25340 );
nand ( n25391 , n25389 , n25390 );
not ( n25392 , n8367 );
not ( n25393 , n14591 );
or ( n25394 , n25392 , n25393 );
not ( n25395 , n8367 );
nand ( n25396 , n25395 , n14596 );
nand ( n25397 , n25394 , n25396 );
and ( n25398 , n25397 , n9302 );
not ( n25399 , n25397 );
and ( n25400 , n25399 , n9294 );
nor ( n25401 , n25398 , n25400 );
buf ( n25402 , n25401 );
not ( n25403 , n25402 );
not ( n25404 , n10301 );
not ( n25405 , n19947 );
xor ( n25406 , n25405 , n19957 );
xor ( n25407 , n25406 , n19964 );
not ( n25408 , n25407 );
not ( n25409 , n25408 );
or ( n25410 , n25404 , n25409 );
or ( n25411 , n25408 , n10301 );
nand ( n25412 , n25410 , n25411 );
buf ( n25413 , n12422 );
and ( n25414 , n25412 , n25413 );
not ( n25415 , n25412 );
not ( n25416 , n12417 );
not ( n25417 , n12405 );
not ( n25418 , n25417 );
or ( n25419 , n25416 , n25418 );
nand ( n25420 , n12405 , n12418 );
nand ( n25421 , n25419 , n25420 );
buf ( n25422 , n25421 );
and ( n25423 , n25415 , n25422 );
nor ( n25424 , n25414 , n25423 );
not ( n25425 , n25424 );
nand ( n25426 , n25403 , n25425 );
not ( n25427 , n25426 );
not ( n25428 , n9391 );
not ( n25429 , n16361 );
or ( n25430 , n25428 , n25429 );
not ( n25431 , n9391 );
nand ( n25432 , n25431 , n16356 );
nand ( n25433 , n25430 , n25432 );
not ( n25434 , n25433 );
buf ( n25435 , n6547 );
buf ( n25436 , n6548 );
buf ( n25437 , n25436 );
not ( n25438 , n25437 );
buf ( n25439 , n6549 );
not ( n25440 , n25439 );
not ( n25441 , n25440 );
or ( n25442 , n25438 , n25441 );
not ( n25443 , n25436 );
buf ( n25444 , n25439 );
nand ( n25445 , n25443 , n25444 );
nand ( n25446 , n25442 , n25445 );
xor ( n25447 , n25435 , n25446 );
buf ( n25448 , n6550 );
buf ( n25449 , n6551 );
not ( n25450 , n25449 );
xor ( n25451 , n25448 , n25450 );
buf ( n25452 , n6552 );
nand ( n25453 , n7478 , n25452 );
xnor ( n25454 , n25451 , n25453 );
xnor ( n25455 , n25447 , n25454 );
not ( n25456 , n25455 );
not ( n25457 , n25456 );
and ( n25458 , n25434 , n25457 );
buf ( n25459 , n25455 );
not ( n25460 , n25459 );
and ( n25461 , n25460 , n25433 );
nor ( n25462 , n25458 , n25461 );
not ( n25463 , n25462 );
not ( n25464 , n25463 );
and ( n25465 , n25427 , n25464 );
and ( n25466 , n25426 , n25463 );
nor ( n25467 , n25465 , n25466 );
and ( n25468 , n25391 , n25467 );
not ( n25469 , n25391 );
not ( n25470 , n25467 );
and ( n25471 , n25469 , n25470 );
nor ( n25472 , n25468 , n25471 );
and ( n25473 , n25303 , n25472 );
not ( n25474 , n25303 );
not ( n25475 , n25472 );
and ( n25476 , n25474 , n25475 );
nor ( n25477 , n25473 , n25476 );
not ( n25478 , n25477 );
not ( n25479 , n25478 );
not ( n25480 , n25479 );
and ( n25481 , n25195 , n25480 );
and ( n25482 , n25194 , n25479 );
nor ( n25483 , n25481 , n25482 );
buf ( n25484 , n13744 );
nor ( n25485 , n25483 , n25484 );
not ( n25486 , n25485 );
and ( n25487 , n10550 , n12200 );
not ( n25488 , n10550 );
not ( n25489 , n12200 );
and ( n25490 , n25488 , n25489 );
nor ( n25491 , n25487 , n25490 );
buf ( n25492 , n6553 );
buf ( n25493 , n6554 );
buf ( n25494 , n25493 );
not ( n25495 , n25494 );
buf ( n25496 , n6555 );
not ( n25497 , n25496 );
not ( n25498 , n25497 );
or ( n25499 , n25495 , n25498 );
not ( n25500 , n25493 );
buf ( n25501 , n25496 );
nand ( n25502 , n25500 , n25501 );
nand ( n25503 , n25499 , n25502 );
xor ( n25504 , n25492 , n25503 );
buf ( n25505 , n6556 );
not ( n25506 , n25505 );
xor ( n25507 , n17415 , n25506 );
buf ( n25508 , n6557 );
nand ( n25509 , n8934 , n25508 );
xnor ( n25510 , n25507 , n25509 );
xnor ( n25511 , n25504 , n25510 );
not ( n25512 , n25511 );
not ( n25513 , n25512 );
and ( n25514 , n25491 , n25513 );
not ( n25515 , n25491 );
not ( n25516 , n25511 );
and ( n25517 , n25515 , n25516 );
nor ( n25518 , n25514 , n25517 );
not ( n25519 , n16098 );
not ( n25520 , n19372 );
and ( n25521 , n25519 , n25520 );
and ( n25522 , n9169 , n19372 );
nor ( n25523 , n25521 , n25522 );
and ( n25524 , n25523 , n16093 );
not ( n25525 , n25523 );
not ( n25526 , n16093 );
and ( n25527 , n25525 , n25526 );
nor ( n25528 , n25524 , n25527 );
nand ( n25529 , n25518 , n25528 );
not ( n25530 , n25529 );
not ( n25531 , n7023 );
not ( n25532 , n21214 );
or ( n25533 , n25531 , n25532 );
nand ( n25534 , n9467 , n7019 );
nand ( n25535 , n25533 , n25534 );
not ( n25536 , n25535 );
buf ( n25537 , n6558 );
nand ( n25538 , n7955 , n25537 );
buf ( n25539 , n6559 );
buf ( n25540 , n25539 );
and ( n25541 , n25538 , n25540 );
not ( n25542 , n25538 );
not ( n25543 , n25539 );
and ( n25544 , n25542 , n25543 );
nor ( n25545 , n25541 , n25544 );
not ( n25546 , n25545 );
buf ( n25547 , n6560 );
nand ( n25548 , n8519 , n25547 );
buf ( n25549 , n6561 );
not ( n25550 , n25549 );
and ( n25551 , n25548 , n25550 );
not ( n25552 , n25548 );
buf ( n25553 , n25549 );
and ( n25554 , n25552 , n25553 );
nor ( n25555 , n25551 , n25554 );
not ( n25556 , n25555 );
or ( n25557 , n25546 , n25556 );
or ( n25558 , n25545 , n25555 );
nand ( n25559 , n25557 , n25558 );
not ( n25560 , n19937 );
buf ( n25561 , n6562 );
not ( n25562 , n25561 );
not ( n25563 , n25562 );
or ( n25564 , n25560 , n25563 );
not ( n25565 , n19936 );
buf ( n25566 , n25561 );
nand ( n25567 , n25565 , n25566 );
nand ( n25568 , n25564 , n25567 );
buf ( n25569 , n6563 );
not ( n25570 , n25569 );
and ( n25571 , n25568 , n25570 );
not ( n25572 , n25568 );
buf ( n25573 , n25569 );
and ( n25574 , n25572 , n25573 );
nor ( n25575 , n25571 , n25574 );
xor ( n25576 , n25559 , n25575 );
buf ( n25577 , n25576 );
not ( n25578 , n25577 );
and ( n25579 , n25536 , n25578 );
and ( n25580 , n25535 , n25577 );
nor ( n25581 , n25579 , n25580 );
not ( n25582 , n25581 );
not ( n25583 , n25582 );
and ( n25584 , n25530 , n25583 );
and ( n25585 , n25529 , n25582 );
nor ( n25586 , n25584 , n25585 );
not ( n25587 , n25586 );
not ( n25588 , n25587 );
not ( n25589 , n17080 );
not ( n25590 , n13343 );
or ( n25591 , n25589 , n25590 );
not ( n25592 , n17080 );
nand ( n25593 , n25592 , n13342 );
nand ( n25594 , n25591 , n25593 );
and ( n25595 , n25594 , n24203 );
not ( n25596 , n25594 );
not ( n25597 , n21577 );
and ( n25598 , n25596 , n25597 );
nor ( n25599 , n25595 , n25598 );
not ( n25600 , n25599 );
not ( n25601 , n11644 );
not ( n25602 , n10331 );
or ( n25603 , n25601 , n25602 );
not ( n25604 , n11644 );
nand ( n25605 , n25604 , n10330 );
nand ( n25606 , n25603 , n25605 );
and ( n25607 , n25606 , n10377 );
not ( n25608 , n25606 );
and ( n25609 , n25608 , n14494 );
nor ( n25610 , n25607 , n25609 );
nand ( n25611 , n25600 , n25610 );
not ( n25612 , n25611 );
not ( n25613 , n8594 );
not ( n25614 , n18897 );
or ( n25615 , n25613 , n25614 );
not ( n25616 , n8594 );
xor ( n25617 , n18877 , n18896 );
buf ( n25618 , n18886 );
xnor ( n25619 , n25617 , n25618 );
nand ( n25620 , n25616 , n25619 );
nand ( n25621 , n25615 , n25620 );
and ( n25622 , n25621 , n18906 );
not ( n25623 , n25621 );
and ( n25624 , n25623 , n18903 );
nor ( n25625 , n25622 , n25624 );
not ( n25626 , n25625 );
and ( n25627 , n25612 , n25626 );
and ( n25628 , n25611 , n25625 );
nor ( n25629 , n25627 , n25628 );
not ( n25630 , n22095 );
not ( n25631 , n9002 );
not ( n25632 , n19109 );
or ( n25633 , n25631 , n25632 );
or ( n25634 , n19109 , n9002 );
nand ( n25635 , n25633 , n25634 );
not ( n25636 , n25635 );
or ( n25637 , n25630 , n25636 );
or ( n25638 , n25635 , n22095 );
nand ( n25639 , n25637 , n25638 );
buf ( n25640 , n25639 );
not ( n25641 , n25640 );
not ( n25642 , n14653 );
buf ( n25643 , n9896 );
not ( n25644 , n25643 );
not ( n25645 , n25644 );
or ( n25646 , n25642 , n25645 );
nand ( n25647 , n25643 , n14649 );
nand ( n25648 , n25646 , n25647 );
buf ( n25649 , n21809 );
not ( n25650 , n25649 );
and ( n25651 , n25648 , n25650 );
not ( n25652 , n25648 );
buf ( n25653 , n20862 );
not ( n25654 , n25653 );
and ( n25655 , n25652 , n25654 );
nor ( n25656 , n25651 , n25655 );
nand ( n25657 , n25641 , n25656 );
not ( n25658 , n25657 );
buf ( n25659 , n16342 );
not ( n25660 , n25659 );
xor ( n25661 , n11341 , n11360 );
not ( n25662 , n11350 );
xnor ( n25663 , n25661 , n25662 );
not ( n25664 , n25663 );
or ( n25665 , n25660 , n25664 );
or ( n25666 , n25663 , n25659 );
nand ( n25667 , n25665 , n25666 );
buf ( n25668 , n6564 );
buf ( n25669 , n25668 );
not ( n25670 , n25669 );
buf ( n25671 , n6565 );
not ( n25672 , n25671 );
not ( n25673 , n25672 );
or ( n25674 , n25670 , n25673 );
not ( n25675 , n25668 );
buf ( n25676 , n25671 );
nand ( n25677 , n25675 , n25676 );
nand ( n25678 , n25674 , n25677 );
buf ( n25679 , n6566 );
not ( n25680 , n25679 );
and ( n25681 , n25678 , n25680 );
not ( n25682 , n25678 );
buf ( n25683 , n25679 );
and ( n25684 , n25682 , n25683 );
nor ( n25685 , n25681 , n25684 );
buf ( n25686 , n6567 );
nand ( n25687 , n7616 , n25686 );
buf ( n25688 , n6568 );
buf ( n25689 , n25688 );
and ( n25690 , n25687 , n25689 );
not ( n25691 , n25687 );
not ( n25692 , n25688 );
and ( n25693 , n25691 , n25692 );
nor ( n25694 , n25690 , n25693 );
xor ( n25695 , n25685 , n25694 );
xnor ( n25696 , n25695 , n22815 );
not ( n25697 , n25696 );
not ( n25698 , n25697 );
and ( n25699 , n25667 , n25698 );
not ( n25700 , n25667 );
and ( n25701 , n25700 , n25697 );
nor ( n25702 , n25699 , n25701 );
not ( n25703 , n25702 );
not ( n25704 , n25703 );
and ( n25705 , n25658 , n25704 );
and ( n25706 , n25657 , n25703 );
nor ( n25707 , n25705 , n25706 );
not ( n25708 , n25707 );
not ( n25709 , n15153 );
not ( n25710 , n17246 );
or ( n25711 , n25709 , n25710 );
not ( n25712 , n15153 );
nand ( n25713 , n25712 , n16719 );
nand ( n25714 , n25711 , n25713 );
and ( n25715 , n25714 , n20703 );
not ( n25716 , n25714 );
not ( n25717 , n20698 );
and ( n25718 , n25716 , n25717 );
nor ( n25719 , n25715 , n25718 );
not ( n25720 , n25719 );
not ( n25721 , n14673 );
not ( n25722 , n25254 );
not ( n25723 , n25722 );
or ( n25724 , n25721 , n25723 );
or ( n25725 , n25722 , n14673 );
nand ( n25726 , n25724 , n25725 );
and ( n25727 , n25726 , n13232 );
not ( n25728 , n25726 );
not ( n25729 , n13229 );
not ( n25730 , n25729 );
and ( n25731 , n25728 , n25730 );
nor ( n25732 , n25727 , n25731 );
nand ( n25733 , n25720 , n25732 );
not ( n25734 , n25733 );
xor ( n25735 , n24389 , n16782 );
xnor ( n25736 , n25735 , n19532 );
not ( n25737 , n25736 );
not ( n25738 , n25737 );
and ( n25739 , n25734 , n25738 );
and ( n25740 , n25733 , n25737 );
nor ( n25741 , n25739 , n25740 );
not ( n25742 , n25741 );
not ( n25743 , n25742 );
or ( n25744 , n25708 , n25743 );
not ( n25745 , n25707 );
nand ( n25746 , n25745 , n25741 );
nand ( n25747 , n25744 , n25746 );
xor ( n25748 , n25629 , n25747 );
not ( n25749 , n25518 );
nand ( n25750 , n25581 , n25749 );
buf ( n25751 , n10406 );
not ( n25752 , n25751 );
not ( n25753 , n22183 );
or ( n25754 , n25752 , n25753 );
or ( n25755 , n22975 , n25751 );
nand ( n25756 , n25754 , n25755 );
and ( n25757 , n25756 , n22980 );
not ( n25758 , n25756 );
and ( n25759 , n25758 , n22984 );
nor ( n25760 , n25757 , n25759 );
not ( n25761 , n25760 );
and ( n25762 , n25750 , n25761 );
not ( n25763 , n25750 );
and ( n25764 , n25763 , n25760 );
nor ( n25765 , n25762 , n25764 );
not ( n25766 , n25765 );
not ( n25767 , n25766 );
not ( n25768 , n7165 );
not ( n25769 , n19805 );
or ( n25770 , n25768 , n25769 );
not ( n25771 , n7165 );
nand ( n25772 , n25771 , n25051 );
nand ( n25773 , n25770 , n25772 );
not ( n25774 , n25063 );
and ( n25775 , n25773 , n25774 );
not ( n25776 , n25773 );
not ( n25777 , n25059 );
not ( n25778 , n25777 );
and ( n25779 , n25776 , n25778 );
nor ( n25780 , n25775 , n25779 );
not ( n25781 , n8301 );
not ( n25782 , n11992 );
not ( n25783 , n25782 );
or ( n25784 , n25781 , n25783 );
or ( n25785 , n25782 , n8301 );
nand ( n25786 , n25784 , n25785 );
and ( n25787 , n25786 , n16488 );
not ( n25788 , n25786 );
buf ( n25789 , n16491 );
and ( n25790 , n25788 , n25789 );
nor ( n25791 , n25787 , n25790 );
buf ( n25792 , n25791 );
nand ( n25793 , n25780 , n25792 );
not ( n25794 , n25793 );
buf ( n25795 , n20630 );
and ( n25796 , n25795 , n23488 );
not ( n25797 , n25795 );
and ( n25798 , n25797 , n23482 );
nor ( n25799 , n25796 , n25798 );
not ( n25800 , n25799 );
not ( n25801 , n24709 );
or ( n25802 , n25800 , n25801 );
not ( n25803 , n24709 );
not ( n25804 , n25803 );
or ( n25805 , n25804 , n25799 );
nand ( n25806 , n25802 , n25805 );
buf ( n25807 , n25806 );
not ( n25808 , n25807 );
and ( n25809 , n25794 , n25808 );
and ( n25810 , n25793 , n25807 );
nor ( n25811 , n25809 , n25810 );
not ( n25812 , n25811 );
not ( n25813 , n25812 );
or ( n25814 , n25767 , n25813 );
nand ( n25815 , n25811 , n25765 );
nand ( n25816 , n25814 , n25815 );
xor ( n25817 , n25748 , n25816 );
not ( n25818 , n25817 );
or ( n25819 , n25588 , n25818 );
not ( n25820 , n25587 );
not ( n25821 , n25747 );
not ( n25822 , n25821 );
not ( n25823 , n25629 );
and ( n25824 , n25816 , n25823 );
not ( n25825 , n25816 );
and ( n25826 , n25825 , n25629 );
nor ( n25827 , n25824 , n25826 );
not ( n25828 , n25827 );
or ( n25829 , n25822 , n25828 );
not ( n25830 , n25827 );
nand ( n25831 , n25830 , n25747 );
nand ( n25832 , n25829 , n25831 );
nand ( n25833 , n25820 , n25832 );
nand ( n25834 , n25819 , n25833 );
buf ( n25835 , n17263 );
and ( n25836 , n25834 , n25835 );
not ( n25837 , n25834 );
not ( n25838 , n17272 );
not ( n25839 , n25838 );
and ( n25840 , n25837 , n25839 );
nor ( n25841 , n25836 , n25840 );
not ( n25842 , n10586 );
not ( n25843 , n12204 );
not ( n25844 , n25843 );
or ( n25845 , n25842 , n25844 );
not ( n25846 , n10586 );
nand ( n25847 , n25846 , n12204 );
nand ( n25848 , n25845 , n25847 );
and ( n25849 , n25848 , n25516 );
not ( n25850 , n25848 );
and ( n25851 , n25850 , n25513 );
nor ( n25852 , n25849 , n25851 );
not ( n25853 , n25852 );
not ( n25854 , n8917 );
not ( n25855 , n18549 );
or ( n25856 , n25854 , n25855 );
or ( n25857 , n18549 , n8917 );
nand ( n25858 , n25856 , n25857 );
not ( n25859 , n20632 );
and ( n25860 , n25858 , n25859 );
not ( n25861 , n25858 );
and ( n25862 , n25861 , n20632 );
nor ( n25863 , n25860 , n25862 );
nand ( n25864 , n25853 , n25863 );
not ( n25865 , n25864 );
not ( n25866 , n15507 );
not ( n25867 , n9912 );
and ( n25868 , n25866 , n25867 );
and ( n25869 , n15507 , n9912 );
nor ( n25870 , n25868 , n25869 );
not ( n25871 , n15548 );
and ( n25872 , n25870 , n25871 );
not ( n25873 , n25870 );
and ( n25874 , n25873 , n15549 );
nor ( n25875 , n25872 , n25874 );
not ( n25876 , n25875 );
and ( n25877 , n25865 , n25876 );
not ( n25878 , n25875 );
not ( n25879 , n25878 );
and ( n25880 , n25864 , n25879 );
nor ( n25881 , n25877 , n25880 );
not ( n25882 , n25881 );
not ( n25883 , n25882 );
not ( n25884 , n19887 );
not ( n25885 , n25884 );
not ( n25886 , n13915 );
not ( n25887 , n24514 );
or ( n25888 , n25886 , n25887 );
or ( n25889 , n24514 , n13915 );
nand ( n25890 , n25888 , n25889 );
not ( n25891 , n25890 );
and ( n25892 , n25885 , n25891 );
and ( n25893 , n25884 , n25890 );
nor ( n25894 , n25892 , n25893 );
not ( n25895 , n25894 );
not ( n25896 , n25895 );
not ( n25897 , n22257 );
not ( n25898 , n9132 );
not ( n25899 , n17978 );
or ( n25900 , n25898 , n25899 );
or ( n25901 , n17978 , n9132 );
nand ( n25902 , n25900 , n25901 );
not ( n25903 , n25902 );
and ( n25904 , n25897 , n25903 );
and ( n25905 , n22257 , n25902 );
nor ( n25906 , n25904 , n25905 );
not ( n25907 , n25696 );
not ( n25908 , n25435 );
and ( n25909 , n25907 , n25908 );
and ( n25910 , n25696 , n25435 );
nor ( n25911 , n25909 , n25910 );
buf ( n25912 , n20330 );
xor ( n25913 , n25911 , n25912 );
nand ( n25914 , n25906 , n25913 );
not ( n25915 , n25914 );
or ( n25916 , n25896 , n25915 );
or ( n25917 , n25914 , n25895 );
nand ( n25918 , n25916 , n25917 );
not ( n25919 , n25918 );
not ( n25920 , n25875 );
not ( n25921 , n25863 );
nand ( n25922 , n25920 , n25921 );
not ( n25923 , n25922 );
not ( n25924 , n24845 );
not ( n25925 , n23790 );
or ( n25926 , n25924 , n25925 );
or ( n25927 , n23790 , n24845 );
nand ( n25928 , n25926 , n25927 );
not ( n25929 , n15119 );
and ( n25930 , n25928 , n25929 );
not ( n25931 , n25928 );
and ( n25932 , n25931 , n15120 );
nor ( n25933 , n25930 , n25932 );
not ( n25934 , n25933 );
not ( n25935 , n25934 );
and ( n25936 , n25923 , n25935 );
nand ( n25937 , n25878 , n25921 );
and ( n25938 , n25937 , n25934 );
nor ( n25939 , n25936 , n25938 );
not ( n25940 , n25939 );
and ( n25941 , n25919 , n25940 );
and ( n25942 , n25918 , n25939 );
nor ( n25943 , n25941 , n25942 );
not ( n25944 , n25943 );
xor ( n25945 , n15659 , n21026 );
xnor ( n25946 , n25945 , n25313 );
not ( n25947 , n8681 );
not ( n25948 , n15886 );
not ( n25949 , n15896 );
or ( n25950 , n25948 , n25949 );
or ( n25951 , n15886 , n15896 );
nand ( n25952 , n25950 , n25951 );
xnor ( n25953 , n25952 , n15877 );
not ( n25954 , n25953 );
or ( n25955 , n25947 , n25954 );
not ( n25956 , n8680 );
nand ( n25957 , n15898 , n25956 );
nand ( n25958 , n25955 , n25957 );
and ( n25959 , n25958 , n15938 );
not ( n25960 , n25958 );
and ( n25961 , n25960 , n15937 );
nor ( n25962 , n25959 , n25961 );
nand ( n25963 , n25946 , n25962 );
not ( n25964 , n12005 );
not ( n25965 , n22633 );
or ( n25966 , n25964 , n25965 );
or ( n25967 , n12005 , n18458 );
nand ( n25968 , n25966 , n25967 );
and ( n25969 , n25968 , n18491 );
not ( n25970 , n25968 );
and ( n25971 , n25970 , n18497 );
nor ( n25972 , n25969 , n25971 );
not ( n25973 , n25972 );
and ( n25974 , n25963 , n25973 );
not ( n25975 , n25963 );
and ( n25976 , n25975 , n25972 );
nor ( n25977 , n25974 , n25976 );
not ( n25978 , n25977 );
and ( n25979 , n25944 , n25978 );
and ( n25980 , n25943 , n25977 );
nor ( n25981 , n25979 , n25980 );
not ( n25982 , n25981 );
not ( n25983 , n25982 );
not ( n25984 , n13366 );
not ( n25985 , n22651 );
or ( n25986 , n25984 , n25985 );
buf ( n25987 , n15647 );
nand ( n25988 , n25987 , n13363 );
nand ( n25989 , n25986 , n25988 );
not ( n25990 , n15599 );
not ( n25991 , n25990 );
not ( n25992 , n15583 );
and ( n25993 , n25991 , n25992 );
and ( n25994 , n25990 , n15583 );
nor ( n25995 , n25993 , n25994 );
buf ( n25996 , n25995 );
and ( n25997 , n25989 , n25996 );
not ( n25998 , n25989 );
and ( n25999 , n25998 , n15604 );
nor ( n26000 , n25997 , n25999 );
not ( n26001 , n26000 );
not ( n26002 , n7679 );
not ( n26003 , n17837 );
not ( n26004 , n26003 );
not ( n26005 , n26004 );
or ( n26006 , n26002 , n26005 );
not ( n26007 , n26003 );
or ( n26008 , n26007 , n7679 );
nand ( n26009 , n26006 , n26008 );
and ( n26010 , n26009 , n17239 );
not ( n26011 , n26009 );
not ( n26012 , n17239 );
and ( n26013 , n26011 , n26012 );
nor ( n26014 , n26010 , n26013 );
nand ( n26015 , n26001 , n26014 );
not ( n26016 , n26015 );
not ( n26017 , n7994 );
not ( n26018 , n17112 );
or ( n26019 , n26017 , n26018 );
or ( n26020 , n17112 , n7994 );
nand ( n26021 , n26019 , n26020 );
not ( n26022 , n26021 );
not ( n26023 , n17126 );
or ( n26024 , n26022 , n26023 );
or ( n26025 , n22339 , n26021 );
nand ( n26026 , n26024 , n26025 );
not ( n26027 , n26026 );
not ( n26028 , n26027 );
not ( n26029 , n26028 );
and ( n26030 , n26016 , n26029 );
and ( n26031 , n26015 , n26028 );
nor ( n26032 , n26030 , n26031 );
not ( n26033 , n26032 );
xor ( n26034 , n10218 , n9780 );
xnor ( n26035 , n26034 , n15843 );
not ( n26036 , n26035 );
xor ( n26037 , n9995 , n7584 );
not ( n26038 , n17873 );
xnor ( n26039 , n26037 , n26038 );
nand ( n26040 , n26036 , n26039 );
and ( n26041 , n10865 , n6638 );
not ( n26042 , n10865 );
and ( n26043 , n26042 , n6634 );
or ( n26044 , n26041 , n26043 );
not ( n26045 , n26044 );
not ( n26046 , n13857 );
or ( n26047 , n26045 , n26046 );
or ( n26048 , n13857 , n26044 );
nand ( n26049 , n26047 , n26048 );
buf ( n26050 , n26049 );
not ( n26051 , n26050 );
and ( n26052 , n26040 , n26051 );
not ( n26053 , n26040 );
and ( n26054 , n26053 , n26050 );
nor ( n26055 , n26052 , n26054 );
not ( n26056 , n26055 );
or ( n26057 , n26033 , n26056 );
or ( n26058 , n26055 , n26032 );
nand ( n26059 , n26057 , n26058 );
not ( n26060 , n26059 );
not ( n26061 , n26060 );
and ( n26062 , n25983 , n26061 );
not ( n26063 , n25981 );
and ( n26064 , n26063 , n26060 );
nor ( n26065 , n26062 , n26064 );
not ( n26066 , n26065 );
or ( n26067 , n25883 , n26066 );
not ( n26068 , n25882 );
not ( n26069 , n26059 );
not ( n26070 , n25981 );
or ( n26071 , n26069 , n26070 );
nand ( n26072 , n25982 , n26060 );
nand ( n26073 , n26071 , n26072 );
nand ( n26074 , n26068 , n26073 );
nand ( n26075 , n26067 , n26074 );
not ( n26076 , n15554 );
not ( n26077 , n16218 );
nand ( n26078 , n26076 , n26077 );
not ( n26079 , n26078 );
not ( n26080 , n21809 );
not ( n26081 , n14644 );
not ( n26082 , n9896 );
not ( n26083 , n26082 );
or ( n26084 , n26081 , n26083 );
not ( n26085 , n9896 );
or ( n26086 , n26085 , n14644 );
nand ( n26087 , n26084 , n26086 );
not ( n26088 , n26087 );
or ( n26089 , n26080 , n26088 );
or ( n26090 , n26087 , n25654 );
nand ( n26091 , n26089 , n26090 );
not ( n26092 , n26091 );
and ( n26093 , n26079 , n26092 );
not ( n26094 , n26091 );
not ( n26095 , n26094 );
and ( n26096 , n26078 , n26095 );
nor ( n26097 , n26093 , n26096 );
not ( n26098 , n26097 );
buf ( n26099 , n23460 );
not ( n26100 , n26099 );
not ( n26101 , n18335 );
or ( n26102 , n26100 , n26101 );
or ( n26103 , n18338 , n26099 );
nand ( n26104 , n26102 , n26103 );
and ( n26105 , n26104 , n18370 );
not ( n26106 , n26104 );
and ( n26107 , n26106 , n18373 );
nor ( n26108 , n26105 , n26107 );
not ( n26109 , n26108 );
not ( n26110 , n26109 );
not ( n26111 , n16052 );
nand ( n26112 , n26111 , n16106 );
not ( n26113 , n26112 );
or ( n26114 , n26110 , n26113 );
or ( n26115 , n26112 , n26109 );
nand ( n26116 , n26114 , n26115 );
not ( n26117 , n26116 );
not ( n26118 , n26117 );
not ( n26119 , n15657 );
nand ( n26120 , n26119 , n15570 );
not ( n26121 , n21515 );
not ( n26122 , n24875 );
and ( n26123 , n8118 , n26122 );
not ( n26124 , n8118 );
and ( n26125 , n26124 , n24875 );
nor ( n26126 , n26123 , n26125 );
not ( n26127 , n26126 );
and ( n26128 , n26121 , n26127 );
not ( n26129 , n26121 );
and ( n26130 , n26129 , n26126 );
nor ( n26131 , n26128 , n26130 );
not ( n26132 , n26131 );
and ( n26133 , n26120 , n26132 );
not ( n26134 , n26120 );
and ( n26135 , n26134 , n26131 );
nor ( n26136 , n26133 , n26135 );
not ( n26137 , n26136 );
not ( n26138 , n26137 );
or ( n26139 , n26118 , n26138 );
nand ( n26140 , n26136 , n26116 );
nand ( n26141 , n26139 , n26140 );
not ( n26142 , n26141 );
or ( n26143 , n26098 , n26142 );
or ( n26144 , n26141 , n26097 );
nand ( n26145 , n26143 , n26144 );
not ( n26146 , n15845 );
not ( n26147 , n15940 );
nand ( n26148 , n26146 , n26147 );
not ( n26149 , n26148 );
xor ( n26150 , n6747 , n11756 );
xnor ( n26151 , n26150 , n14061 );
not ( n26152 , n26151 );
or ( n26153 , n26149 , n26152 );
or ( n26154 , n26151 , n26148 );
nand ( n26155 , n26153 , n26154 );
not ( n26156 , n26155 );
nand ( n26157 , n15992 , n16023 );
not ( n26158 , n26157 );
not ( n26159 , n17641 );
not ( n26160 , n24003 );
or ( n26161 , n26159 , n26160 );
or ( n26162 , n24003 , n17641 );
nand ( n26163 , n26161 , n26162 );
and ( n26164 , n26163 , n20809 );
not ( n26165 , n26163 );
not ( n26166 , n20755 );
and ( n26167 , n26165 , n26166 );
or ( n26168 , n26164 , n26167 );
not ( n26169 , n26168 );
not ( n26170 , n26169 );
and ( n26171 , n26158 , n26170 );
and ( n26172 , n26157 , n26169 );
nor ( n26173 , n26171 , n26172 );
not ( n26174 , n26173 );
or ( n26175 , n26156 , n26174 );
or ( n26176 , n26173 , n26155 );
nand ( n26177 , n26175 , n26176 );
not ( n26178 , n26177 );
and ( n26179 , n26145 , n26178 );
not ( n26180 , n26145 );
and ( n26181 , n26180 , n26177 );
nor ( n26182 , n26179 , n26181 );
buf ( n26183 , n26182 );
not ( n26184 , n26183 );
and ( n26185 , n26075 , n26184 );
not ( n26186 , n26075 );
and ( n26187 , n26186 , n26183 );
nor ( n26188 , n26185 , n26187 );
not ( n26189 , n26188 );
nand ( n26190 , n25841 , n26189 );
or ( n26191 , n25486 , n26190 );
not ( n26192 , n26189 );
not ( n26193 , n25483 );
not ( n26194 , n26193 );
or ( n26195 , n26192 , n26194 );
buf ( n26196 , n22058 );
nor ( n26197 , n25841 , n26196 );
nand ( n26198 , n26195 , n26197 );
nand ( n26199 , n13766 , n9753 );
nand ( n26200 , n26191 , n26198 , n26199 );
buf ( n26201 , n26200 );
buf ( n26202 , n26201 );
buf ( n26203 , n11775 );
not ( n26204 , n26203 );
not ( n26205 , n11772 );
and ( n26206 , n26204 , n26205 );
and ( n26207 , n26203 , n11772 );
nor ( n26208 , n26206 , n26207 );
not ( n26209 , n26208 );
buf ( n26210 , n8488 );
not ( n26211 , n26210 );
or ( n26212 , n26209 , n26211 );
or ( n26213 , n26210 , n26208 );
nand ( n26214 , n26212 , n26213 );
and ( n26215 , n26214 , n8532 );
not ( n26216 , n26214 );
not ( n26217 , n8532 );
and ( n26218 , n26216 , n26217 );
nor ( n26219 , n26215 , n26218 );
not ( n26220 , n26219 );
xor ( n26221 , n13004 , n23694 );
xnor ( n26222 , n26221 , n16442 );
nand ( n26223 , n26220 , n26222 );
not ( n26224 , n26223 );
not ( n26225 , n9489 );
not ( n26226 , n6845 );
not ( n26227 , n16533 );
or ( n26228 , n26226 , n26227 );
or ( n26229 , n16538 , n6845 );
nand ( n26230 , n26228 , n26229 );
not ( n26231 , n26230 );
or ( n26232 , n26225 , n26231 );
or ( n26233 , n26230 , n9489 );
nand ( n26234 , n26232 , n26233 );
not ( n26235 , n26234 );
not ( n26236 , n26235 );
not ( n26237 , n26236 );
and ( n26238 , n26224 , n26237 );
and ( n26239 , n26223 , n26236 );
nor ( n26240 , n26238 , n26239 );
not ( n26241 , n26240 );
not ( n26242 , n14429 );
not ( n26243 , n18031 );
and ( n26244 , n26242 , n26243 );
and ( n26245 , n14429 , n18031 );
nor ( n26246 , n26244 , n26245 );
and ( n26247 , n26246 , n20518 );
not ( n26248 , n26246 );
and ( n26249 , n26248 , n21227 );
nor ( n26250 , n26247 , n26249 );
buf ( n26251 , n26250 );
not ( n26252 , n26251 );
xor ( n26253 , n10349 , n25421 );
xnor ( n26254 , n26253 , n12468 );
buf ( n26255 , n7614 );
not ( n26256 , n26255 );
not ( n26257 , n10941 );
or ( n26258 , n26256 , n26257 );
or ( n26259 , n10941 , n26255 );
nand ( n26260 , n26258 , n26259 );
nor ( n26261 , n19390 , n26260 );
not ( n26262 , n26261 );
nand ( n26263 , n19391 , n26260 );
nand ( n26264 , n26262 , n26263 );
nand ( n26265 , n26254 , n26264 );
not ( n26266 , n26265 );
or ( n26267 , n26252 , n26266 );
or ( n26268 , n26265 , n26251 );
nand ( n26269 , n26267 , n26268 );
not ( n26270 , n26269 );
buf ( n26271 , n20267 );
not ( n26272 , n26271 );
not ( n26273 , n22214 );
or ( n26274 , n26272 , n26273 );
or ( n26275 , n22214 , n26271 );
nand ( n26276 , n26274 , n26275 );
and ( n26277 , n26276 , n23302 );
not ( n26278 , n26276 );
and ( n26279 , n26278 , n23303 );
nor ( n26280 , n26277 , n26279 );
not ( n26281 , n12958 );
not ( n26282 , n16901 );
or ( n26283 , n26281 , n26282 );
or ( n26284 , n16901 , n12958 );
nand ( n26285 , n26283 , n26284 );
and ( n26286 , n26285 , n14537 );
not ( n26287 , n26285 );
and ( n26288 , n26287 , n22535 );
nor ( n26289 , n26286 , n26288 );
nand ( n26290 , n26280 , n26289 );
not ( n26291 , n26290 );
not ( n26292 , n25459 );
nand ( n26293 , n16361 , n9356 );
not ( n26294 , n26293 );
nor ( n26295 , n16361 , n9356 );
nor ( n26296 , n26294 , n26295 );
not ( n26297 , n26296 );
or ( n26298 , n26292 , n26297 );
not ( n26299 , n25456 );
or ( n26300 , n26299 , n26296 );
nand ( n26301 , n26298 , n26300 );
not ( n26302 , n26301 );
and ( n26303 , n26291 , n26302 );
not ( n26304 , n26289 );
not ( n26305 , n26304 );
nand ( n26306 , n26305 , n26280 );
and ( n26307 , n26306 , n26301 );
nor ( n26308 , n26303 , n26307 );
not ( n26309 , n26308 );
or ( n26310 , n26270 , n26309 );
or ( n26311 , n26308 , n26269 );
nand ( n26312 , n26310 , n26311 );
buf ( n26313 , n20232 );
not ( n26314 , n26313 );
xor ( n26315 , n15367 , n26314 );
xnor ( n26316 , n26315 , n13500 );
not ( n26317 , n7488 );
not ( n26318 , n26317 );
not ( n26319 , n26318 );
not ( n26320 , n13812 );
not ( n26321 , n13617 );
not ( n26322 , n26321 );
or ( n26323 , n26320 , n26322 );
or ( n26324 , n17672 , n13812 );
nand ( n26325 , n26323 , n26324 );
not ( n26326 , n26325 );
or ( n26327 , n26319 , n26326 );
or ( n26328 , n26325 , n7489 );
nand ( n26329 , n26327 , n26328 );
not ( n26330 , n26329 );
nand ( n26331 , n26316 , n26330 );
not ( n26332 , n18780 );
not ( n26333 , n9038 );
not ( n26334 , n22089 );
or ( n26335 , n26333 , n26334 );
or ( n26336 , n22089 , n9038 );
nand ( n26337 , n26335 , n26336 );
not ( n26338 , n26337 );
and ( n26339 , n26332 , n26338 );
and ( n26340 , n18780 , n26337 );
nor ( n26341 , n26339 , n26340 );
and ( n26342 , n26331 , n26341 );
not ( n26343 , n26331 );
not ( n26344 , n26341 );
and ( n26345 , n26343 , n26344 );
nor ( n26346 , n26342 , n26345 );
not ( n26347 , n26346 );
and ( n26348 , n26312 , n26347 );
not ( n26349 , n26312 );
and ( n26350 , n26349 , n26346 );
nor ( n26351 , n26348 , n26350 );
not ( n26352 , n19026 );
not ( n26353 , n9306 );
and ( n26354 , n26352 , n26353 );
and ( n26355 , n19026 , n9306 );
nor ( n26356 , n26354 , n26355 );
and ( n26357 , n26356 , n15843 );
not ( n26358 , n26356 );
and ( n26359 , n26358 , n15842 );
nor ( n26360 , n26357 , n26359 );
not ( n26361 , n26360 );
nand ( n26362 , n26219 , n26235 );
not ( n26363 , n26362 );
or ( n26364 , n26361 , n26363 );
or ( n26365 , n26362 , n26360 );
nand ( n26366 , n26364 , n26365 );
not ( n26367 , n26366 );
not ( n26368 , n21686 );
not ( n26369 , n11822 );
or ( n26370 , n26368 , n26369 );
or ( n26371 , n13403 , n21686 );
nand ( n26372 , n26370 , n26371 );
xnor ( n26373 , n26372 , n11868 );
not ( n26374 , n17087 );
not ( n26375 , n13343 );
or ( n26376 , n26374 , n26375 );
not ( n26377 , n17087 );
nand ( n26378 , n26377 , n17698 );
nand ( n26379 , n26376 , n26378 );
not ( n26380 , n25597 );
and ( n26381 , n26379 , n26380 );
not ( n26382 , n26379 );
and ( n26383 , n26382 , n21572 );
nor ( n26384 , n26381 , n26383 );
not ( n26385 , n26384 );
nand ( n26386 , n26373 , n26385 );
not ( n26387 , n26386 );
buf ( n26388 , n9606 );
not ( n26389 , n26388 );
not ( n26390 , n13708 );
or ( n26391 , n26389 , n26390 );
or ( n26392 , n13708 , n26388 );
nand ( n26393 , n26391 , n26392 );
not ( n26394 , n26393 );
not ( n26395 , n22963 );
and ( n26396 , n26394 , n26395 );
and ( n26397 , n26393 , n22960 );
nor ( n26398 , n26396 , n26397 );
not ( n26399 , n26398 );
not ( n26400 , n26399 );
and ( n26401 , n26387 , n26400 );
and ( n26402 , n26386 , n26399 );
nor ( n26403 , n26401 , n26402 );
not ( n26404 , n26403 );
or ( n26405 , n26367 , n26404 );
or ( n26406 , n26403 , n26366 );
nand ( n26407 , n26405 , n26406 );
not ( n26408 , n26407 );
and ( n26409 , n26351 , n26408 );
not ( n26410 , n26351 );
and ( n26411 , n26410 , n26407 );
nor ( n26412 , n26409 , n26411 );
buf ( n26413 , n26412 );
not ( n26414 , n26413 );
or ( n26415 , n26241 , n26414 );
or ( n26416 , n26413 , n26240 );
nand ( n26417 , n26415 , n26416 );
not ( n26418 , n10667 );
not ( n26419 , n20430 );
or ( n26420 , n26418 , n26419 );
nand ( n26421 , n20436 , n10663 );
nand ( n26422 , n26420 , n26421 );
not ( n26423 , n26422 );
not ( n26424 , n22232 );
and ( n26425 , n26423 , n26424 );
not ( n26426 , n19452 );
and ( n26427 , n26422 , n26426 );
nor ( n26428 , n26425 , n26427 );
not ( n26429 , n26428 );
not ( n26430 , n18066 );
not ( n26431 , n14429 );
or ( n26432 , n26430 , n26431 );
not ( n26433 , n18066 );
not ( n26434 , n14429 );
nand ( n26435 , n26433 , n26434 );
nand ( n26436 , n26432 , n26435 );
and ( n26437 , n26436 , n20518 );
not ( n26438 , n26436 );
and ( n26439 , n26438 , n21227 );
nor ( n26440 , n26437 , n26439 );
nand ( n26441 , n26429 , n26440 );
not ( n26442 , n26441 );
not ( n26443 , n11810 );
not ( n26444 , n25995 );
or ( n26445 , n26443 , n26444 );
not ( n26446 , n11810 );
nand ( n26447 , n26446 , n15603 );
nand ( n26448 , n26445 , n26447 );
buf ( n26449 , n13837 );
and ( n26450 , n26448 , n26449 );
not ( n26451 , n26448 );
not ( n26452 , n26449 );
and ( n26453 , n26451 , n26452 );
nor ( n26454 , n26450 , n26453 );
not ( n26455 , n26454 );
and ( n26456 , n26442 , n26455 );
nand ( n26457 , n26429 , n26440 );
and ( n26458 , n26457 , n26454 );
nor ( n26459 , n26456 , n26458 );
not ( n26460 , n26459 );
not ( n26461 , n26460 );
not ( n26462 , n9489 );
buf ( n26463 , n6860 );
not ( n26464 , n26463 );
not ( n26465 , n16537 );
or ( n26466 , n26464 , n26465 );
or ( n26467 , n16537 , n26463 );
nand ( n26468 , n26466 , n26467 );
not ( n26469 , n26468 );
and ( n26470 , n26462 , n26469 );
and ( n26471 , n9489 , n26468 );
nor ( n26472 , n26470 , n26471 );
not ( n26473 , n19222 );
not ( n26474 , n9031 );
or ( n26475 , n26473 , n26474 );
not ( n26476 , n19222 );
not ( n26477 , n9031 );
nand ( n26478 , n26476 , n26477 );
nand ( n26479 , n26475 , n26478 );
and ( n26480 , n26479 , n9075 );
not ( n26481 , n26479 );
and ( n26482 , n26481 , n9076 );
nor ( n26483 , n26480 , n26482 );
nand ( n26484 , n26472 , n26483 );
not ( n26485 , n26484 );
xor ( n26486 , n24967 , n13396 );
xnor ( n26487 , n26486 , n23201 );
not ( n26488 , n26487 );
or ( n26489 , n26485 , n26488 );
or ( n26490 , n26487 , n26484 );
nand ( n26491 , n26489 , n26490 );
not ( n26492 , n26491 );
not ( n26493 , n26492 );
or ( n26494 , n26461 , n26493 );
nand ( n26495 , n26491 , n26459 );
nand ( n26496 , n26494 , n26495 );
not ( n26497 , n20932 );
not ( n26498 , n9393 );
not ( n26499 , n26498 );
or ( n26500 , n26497 , n26499 );
not ( n26501 , n20932 );
nand ( n26502 , n26501 , n9393 );
nand ( n26503 , n26500 , n26502 );
and ( n26504 , n26503 , n9405 );
not ( n26505 , n26503 );
and ( n26506 , n26505 , n7672 );
nor ( n26507 , n26504 , n26506 );
not ( n26508 , n26507 );
not ( n26509 , n23342 );
not ( n26510 , n7520 );
or ( n26511 , n26509 , n26510 );
not ( n26512 , n23342 );
buf ( n26513 , n7499 );
xor ( n26514 , n26513 , n7509 );
xnor ( n26515 , n26514 , n7519 );
nand ( n26516 , n26512 , n26515 );
nand ( n26517 , n26511 , n26516 );
and ( n26518 , n26517 , n18550 );
not ( n26519 , n26517 );
not ( n26520 , n18550 );
and ( n26521 , n26519 , n26520 );
nor ( n26522 , n26518 , n26521 );
not ( n26523 , n26522 );
nand ( n26524 , n26508 , n26523 );
not ( n26525 , n26524 );
not ( n26526 , n18403 );
buf ( n26527 , n9157 );
not ( n26528 , n26527 );
not ( n26529 , n17979 );
or ( n26530 , n26528 , n26529 );
or ( n26531 , n17979 , n26527 );
nand ( n26532 , n26530 , n26531 );
and ( n26533 , n26526 , n26532 );
not ( n26534 , n26526 );
not ( n26535 , n26532 );
and ( n26536 , n26534 , n26535 );
nor ( n26537 , n26533 , n26536 );
not ( n26538 , n26537 );
and ( n26539 , n26525 , n26538 );
and ( n26540 , n26524 , n26537 );
nor ( n26541 , n26539 , n26540 );
not ( n26542 , n26541 );
and ( n26543 , n26496 , n26542 );
not ( n26544 , n26496 );
and ( n26545 , n26544 , n26541 );
nor ( n26546 , n26543 , n26545 );
buf ( n26547 , n26546 );
not ( n26548 , n25511 );
not ( n26549 , n13027 );
and ( n26550 , n26548 , n26549 );
and ( n26551 , n25513 , n13027 );
nor ( n26552 , n26550 , n26551 );
and ( n26553 , n23108 , n23126 );
not ( n26554 , n23108 );
and ( n26555 , n26554 , n23127 );
nor ( n26556 , n26553 , n26555 );
buf ( n26557 , n26556 );
and ( n26558 , n26552 , n26557 );
not ( n26559 , n26552 );
not ( n26560 , n26557 );
and ( n26561 , n26559 , n26560 );
nor ( n26562 , n26558 , n26561 );
not ( n26563 , n26562 );
not ( n26564 , n8114 );
not ( n26565 , n24876 );
or ( n26566 , n26564 , n26565 );
buf ( n26567 , n24875 );
nand ( n26568 , n26567 , n8110 );
nand ( n26569 , n26566 , n26568 );
and ( n26570 , n26569 , n26121 );
not ( n26571 , n26569 );
not ( n26572 , n21514 );
not ( n26573 , n26572 );
and ( n26574 , n26571 , n26573 );
nor ( n26575 , n26570 , n26574 );
not ( n26576 , n26575 );
nand ( n26577 , n26563 , n26576 );
not ( n26578 , n26577 );
not ( n26579 , n13564 );
and ( n26580 , n13568 , n26579 );
not ( n26581 , n13568 );
and ( n26582 , n26581 , n13565 );
nor ( n26583 , n26580 , n26582 );
not ( n26584 , n26583 );
not ( n26585 , n7628 );
or ( n26586 , n26584 , n26585 );
not ( n26587 , n7628 );
not ( n26588 , n26583 );
nand ( n26589 , n26587 , n26588 );
nand ( n26590 , n26586 , n26589 );
buf ( n26591 , n6569 );
buf ( n26592 , n26591 );
not ( n26593 , n26592 );
buf ( n26594 , n6570 );
not ( n26595 , n26594 );
not ( n26596 , n26595 );
or ( n26597 , n26593 , n26596 );
not ( n26598 , n26591 );
buf ( n26599 , n26594 );
nand ( n26600 , n26598 , n26599 );
nand ( n26601 , n26597 , n26600 );
buf ( n26602 , n6571 );
buf ( n26603 , n26602 );
and ( n26604 , n26601 , n26603 );
not ( n26605 , n26601 );
not ( n26606 , n26602 );
and ( n26607 , n26605 , n26606 );
nor ( n26608 , n26604 , n26607 );
buf ( n26609 , n6572 );
nand ( n26610 , n7133 , n26609 );
buf ( n26611 , n6573 );
not ( n26612 , n26611 );
and ( n26613 , n26610 , n26612 );
not ( n26614 , n26610 );
buf ( n26615 , n26611 );
and ( n26616 , n26614 , n26615 );
nor ( n26617 , n26613 , n26616 );
xor ( n26618 , n26608 , n26617 );
xnor ( n26619 , n26618 , n25215 );
buf ( n26620 , n26619 );
and ( n26621 , n26590 , n26620 );
not ( n26622 , n26590 );
not ( n26623 , n26620 );
and ( n26624 , n26622 , n26623 );
nor ( n26625 , n26621 , n26624 );
not ( n26626 , n26625 );
not ( n26627 , n26626 );
and ( n26628 , n26578 , n26627 );
and ( n26629 , n26577 , n26626 );
nor ( n26630 , n26628 , n26629 );
not ( n26631 , n26630 );
not ( n26632 , n6689 );
buf ( n26633 , n14101 );
not ( n26634 , n26633 );
or ( n26635 , n26632 , n26634 );
not ( n26636 , n20697 );
or ( n26637 , n26636 , n6689 );
nand ( n26638 , n26635 , n26637 );
and ( n26639 , n26638 , n14061 );
not ( n26640 , n26638 );
and ( n26641 , n26640 , n11778 );
nor ( n26642 , n26639 , n26641 );
not ( n26643 , n26642 );
not ( n26644 , n17882 );
not ( n26645 , n26644 );
not ( n26646 , n13666 );
or ( n26647 , n26645 , n26646 );
or ( n26648 , n13666 , n26644 );
nand ( n26649 , n26647 , n26648 );
and ( n26650 , n26649 , n13709 );
not ( n26651 , n26649 );
not ( n26652 , n13709 );
and ( n26653 , n26651 , n26652 );
nor ( n26654 , n26650 , n26653 );
nand ( n26655 , n26643 , n26654 );
buf ( n26656 , n13826 );
not ( n26657 , n26656 );
not ( n26658 , n13618 );
or ( n26659 , n26657 , n26658 );
not ( n26660 , n17672 );
or ( n26661 , n26660 , n26656 );
nand ( n26662 , n26659 , n26661 );
and ( n26663 , n26662 , n7495 );
not ( n26664 , n26662 );
and ( n26665 , n26664 , n13576 );
nor ( n26666 , n26663 , n26665 );
not ( n26667 , n26666 );
and ( n26668 , n26655 , n26667 );
not ( n26669 , n26655 );
and ( n26670 , n26669 , n26666 );
nor ( n26671 , n26668 , n26670 );
not ( n26672 , n26671 );
and ( n26673 , n26631 , n26672 );
and ( n26674 , n26630 , n26671 );
nor ( n26675 , n26673 , n26674 );
buf ( n26676 , n26675 );
xor ( n26677 , n26547 , n26676 );
buf ( n26678 , n26677 );
and ( n26679 , n26417 , n26678 );
not ( n26680 , n26417 );
not ( n26681 , n26675 );
not ( n26682 , n26546 );
or ( n26683 , n26681 , n26682 );
not ( n26684 , n26546 );
not ( n26685 , n26675 );
nand ( n26686 , n26684 , n26685 );
nand ( n26687 , n26683 , n26686 );
buf ( n26688 , n26687 );
and ( n26689 , n26680 , n26688 );
nor ( n26690 , n26679 , n26689 );
not ( n26691 , n19016 );
nand ( n26692 , n26690 , n26691 );
not ( n26693 , n20809 );
not ( n26694 , n20794 );
buf ( n26695 , n17655 );
not ( n26696 , n26695 );
and ( n26697 , n26694 , n26696 );
not ( n26698 , n24003 );
and ( n26699 , n26698 , n26695 );
nor ( n26700 , n26697 , n26699 );
not ( n26701 , n26700 );
and ( n26702 , n26693 , n26701 );
and ( n26703 , n24013 , n26700 );
nor ( n26704 , n26702 , n26703 );
nand ( n26705 , n26704 , n16814 );
not ( n26706 , n14382 );
not ( n26707 , n24685 );
or ( n26708 , n26706 , n26707 );
not ( n26709 , n14382 );
not ( n26710 , n24684 );
not ( n26711 , n26710 );
nand ( n26712 , n26709 , n26711 );
nand ( n26713 , n26708 , n26712 );
buf ( n26714 , n6574 );
buf ( n26715 , n26714 );
not ( n26716 , n26715 );
buf ( n26717 , n6575 );
not ( n26718 , n26717 );
not ( n26719 , n26718 );
or ( n26720 , n26716 , n26719 );
not ( n26721 , n26714 );
buf ( n26722 , n26717 );
nand ( n26723 , n26721 , n26722 );
nand ( n26724 , n26720 , n26723 );
and ( n26725 , n26724 , n10769 );
not ( n26726 , n26724 );
not ( n26727 , n10768 );
and ( n26728 , n26726 , n26727 );
nor ( n26729 , n26725 , n26728 );
buf ( n26730 , n6576 );
nand ( n26731 , n8344 , n26730 );
buf ( n26732 , n6577 );
buf ( n26733 , n26732 );
and ( n26734 , n26731 , n26733 );
not ( n26735 , n26731 );
not ( n26736 , n26732 );
and ( n26737 , n26735 , n26736 );
nor ( n26738 , n26734 , n26737 );
xor ( n26739 , n26729 , n26738 );
xor ( n26740 , n26739 , n23630 );
buf ( n26741 , n26740 );
not ( n26742 , n26741 );
and ( n26743 , n26713 , n26742 );
not ( n26744 , n26713 );
not ( n26745 , n26740 );
not ( n26746 , n26745 );
and ( n26747 , n26744 , n26746 );
nor ( n26748 , n26743 , n26747 );
and ( n26749 , n26705 , n26748 );
not ( n26750 , n26705 );
not ( n26751 , n26748 );
and ( n26752 , n26750 , n26751 );
nor ( n26753 , n26749 , n26752 );
not ( n26754 , n26753 );
not ( n26755 , n26754 );
not ( n26756 , n18395 );
not ( n26757 , n16997 );
or ( n26758 , n26756 , n26757 );
or ( n26759 , n16997 , n18395 );
nand ( n26760 , n26758 , n26759 );
xnor ( n26761 , n26760 , n17044 );
not ( n26762 , n26761 );
not ( n26763 , n11503 );
not ( n26764 , n18792 );
buf ( n26765 , n21917 );
not ( n26766 , n26765 );
and ( n26767 , n26764 , n26766 );
and ( n26768 , n13032 , n26765 );
nor ( n26769 , n26767 , n26768 );
xor ( n26770 , n26763 , n26769 );
nand ( n26771 , n26762 , n26770 );
not ( n26772 , n26771 );
not ( n26773 , n16551 );
and ( n26774 , n26772 , n26773 );
and ( n26775 , n26771 , n16551 );
nor ( n26776 , n26774 , n26775 );
not ( n26777 , n26776 );
buf ( n26778 , n15897 );
not ( n26779 , n26778 );
not ( n26780 , n10815 );
xor ( n26781 , n26780 , n10827 );
xnor ( n26782 , n26781 , n10843 );
not ( n26783 , n26782 );
or ( n26784 , n26779 , n26783 );
or ( n26785 , n26782 , n26778 );
nand ( n26786 , n26784 , n26785 );
and ( n26787 , n26786 , n22288 );
not ( n26788 , n26786 );
and ( n26789 , n26788 , n25034 );
nor ( n26790 , n26787 , n26789 );
not ( n26791 , n7297 );
not ( n26792 , n26791 );
not ( n26793 , n26792 );
not ( n26794 , n21056 );
or ( n26795 , n26793 , n26794 );
or ( n26796 , n21056 , n26792 );
nand ( n26797 , n26795 , n26796 );
and ( n26798 , n26797 , n21104 );
not ( n26799 , n26797 );
and ( n26800 , n26799 , n21098 );
nor ( n26801 , n26798 , n26800 );
not ( n26802 , n26801 );
nand ( n26803 , n26790 , n26802 );
not ( n26804 , n16724 );
and ( n26805 , n26803 , n26804 );
not ( n26806 , n26803 );
and ( n26807 , n26806 , n16724 );
nor ( n26808 , n26805 , n26807 );
not ( n26809 , n26808 );
or ( n26810 , n26777 , n26809 );
or ( n26811 , n26808 , n26776 );
nand ( n26812 , n26810 , n26811 );
not ( n26813 , n26704 );
nand ( n26814 , n26813 , n26751 );
not ( n26815 , n16798 );
and ( n26816 , n26814 , n26815 );
not ( n26817 , n26814 );
and ( n26818 , n26817 , n16798 );
nor ( n26819 , n26816 , n26818 );
and ( n26820 , n26812 , n26819 );
not ( n26821 , n26812 );
not ( n26822 , n26819 );
and ( n26823 , n26821 , n26822 );
nor ( n26824 , n26820 , n26823 );
not ( n26825 , n26824 );
buf ( n26826 , n19479 );
not ( n26827 , n26826 );
not ( n26828 , n14242 );
or ( n26829 , n26827 , n26828 );
or ( n26830 , n14242 , n26826 );
nand ( n26831 , n26829 , n26830 );
and ( n26832 , n26831 , n14293 );
not ( n26833 , n26831 );
and ( n26834 , n26833 , n14290 );
nor ( n26835 , n26832 , n26834 );
not ( n26836 , n26835 );
buf ( n26837 , n25509 );
buf ( n26838 , n25505 );
and ( n26839 , n26837 , n26838 );
not ( n26840 , n26837 );
and ( n26841 , n26840 , n25506 );
nor ( n26842 , n26839 , n26841 );
not ( n26843 , n26842 );
not ( n26844 , n26843 );
not ( n26845 , n19646 );
or ( n26846 , n26844 , n26845 );
nand ( n26847 , n21206 , n26842 );
nand ( n26848 , n26846 , n26847 );
buf ( n26849 , n24440 );
and ( n26850 , n26848 , n26849 );
not ( n26851 , n26848 );
not ( n26852 , n26849 );
and ( n26853 , n26851 , n26852 );
nor ( n26854 , n26850 , n26853 );
not ( n26855 , n26854 );
nand ( n26856 , n26836 , n26855 );
not ( n26857 , n16291 );
and ( n26858 , n26856 , n26857 );
not ( n26859 , n26856 );
and ( n26860 , n26859 , n16291 );
nor ( n26861 , n26858 , n26860 );
not ( n26862 , n26861 );
buf ( n26863 , n8132 );
not ( n26864 , n26863 );
not ( n26865 , n26864 );
not ( n26866 , n24876 );
or ( n26867 , n26865 , n26866 );
nand ( n26868 , n26567 , n26863 );
nand ( n26869 , n26867 , n26868 );
and ( n26870 , n26869 , n26121 );
not ( n26871 , n26869 );
and ( n26872 , n26871 , n26573 );
nor ( n26873 , n26870 , n26872 );
buf ( n26874 , n8221 );
not ( n26875 , n26874 );
not ( n26876 , n20584 );
or ( n26877 , n26875 , n26876 );
or ( n26878 , n6961 , n26874 );
nand ( n26879 , n26877 , n26878 );
buf ( n26880 , n19187 );
and ( n26881 , n26879 , n26880 );
not ( n26882 , n26879 );
and ( n26883 , n26882 , n19174 );
nor ( n26884 , n26881 , n26883 );
nand ( n26885 , n26873 , n26884 );
not ( n26886 , n26885 );
not ( n26887 , n16379 );
and ( n26888 , n26886 , n26887 );
and ( n26889 , n26885 , n16379 );
nor ( n26890 , n26888 , n26889 );
not ( n26891 , n26890 );
and ( n26892 , n26862 , n26891 );
and ( n26893 , n26861 , n26890 );
nor ( n26894 , n26892 , n26893 );
not ( n26895 , n26894 );
and ( n26896 , n26825 , n26895 );
and ( n26897 , n26824 , n26894 );
nor ( n26898 , n26896 , n26897 );
not ( n26899 , n26898 );
or ( n26900 , n26755 , n26899 );
not ( n26901 , n26754 );
not ( n26902 , n26894 );
not ( n26903 , n26824 );
or ( n26904 , n26902 , n26903 );
not ( n26905 , n26824 );
not ( n26906 , n26894 );
nand ( n26907 , n26905 , n26906 );
nand ( n26908 , n26904 , n26907 );
nand ( n26909 , n26901 , n26908 );
nand ( n26910 , n26900 , n26909 );
not ( n26911 , n15512 );
xor ( n26912 , n7287 , n7308 );
xnor ( n26913 , n26912 , n26791 );
not ( n26914 , n26913 );
not ( n26915 , n26914 );
or ( n26916 , n26911 , n26915 );
or ( n26917 , n25121 , n15512 );
nand ( n26918 , n26916 , n26917 );
and ( n26919 , n26918 , n25127 );
not ( n26920 , n26918 );
and ( n26921 , n26920 , n25128 );
nor ( n26922 , n26919 , n26921 );
not ( n26923 , n26922 );
not ( n26924 , n13165 );
not ( n26925 , n7065 );
not ( n26926 , n21191 );
or ( n26927 , n26925 , n26926 );
or ( n26928 , n21191 , n7065 );
nand ( n26929 , n26927 , n26928 );
not ( n26930 , n26929 );
or ( n26931 , n26924 , n26930 );
not ( n26932 , n26929 );
nand ( n26933 , n26932 , n13157 );
nand ( n26934 , n26931 , n26933 );
nand ( n26935 , n26923 , n26934 );
not ( n26936 , n26935 );
buf ( n26937 , n6813 );
not ( n26938 , n26937 );
not ( n26939 , n16491 );
or ( n26940 , n26938 , n26939 );
not ( n26941 , n16488 );
or ( n26942 , n26941 , n26937 );
nand ( n26943 , n26940 , n26942 );
buf ( n26944 , n16536 );
and ( n26945 , n26943 , n26944 );
not ( n26946 , n26943 );
and ( n26947 , n26946 , n16539 );
nor ( n26948 , n26945 , n26947 );
not ( n26949 , n26948 );
not ( n26950 , n26949 );
and ( n26951 , n26936 , n26950 );
and ( n26952 , n26935 , n26949 );
nor ( n26953 , n26951 , n26952 );
not ( n26954 , n26953 );
not ( n26955 , n9279 );
not ( n26956 , n12901 );
or ( n26957 , n26955 , n26956 );
or ( n26958 , n12901 , n9279 );
nand ( n26959 , n26957 , n26958 );
buf ( n26960 , n19026 );
and ( n26961 , n26959 , n26960 );
not ( n26962 , n26959 );
buf ( n26963 , n15830 );
and ( n26964 , n26962 , n26963 );
nor ( n26965 , n26961 , n26964 );
not ( n26966 , n12242 );
not ( n26967 , n9543 );
or ( n26968 , n26966 , n26967 );
or ( n26969 , n9543 , n12242 );
nand ( n26970 , n26968 , n26969 );
and ( n26971 , n26970 , n7256 );
not ( n26972 , n26970 );
and ( n26973 , n26972 , n7255 );
nor ( n26974 , n26971 , n26973 );
not ( n26975 , n26974 );
nand ( n26976 , n26965 , n26975 );
not ( n26977 , n13228 );
not ( n26978 , n9237 );
and ( n26979 , n26977 , n26978 );
and ( n26980 , n13228 , n9237 );
nor ( n26981 , n26979 , n26980 );
buf ( n26982 , n11592 );
xor ( n26983 , n26981 , n26982 );
buf ( n26984 , n26983 );
and ( n26985 , n26976 , n26984 );
not ( n26986 , n26976 );
not ( n26987 , n26984 );
and ( n26988 , n26986 , n26987 );
nor ( n26989 , n26985 , n26988 );
not ( n26990 , n26989 );
or ( n26991 , n26954 , n26990 );
or ( n26992 , n26989 , n26953 );
nand ( n26993 , n26991 , n26992 );
not ( n26994 , n20062 );
not ( n26995 , n26994 );
not ( n26996 , n21411 );
and ( n26997 , n26995 , n26996 );
and ( n26998 , n20057 , n21411 );
nor ( n26999 , n26997 , n26998 );
and ( n27000 , n26999 , n24392 );
not ( n27001 , n26999 );
buf ( n27002 , n24390 );
not ( n27003 , n27002 );
and ( n27004 , n27001 , n27003 );
nor ( n27005 , n27000 , n27004 );
buf ( n27006 , n27005 );
not ( n27007 , n27006 );
xor ( n27008 , n7339 , n9950 );
not ( n27009 , n9974 );
xnor ( n27010 , n27008 , n27009 );
nand ( n27011 , n27007 , n27010 );
not ( n27012 , n16285 );
buf ( n27013 , n18581 );
and ( n27014 , n27013 , n19670 );
not ( n27015 , n27013 );
xor ( n27016 , n11847 , n11856 );
not ( n27017 , n11866 );
xnor ( n27018 , n27016 , n27017 );
and ( n27019 , n27015 , n27018 );
nor ( n27020 , n27014 , n27019 );
not ( n27021 , n27020 );
and ( n27022 , n27012 , n27021 );
and ( n27023 , n16285 , n27020 );
nor ( n27024 , n27022 , n27023 );
and ( n27025 , n27011 , n27024 );
not ( n27026 , n27011 );
not ( n27027 , n27024 );
and ( n27028 , n27026 , n27027 );
nor ( n27029 , n27025 , n27028 );
and ( n27030 , n26993 , n27029 );
not ( n27031 , n26993 );
not ( n27032 , n27029 );
and ( n27033 , n27031 , n27032 );
nor ( n27034 , n27030 , n27033 );
not ( n27035 , n27034 );
not ( n27036 , n11924 );
and ( n27037 , n10272 , n13317 );
not ( n27038 , n10272 );
and ( n27039 , n27038 , n13318 );
or ( n27040 , n27037 , n27039 );
not ( n27041 , n27040 );
and ( n27042 , n27036 , n27041 );
and ( n27043 , n11924 , n27040 );
nor ( n27044 , n27042 , n27043 );
not ( n27045 , n27044 );
not ( n27046 , n27045 );
xor ( n27047 , n10476 , n14056 );
xnor ( n27048 , n27047 , n8074 );
not ( n27049 , n10557 );
not ( n27050 , n12200 );
or ( n27051 , n27049 , n27050 );
or ( n27052 , n25843 , n10557 );
nand ( n27053 , n27051 , n27052 );
and ( n27054 , n27053 , n25512 );
not ( n27055 , n27053 );
and ( n27056 , n27055 , n25513 );
or ( n27057 , n27054 , n27056 );
not ( n27058 , n27057 );
nand ( n27059 , n27048 , n27058 );
not ( n27060 , n27059 );
or ( n27061 , n27046 , n27060 );
or ( n27062 , n27059 , n27045 );
nand ( n27063 , n27061 , n27062 );
not ( n27064 , n27063 );
not ( n27065 , n11332 );
not ( n27066 , n25202 );
or ( n27067 , n27065 , n27066 );
or ( n27068 , n25202 , n11332 );
nand ( n27069 , n27067 , n27068 );
not ( n27070 , n27069 );
not ( n27071 , n23923 );
and ( n27072 , n27070 , n27071 );
and ( n27073 , n27069 , n23923 );
nor ( n27074 , n27072 , n27073 );
xor ( n27075 , n14065 , n26210 );
not ( n27076 , n21783 );
xnor ( n27077 , n27075 , n27076 );
nand ( n27078 , n27074 , n27077 );
not ( n27079 , n27078 );
not ( n27080 , n17810 );
not ( n27081 , n27080 );
xor ( n27082 , n27081 , n20686 );
xnor ( n27083 , n27082 , n12089 );
not ( n27084 , n27083 );
and ( n27085 , n27079 , n27084 );
not ( n27086 , n27074 );
not ( n27087 , n27086 );
nand ( n27088 , n27087 , n27077 );
and ( n27089 , n27088 , n27083 );
nor ( n27090 , n27085 , n27089 );
not ( n27091 , n27090 );
or ( n27092 , n27064 , n27091 );
or ( n27093 , n27090 , n27063 );
nand ( n27094 , n27092 , n27093 );
not ( n27095 , n27094 );
not ( n27096 , n27095 );
or ( n27097 , n27035 , n27096 );
not ( n27098 , n27034 );
nand ( n27099 , n27094 , n27098 );
nand ( n27100 , n27097 , n27099 );
not ( n27101 , n27100 );
not ( n27102 , n27101 );
and ( n27103 , n26910 , n27102 );
not ( n27104 , n26910 );
not ( n27105 , n27101 );
not ( n27106 , n27105 );
and ( n27107 , n27104 , n27106 );
nor ( n27108 , n27103 , n27107 );
or ( n27109 , n11062 , n17317 );
buf ( n27110 , n11017 );
not ( n27111 , n27110 );
and ( n27112 , n27109 , n27111 );
not ( n27113 , n27109 );
and ( n27114 , n27113 , n27110 );
nor ( n27115 , n27112 , n27114 );
not ( n27116 , n27115 );
not ( n27117 , n27116 );
not ( n27118 , n11750 );
or ( n27119 , n27117 , n27118 );
not ( n27120 , n27116 );
nand ( n27121 , n27120 , n11739 );
nand ( n27122 , n27119 , n27121 );
and ( n27123 , n27122 , n23812 );
not ( n27124 , n27122 );
buf ( n27125 , n23811 );
and ( n27126 , n27124 , n27125 );
nor ( n27127 , n27123 , n27126 );
nand ( n27128 , n27108 , n27127 );
or ( n27129 , n26692 , n27128 );
not ( n27130 , n27108 );
not ( n27131 , n26690 );
or ( n27132 , n27130 , n27131 );
buf ( n27133 , n22058 );
nor ( n27134 , n27127 , n27133 );
nand ( n27135 , n27132 , n27134 );
nand ( n27136 , n13766 , n16503 );
nand ( n27137 , n27129 , n27135 , n27136 );
buf ( n27138 , n27137 );
buf ( n27139 , n27138 );
not ( n27140 , n21933 );
not ( n27141 , n10641 );
or ( n27142 , n27140 , n27141 );
not ( n27143 , n21933 );
nand ( n27144 , n27143 , n10640 );
nand ( n27145 , n27142 , n27144 );
and ( n27146 , n27145 , n18794 );
not ( n27147 , n27145 );
and ( n27148 , n27147 , n18793 );
nor ( n27149 , n27146 , n27148 );
nand ( n27150 , n27149 , n24892 );
not ( n27151 , n27150 );
not ( n27152 , n12599 );
not ( n27153 , n23005 );
or ( n27154 , n27152 , n27153 );
or ( n27155 , n23005 , n12599 );
nand ( n27156 , n27154 , n27155 );
and ( n27157 , n27156 , n16184 );
not ( n27158 , n27156 );
and ( n27159 , n27158 , n16183 );
nor ( n27160 , n27157 , n27159 );
not ( n27161 , n27160 );
not ( n27162 , n27161 );
and ( n27163 , n27151 , n27162 );
and ( n27164 , n27150 , n27161 );
nor ( n27165 , n27163 , n27164 );
not ( n27166 , n27165 );
not ( n27167 , n6916 );
not ( n27168 , n23245 );
or ( n27169 , n27167 , n27168 );
not ( n27170 , n6916 );
not ( n27171 , n23244 );
nand ( n27172 , n27170 , n27171 );
nand ( n27173 , n27169 , n27172 );
not ( n27174 , n13324 );
and ( n27175 , n27173 , n27174 );
not ( n27176 , n27173 );
and ( n27177 , n27176 , n13324 );
nor ( n27178 , n27175 , n27177 );
not ( n27179 , n9219 );
not ( n27180 , n21162 );
and ( n27181 , n27179 , n27180 );
and ( n27182 , n9219 , n21162 );
nor ( n27183 , n27181 , n27182 );
and ( n27184 , n27183 , n15286 );
not ( n27185 , n27183 );
and ( n27186 , n27185 , n15282 );
nor ( n27187 , n27184 , n27186 );
nand ( n27188 , n27178 , n27187 );
not ( n27189 , n27188 );
not ( n27190 , n24951 );
or ( n27191 , n27189 , n27190 );
or ( n27192 , n24951 , n27188 );
nand ( n27193 , n27191 , n27192 );
not ( n27194 , n27193 );
not ( n27195 , n27194 );
not ( n27196 , n9489 );
not ( n27197 , n6834 );
not ( n27198 , n16536 );
or ( n27199 , n27197 , n27198 );
or ( n27200 , n16536 , n6834 );
nand ( n27201 , n27199 , n27200 );
not ( n27202 , n27201 );
and ( n27203 , n27196 , n27202 );
and ( n27204 , n9489 , n27201 );
nor ( n27205 , n27203 , n27204 );
buf ( n27206 , n18232 );
xor ( n27207 , n27206 , n14212 );
xnor ( n27208 , n27207 , n13902 );
nand ( n27209 , n27205 , n27208 );
not ( n27210 , n27209 );
not ( n27211 , n24920 );
and ( n27212 , n27210 , n27211 );
and ( n27213 , n27209 , n24920 );
nor ( n27214 , n27212 , n27213 );
not ( n27215 , n27214 );
not ( n27216 , n27215 );
or ( n27217 , n27195 , n27216 );
nand ( n27218 , n27214 , n27193 );
nand ( n27219 , n27217 , n27218 );
not ( n27220 , n27149 );
nand ( n27221 , n27160 , n27220 );
not ( n27222 , n27221 );
buf ( n27223 , n24883 );
not ( n27224 , n27223 );
and ( n27225 , n27222 , n27224 );
and ( n27226 , n27221 , n27223 );
nor ( n27227 , n27225 , n27226 );
not ( n27228 , n27227 );
and ( n27229 , n27219 , n27228 );
not ( n27230 , n27219 );
and ( n27231 , n27230 , n27227 );
nor ( n27232 , n27229 , n27231 );
not ( n27233 , n13571 );
not ( n27234 , n27233 );
not ( n27235 , n8458 );
not ( n27236 , n10060 );
or ( n27237 , n27235 , n27236 );
not ( n27238 , n8458 );
not ( n27239 , n10059 );
buf ( n27240 , n27239 );
nand ( n27241 , n27238 , n27240 );
nand ( n27242 , n27237 , n27241 );
not ( n27243 , n27242 );
or ( n27244 , n27234 , n27243 );
or ( n27245 , n27233 , n27242 );
nand ( n27246 , n27244 , n27245 );
not ( n27247 , n22587 );
not ( n27248 , n21030 );
or ( n27249 , n27247 , n27248 );
or ( n27250 , n21026 , n22587 );
nand ( n27251 , n27249 , n27250 );
not ( n27252 , n27251 );
not ( n27253 , n7425 );
and ( n27254 , n27252 , n27253 );
and ( n27255 , n27251 , n21037 );
nor ( n27256 , n27254 , n27255 );
nand ( n27257 , n27246 , n27256 );
not ( n27258 , n27257 );
not ( n27259 , n24722 );
and ( n27260 , n27258 , n27259 );
and ( n27261 , n27257 , n24722 );
nor ( n27262 , n27260 , n27261 );
not ( n27263 , n27262 );
not ( n27264 , n27263 );
not ( n27265 , n24643 );
not ( n27266 , n15476 );
not ( n27267 , n7334 );
or ( n27268 , n27266 , n27267 );
or ( n27269 , n7334 , n15476 );
nand ( n27270 , n27268 , n27269 );
buf ( n27271 , n25121 );
not ( n27272 , n27271 );
and ( n27273 , n27270 , n27272 );
not ( n27274 , n27270 );
and ( n27275 , n27274 , n27271 );
nor ( n27276 , n27273 , n27275 );
nand ( n27277 , n27276 , n24610 );
not ( n27278 , n27277 );
or ( n27279 , n27265 , n27278 );
or ( n27280 , n27277 , n24643 );
nand ( n27281 , n27279 , n27280 );
not ( n27282 , n27281 );
not ( n27283 , n27282 );
or ( n27284 , n27264 , n27283 );
nand ( n27285 , n27281 , n27262 );
nand ( n27286 , n27284 , n27285 );
not ( n27287 , n27286 );
and ( n27288 , n27232 , n27287 );
not ( n27289 , n27232 );
and ( n27290 , n27289 , n27286 );
nor ( n27291 , n27288 , n27290 );
not ( n27292 , n27291 );
not ( n27293 , n27292 );
or ( n27294 , n27166 , n27293 );
not ( n27295 , n27291 );
not ( n27296 , n27165 );
not ( n27297 , n27296 );
or ( n27298 , n27295 , n27297 );
nand ( n27299 , n27294 , n27298 );
not ( n27300 , n27299 );
buf ( n27301 , n13388 );
not ( n27302 , n27301 );
not ( n27303 , n22651 );
or ( n27304 , n27302 , n27303 );
not ( n27305 , n27301 );
nand ( n27306 , n27305 , n15647 );
nand ( n27307 , n27304 , n27306 );
and ( n27308 , n27307 , n15604 );
not ( n27309 , n27307 );
and ( n27310 , n27309 , n25996 );
nor ( n27311 , n27308 , n27310 );
not ( n27312 , n27311 );
not ( n27313 , n19799 );
not ( n27314 , n11281 );
or ( n27315 , n27313 , n27314 );
not ( n27316 , n19799 );
nand ( n27317 , n27316 , n6873 );
nand ( n27318 , n27315 , n27317 );
and ( n27319 , n27318 , n11287 );
not ( n27320 , n27318 );
and ( n27321 , n27320 , n11284 );
nor ( n27322 , n27319 , n27321 );
nand ( n27323 , n27312 , n27322 );
and ( n27324 , n27323 , n24334 );
not ( n27325 , n27323 );
and ( n27326 , n27325 , n24333 );
nor ( n27327 , n27324 , n27326 );
not ( n27328 , n27327 );
not ( n27329 , n27328 );
not ( n27330 , n12994 );
not ( n27331 , n16425 );
not ( n27332 , n16437 );
xor ( n27333 , n27331 , n27332 );
xnor ( n27334 , n27333 , n16440 );
not ( n27335 , n27334 );
or ( n27336 , n27330 , n27335 );
or ( n27337 , n27334 , n12994 );
nand ( n27338 , n27336 , n27337 );
and ( n27339 , n27338 , n23257 );
not ( n27340 , n27338 );
and ( n27341 , n27340 , n23258 );
nor ( n27342 , n27339 , n27341 );
buf ( n27343 , n6943 );
not ( n27344 , n27343 );
not ( n27345 , n27171 );
or ( n27346 , n27344 , n27345 );
or ( n27347 , n27171 , n27343 );
nand ( n27348 , n27346 , n27347 );
and ( n27349 , n27348 , n13320 );
not ( n27350 , n27348 );
and ( n27351 , n27350 , n13324 );
nor ( n27352 , n27349 , n27351 );
not ( n27353 , n27352 );
nand ( n27354 , n27342 , n27353 );
buf ( n27355 , n24396 );
xor ( n27356 , n27354 , n27355 );
not ( n27357 , n27356 );
not ( n27358 , n27357 );
or ( n27359 , n27329 , n27358 );
nand ( n27360 , n27356 , n27327 );
nand ( n27361 , n27359 , n27360 );
xor ( n27362 , n8579 , n18898 );
xnor ( n27363 , n27362 , n13218 );
not ( n27364 , n8482 );
not ( n27365 , n10061 );
or ( n27366 , n27364 , n27365 );
not ( n27367 , n8482 );
not ( n27368 , n10060 );
nand ( n27369 , n27367 , n27368 );
nand ( n27370 , n27366 , n27369 );
and ( n27371 , n27370 , n13571 );
not ( n27372 , n27370 );
and ( n27373 , n27372 , n16377 );
nor ( n27374 , n27371 , n27373 );
nand ( n27375 , n27363 , n27374 );
not ( n27376 , n27375 );
not ( n27377 , n24450 );
and ( n27378 , n27376 , n27377 );
and ( n27379 , n27375 , n24450 );
nor ( n27380 , n27378 , n27379 );
and ( n27381 , n27361 , n27380 );
not ( n27382 , n27361 );
not ( n27383 , n27380 );
and ( n27384 , n27382 , n27383 );
nor ( n27385 , n27381 , n27384 );
not ( n27386 , n27385 );
not ( n27387 , n24533 );
not ( n27388 , n27387 );
not ( n27389 , n27388 );
buf ( n27390 , n15392 );
not ( n27391 , n27390 );
not ( n27392 , n15389 );
and ( n27393 , n27391 , n27392 );
and ( n27394 , n27390 , n15389 );
nor ( n27395 , n27393 , n27394 );
and ( n27396 , n27395 , n20232 );
not ( n27397 , n27395 );
not ( n27398 , n13457 );
and ( n27399 , n27397 , n27398 );
nor ( n27400 , n27396 , n27399 );
not ( n27401 , n20284 );
and ( n27402 , n27400 , n27401 );
not ( n27403 , n27400 );
and ( n27404 , n27403 , n20284 );
nor ( n27405 , n27402 , n27404 );
not ( n27406 , n27405 );
not ( n27407 , n14005 );
buf ( n27408 , n27407 );
xor ( n27409 , n14796 , n27408 );
xnor ( n27410 , n27409 , n9630 );
not ( n27411 , n27410 );
nand ( n27412 , n27406 , n27411 );
not ( n27413 , n27412 );
or ( n27414 , n27389 , n27413 );
or ( n27415 , n27412 , n27388 );
nand ( n27416 , n27414 , n27415 );
not ( n27417 , n27416 );
buf ( n27418 , n11103 );
buf ( n27419 , n18737 );
xor ( n27420 , n27418 , n27419 );
xnor ( n27421 , n27420 , n18780 );
not ( n27422 , n27421 );
buf ( n27423 , n21944 );
not ( n27424 , n27423 );
not ( n27425 , n27424 );
not ( n27426 , n10641 );
or ( n27427 , n27425 , n27426 );
nand ( n27428 , n18788 , n27423 );
nand ( n27429 , n27427 , n27428 );
buf ( n27430 , n25351 );
xnor ( n27431 , n27429 , n27430 );
not ( n27432 , n27431 );
nand ( n27433 , n27422 , n27432 );
not ( n27434 , n27433 );
not ( n27435 , n24552 );
and ( n27436 , n27434 , n27435 );
and ( n27437 , n27433 , n24552 );
nor ( n27438 , n27436 , n27437 );
not ( n27439 , n27438 );
or ( n27440 , n27417 , n27439 );
or ( n27441 , n27438 , n27416 );
nand ( n27442 , n27440 , n27441 );
not ( n27443 , n27442 );
or ( n27444 , n27386 , n27443 );
or ( n27445 , n27442 , n27385 );
nand ( n27446 , n27444 , n27445 );
buf ( n27447 , n27446 );
not ( n27448 , n27447 );
not ( n27449 , n27448 );
and ( n27450 , n27300 , n27449 );
not ( n27451 , n27447 );
and ( n27452 , n27299 , n27451 );
nor ( n27453 , n27450 , n27452 );
not ( n27454 , n27453 );
not ( n27455 , n10779 );
not ( n27456 , n27408 );
or ( n27457 , n27455 , n27456 );
nand ( n27458 , n14007 , n10775 );
nand ( n27459 , n27457 , n27458 );
not ( n27460 , n24834 );
and ( n27461 , n27459 , n27460 );
not ( n27462 , n27459 );
and ( n27463 , n27462 , n24834 );
nor ( n27464 , n27461 , n27463 );
not ( n27465 , n27464 );
nand ( n27466 , n27465 , n23055 );
not ( n27467 , n27466 );
not ( n27468 , n14832 );
not ( n27469 , n23386 );
or ( n27470 , n27468 , n27469 );
or ( n27471 , n23386 , n14832 );
nand ( n27472 , n27470 , n27471 );
and ( n27473 , n27472 , n8951 );
not ( n27474 , n27472 );
not ( n27475 , n20971 );
and ( n27476 , n27474 , n27475 );
nor ( n27477 , n27473 , n27476 );
not ( n27478 , n27477 );
not ( n27479 , n27478 );
and ( n27480 , n27467 , n27479 );
and ( n27481 , n27466 , n27478 );
nor ( n27482 , n27480 , n27481 );
buf ( n27483 , n27482 );
not ( n27484 , n27483 );
not ( n27485 , n23000 );
not ( n27486 , n27485 );
xor ( n27487 , n15066 , n11310 );
xor ( n27488 , n27487 , n11317 );
buf ( n27489 , n27488 );
xor ( n27490 , n8041 , n27489 );
xnor ( n27491 , n27490 , n12587 );
not ( n27492 , n27491 );
not ( n27493 , n20727 );
xor ( n27494 , n18572 , n18591 );
xor ( n27495 , n27494 , n18581 );
not ( n27496 , n27495 );
not ( n27497 , n27496 );
or ( n27498 , n27493 , n27497 );
or ( n27499 , n23310 , n20727 );
nand ( n27500 , n27498 , n27499 );
and ( n27501 , n27500 , n18645 );
not ( n27502 , n27500 );
and ( n27503 , n27502 , n18651 );
nor ( n27504 , n27501 , n27503 );
not ( n27505 , n27504 );
nand ( n27506 , n27492 , n27505 );
not ( n27507 , n27506 );
or ( n27508 , n27486 , n27507 );
nand ( n27509 , n27492 , n27505 );
or ( n27510 , n27509 , n27485 );
nand ( n27511 , n27508 , n27510 );
not ( n27512 , n27511 );
nand ( n27513 , n27464 , n27477 );
and ( n27514 , n27513 , n23024 );
not ( n27515 , n27513 );
and ( n27516 , n27515 , n23023 );
nor ( n27517 , n27514 , n27516 );
not ( n27518 , n27517 );
and ( n27519 , n27512 , n27518 );
and ( n27520 , n27511 , n27517 );
nor ( n27521 , n27519 , n27520 );
not ( n27522 , n27521 );
not ( n27523 , n22933 );
buf ( n27524 , n10237 );
not ( n27525 , n27524 );
not ( n27526 , n9651 );
not ( n27527 , n9343 );
or ( n27528 , n27526 , n27527 );
or ( n27529 , n9343 , n9651 );
nand ( n27530 , n27528 , n27529 );
not ( n27531 , n27530 );
or ( n27532 , n27525 , n27531 );
not ( n27533 , n27530 );
not ( n27534 , n10237 );
nand ( n27535 , n27533 , n27534 );
nand ( n27536 , n27532 , n27535 );
nand ( n27537 , n27536 , n22728 );
not ( n27538 , n27537 );
or ( n27539 , n27523 , n27538 );
or ( n27540 , n27537 , n22933 );
nand ( n27541 , n27539 , n27540 );
not ( n27542 , n27541 );
xor ( n27543 , n16919 , n20564 );
and ( n27544 , n27543 , n13500 );
not ( n27545 , n27543 );
and ( n27546 , n27545 , n13499 );
nor ( n27547 , n27544 , n27546 );
buf ( n27548 , n19897 );
not ( n27549 , n27548 );
not ( n27550 , n19819 );
or ( n27551 , n27549 , n27550 );
or ( n27552 , n19819 , n27548 );
nand ( n27553 , n27551 , n27552 );
and ( n27554 , n27553 , n19110 );
not ( n27555 , n27553 );
and ( n27556 , n27555 , n19829 );
nor ( n27557 , n27554 , n27556 );
not ( n27558 , n27557 );
nand ( n27559 , n27547 , n27558 );
not ( n27560 , n27559 );
not ( n27561 , n22867 );
and ( n27562 , n27560 , n27561 );
and ( n27563 , n27559 , n22867 );
nor ( n27564 , n27562 , n27563 );
not ( n27565 , n27564 );
or ( n27566 , n27542 , n27565 );
or ( n27567 , n27564 , n27541 );
nand ( n27568 , n27566 , n27567 );
xor ( n27569 , n12123 , n11059 );
xnor ( n27570 , n27569 , n8612 );
not ( n27571 , n27570 );
not ( n27572 , n13143 );
not ( n27573 , n15286 );
or ( n27574 , n27572 , n27573 );
not ( n27575 , n13143 );
nand ( n27576 , n27575 , n15282 );
nand ( n27577 , n27574 , n27576 );
and ( n27578 , n27577 , n15328 );
not ( n27579 , n27577 );
and ( n27580 , n27579 , n15334 );
nor ( n27581 , n27578 , n27580 );
nand ( n27582 , n27571 , n27581 );
not ( n27583 , n27582 );
not ( n27584 , n22912 );
and ( n27585 , n27583 , n27584 );
not ( n27586 , n27581 );
not ( n27587 , n27586 );
nand ( n27588 , n27587 , n27571 );
and ( n27589 , n27588 , n22912 );
nor ( n27590 , n27585 , n27589 );
not ( n27591 , n27590 );
and ( n27592 , n27568 , n27591 );
not ( n27593 , n27568 );
and ( n27594 , n27593 , n27590 );
nor ( n27595 , n27592 , n27594 );
not ( n27596 , n27595 );
or ( n27597 , n27522 , n27596 );
not ( n27598 , n27595 );
not ( n27599 , n27521 );
nand ( n27600 , n27598 , n27599 );
nand ( n27601 , n27597 , n27600 );
not ( n27602 , n27601 );
or ( n27603 , n27484 , n27602 );
or ( n27604 , n27601 , n27483 );
nand ( n27605 , n27603 , n27604 );
not ( n27606 , n27605 );
not ( n27607 , n7715 );
not ( n27608 , n9895 );
and ( n27609 , n27607 , n27608 );
and ( n27610 , n7715 , n9895 );
nor ( n27611 , n27609 , n27610 );
xor ( n27612 , n15205 , n27611 );
not ( n27613 , n27612 );
not ( n27614 , n16510 );
not ( n27615 , n12270 );
or ( n27616 , n27614 , n27615 );
or ( n27617 , n12270 , n16510 );
nand ( n27618 , n27616 , n27617 );
not ( n27619 , n19342 );
and ( n27620 , n27618 , n27619 );
not ( n27621 , n27618 );
not ( n27622 , n19346 );
and ( n27623 , n27621 , n27622 );
nor ( n27624 , n27620 , n27623 );
nand ( n27625 , n27613 , n27624 );
and ( n27626 , n27625 , n23217 );
not ( n27627 , n27625 );
and ( n27628 , n27627 , n23218 );
nor ( n27629 , n27626 , n27628 );
xor ( n27630 , n22172 , n24227 );
xnor ( n27631 , n27630 , n19209 );
not ( n27632 , n12522 );
not ( n27633 , n26740 );
or ( n27634 , n27632 , n27633 );
not ( n27635 , n12522 );
xor ( n27636 , n26729 , n26738 );
xor ( n27637 , n27636 , n23630 );
not ( n27638 , n27637 );
nand ( n27639 , n27635 , n27638 );
nand ( n27640 , n27634 , n27639 );
not ( n27641 , n15898 );
not ( n27642 , n27641 );
and ( n27643 , n27640 , n27642 );
not ( n27644 , n27640 );
buf ( n27645 , n25953 );
and ( n27646 , n27644 , n27645 );
nor ( n27647 , n27643 , n27646 );
not ( n27648 , n27647 );
nand ( n27649 , n27631 , n27648 );
not ( n27650 , n23095 );
and ( n27651 , n27649 , n27650 );
not ( n27652 , n27649 );
and ( n27653 , n27652 , n23095 );
nor ( n27654 , n27651 , n27653 );
xor ( n27655 , n27629 , n27654 );
not ( n27656 , n12384 );
not ( n27657 , n16948 );
or ( n27658 , n27656 , n27657 );
or ( n27659 , n17592 , n12384 );
nand ( n27660 , n27658 , n27659 );
and ( n27661 , n27660 , n15370 );
not ( n27662 , n27660 );
and ( n27663 , n27662 , n16955 );
nor ( n27664 , n27661 , n27663 );
not ( n27665 , n27664 );
not ( n27666 , n7249 );
not ( n27667 , n25060 );
not ( n27668 , n27667 );
or ( n27669 , n27666 , n27668 );
not ( n27670 , n7249 );
nand ( n27671 , n27670 , n25060 );
nand ( n27672 , n27669 , n27671 );
not ( n27673 , n22145 );
and ( n27674 , n27672 , n27673 );
not ( n27675 , n27672 );
not ( n27676 , n22141 );
and ( n27677 , n27675 , n27676 );
nor ( n27678 , n27674 , n27677 );
not ( n27679 , n27678 );
nand ( n27680 , n27665 , n27679 );
not ( n27681 , n27680 );
not ( n27682 , n27681 );
not ( n27683 , n23260 );
not ( n27684 , n27683 );
or ( n27685 , n27682 , n27684 );
nand ( n27686 , n23260 , n27680 );
nand ( n27687 , n27685 , n27686 );
xor ( n27688 , n27655 , n27687 );
not ( n27689 , n27688 );
not ( n27690 , n7398 );
not ( n27691 , n13946 );
or ( n27692 , n27690 , n27691 );
nand ( n27693 , n15061 , n7395 );
nand ( n27694 , n27692 , n27693 );
and ( n27695 , n27694 , n27009 );
not ( n27696 , n27694 );
and ( n27697 , n27696 , n9974 );
nor ( n27698 , n27695 , n27697 );
buf ( n27699 , n25449 );
and ( n27700 , n25453 , n27699 );
not ( n27701 , n25453 );
and ( n27702 , n27701 , n25450 );
nor ( n27703 , n27700 , n27702 );
and ( n27704 , n27703 , n25697 );
not ( n27705 , n27703 );
buf ( n27706 , n25696 );
and ( n27707 , n27705 , n27706 );
or ( n27708 , n27704 , n27707 );
buf ( n27709 , n25912 );
and ( n27710 , n27708 , n27709 );
not ( n27711 , n27708 );
not ( n27712 , n27709 );
and ( n27713 , n27711 , n27712 );
nor ( n27714 , n27710 , n27713 );
not ( n27715 , n27714 );
nand ( n27716 , n27698 , n27715 );
not ( n27717 , n27716 );
not ( n27718 , n23401 );
or ( n27719 , n27717 , n27718 );
or ( n27720 , n23401 , n27716 );
nand ( n27721 , n27719 , n27720 );
not ( n27722 , n27721 );
not ( n27723 , n27722 );
xor ( n27724 , n13107 , n8441 );
xnor ( n27725 , n27724 , n21521 );
buf ( n27726 , n11669 );
not ( n27727 , n27726 );
not ( n27728 , n22919 );
or ( n27729 , n27727 , n27728 );
or ( n27730 , n22919 , n27726 );
nand ( n27731 , n27729 , n27730 );
and ( n27732 , n27731 , n14494 );
not ( n27733 , n27731 );
and ( n27734 , n27733 , n10377 );
nor ( n27735 , n27732 , n27734 );
not ( n27736 , n27735 );
nand ( n27737 , n27725 , n27736 );
not ( n27738 , n27737 );
not ( n27739 , n23389 );
and ( n27740 , n27738 , n27739 );
nand ( n27741 , n27725 , n27736 );
and ( n27742 , n27741 , n23389 );
nor ( n27743 , n27740 , n27742 );
not ( n27744 , n27743 );
not ( n27745 , n27744 );
or ( n27746 , n27723 , n27745 );
nand ( n27747 , n27743 , n27721 );
nand ( n27748 , n27746 , n27747 );
and ( n27749 , n27689 , n27748 );
not ( n27750 , n27689 );
not ( n27751 , n27748 );
and ( n27752 , n27750 , n27751 );
nor ( n27753 , n27749 , n27752 );
buf ( n27754 , n27753 );
not ( n27755 , n27754 );
and ( n27756 , n27606 , n27755 );
and ( n27757 , n27605 , n27754 );
nor ( n27758 , n27756 , n27757 );
nand ( n27759 , n27454 , n27758 );
not ( n27760 , n16874 );
not ( n27761 , n21873 );
or ( n27762 , n27760 , n27761 );
or ( n27763 , n21873 , n16874 );
nand ( n27764 , n27762 , n27763 );
and ( n27765 , n27764 , n19658 );
not ( n27766 , n27764 );
not ( n27767 , n19658 );
and ( n27768 , n27766 , n27767 );
nor ( n27769 , n27765 , n27768 );
not ( n27770 , n20545 );
not ( n27771 , n11717 );
or ( n27772 , n27770 , n27771 );
or ( n27773 , n11717 , n20545 );
nand ( n27774 , n27772 , n27773 );
and ( n27775 , n27774 , n21834 );
not ( n27776 , n27774 );
and ( n27777 , n27776 , n21828 );
nor ( n27778 , n27775 , n27777 );
nand ( n27779 , n27769 , n27778 );
not ( n27780 , n27779 );
buf ( n27781 , n8886 );
xor ( n27782 , n27781 , n10463 );
not ( n27783 , n11180 );
not ( n27784 , n10418 );
or ( n27785 , n27783 , n27784 );
nand ( n27786 , n27785 , n11184 );
not ( n27787 , n27786 );
xnor ( n27788 , n27782 , n27787 );
not ( n27789 , n27788 );
not ( n27790 , n27789 );
or ( n27791 , n27780 , n27790 );
or ( n27792 , n27789 , n27779 );
nand ( n27793 , n27791 , n27792 );
not ( n27794 , n27793 );
and ( n27795 , n10234 , n10231 );
not ( n27796 , n10234 );
buf ( n27797 , n10230 );
and ( n27798 , n27796 , n27797 );
nor ( n27799 , n27795 , n27798 );
xor ( n27800 , n27799 , n19129 );
xnor ( n27801 , n27800 , n15843 );
not ( n27802 , n27801 );
xor ( n27803 , n21726 , n21733 );
xnor ( n27804 , n27803 , n21740 );
buf ( n27805 , n27804 );
not ( n27806 , n27805 );
buf ( n27807 , n16707 );
not ( n27808 , n27807 );
and ( n27809 , n27806 , n27808 );
and ( n27810 , n27805 , n27807 );
nor ( n27811 , n27809 , n27810 );
and ( n27812 , n27811 , n21780 );
not ( n27813 , n27811 );
not ( n27814 , n21780 );
and ( n27815 , n27813 , n27814 );
nor ( n27816 , n27812 , n27815 );
not ( n27817 , n27816 );
buf ( n27818 , n24758 );
and ( n27819 , n18108 , n27818 );
not ( n27820 , n18108 );
and ( n27821 , n27820 , n24759 );
nor ( n27822 , n27819 , n27821 );
and ( n27823 , n27822 , n25987 );
not ( n27824 , n27822 );
not ( n27825 , n22651 );
not ( n27826 , n27825 );
and ( n27827 , n27824 , n27826 );
nor ( n27828 , n27823 , n27827 );
nand ( n27829 , n27817 , n27828 );
not ( n27830 , n27829 );
or ( n27831 , n27802 , n27830 );
nand ( n27832 , n27828 , n27817 );
or ( n27833 , n27832 , n27801 );
nand ( n27834 , n27831 , n27833 );
not ( n27835 , n27834 );
not ( n27836 , n27769 );
nand ( n27837 , n27788 , n27836 );
not ( n27838 , n27837 );
not ( n27839 , n7309 );
not ( n27840 , n18187 );
or ( n27841 , n27839 , n27840 );
not ( n27842 , n7309 );
nand ( n27843 , n27842 , n21057 );
nand ( n27844 , n27841 , n27843 );
and ( n27845 , n27844 , n21105 );
not ( n27846 , n27844 );
and ( n27847 , n27846 , n21098 );
nor ( n27848 , n27845 , n27847 );
not ( n27849 , n27848 );
not ( n27850 , n27849 );
and ( n27851 , n27838 , n27850 );
and ( n27852 , n27837 , n27849 );
nor ( n27853 , n27851 , n27852 );
not ( n27854 , n27853 );
or ( n27855 , n27835 , n27854 );
or ( n27856 , n27853 , n27834 );
nand ( n27857 , n27855 , n27856 );
not ( n27858 , n21155 );
not ( n27859 , n10854 );
or ( n27860 , n27858 , n27859 );
not ( n27861 , n21155 );
nand ( n27862 , n27861 , n9220 );
nand ( n27863 , n27860 , n27862 );
and ( n27864 , n27863 , n15287 );
not ( n27865 , n27863 );
and ( n27866 , n27865 , n10896 );
nor ( n27867 , n27864 , n27866 );
not ( n27868 , n18950 );
not ( n27869 , n27868 );
xor ( n27870 , n7124 , n7130 );
xnor ( n27871 , n27870 , n7143 );
not ( n27872 , n27871 );
not ( n27873 , n27872 );
or ( n27874 , n27869 , n27873 );
not ( n27875 , n7144 );
or ( n27876 , n27875 , n27868 );
nand ( n27877 , n27874 , n27876 );
and ( n27878 , n27877 , n15850 );
not ( n27879 , n27877 );
and ( n27880 , n27879 , n20505 );
nor ( n27881 , n27878 , n27880 );
nand ( n27882 , n27867 , n27881 );
not ( n27883 , n27882 );
buf ( n27884 , n15490 );
not ( n27885 , n27884 );
not ( n27886 , n7335 );
or ( n27887 , n27885 , n27886 );
or ( n27888 , n7335 , n27884 );
nand ( n27889 , n27887 , n27888 );
and ( n27890 , n27889 , n7312 );
not ( n27891 , n27889 );
and ( n27892 , n27891 , n27271 );
nor ( n27893 , n27890 , n27892 );
not ( n27894 , n27893 );
and ( n27895 , n27883 , n27894 );
and ( n27896 , n27882 , n27893 );
nor ( n27897 , n27895 , n27896 );
not ( n27898 , n27897 );
buf ( n27899 , n13933 );
not ( n27900 , n27899 );
not ( n27901 , n27900 );
not ( n27902 , n24514 );
or ( n27903 , n27901 , n27902 );
not ( n27904 , n24514 );
nand ( n27905 , n27904 , n27899 );
nand ( n27906 , n27903 , n27905 );
not ( n27907 , n27906 );
not ( n27908 , n24522 );
or ( n27909 , n27907 , n27908 );
or ( n27910 , n19889 , n27906 );
nand ( n27911 , n27909 , n27910 );
not ( n27912 , n27911 );
not ( n27913 , n13552 );
not ( n27914 , n7628 );
or ( n27915 , n27913 , n27914 );
or ( n27916 , n7628 , n13552 );
nand ( n27917 , n27915 , n27916 );
and ( n27918 , n27917 , n26620 );
not ( n27919 , n27917 );
and ( n27920 , n27919 , n26623 );
nor ( n27921 , n27918 , n27920 );
not ( n27922 , n27921 );
buf ( n27923 , n14461 );
not ( n27924 , n27923 );
not ( n27925 , n10697 );
or ( n27926 , n27924 , n27925 );
not ( n27927 , n24190 );
or ( n27928 , n27927 , n27923 );
nand ( n27929 , n27926 , n27928 );
not ( n27930 , n27929 );
buf ( n27931 , n10739 );
not ( n27932 , n27931 );
and ( n27933 , n27930 , n27932 );
and ( n27934 , n27931 , n27929 );
nor ( n27935 , n27933 , n27934 );
nand ( n27936 , n27922 , n27935 );
not ( n27937 , n27936 );
or ( n27938 , n27912 , n27937 );
or ( n27939 , n27936 , n27911 );
nand ( n27940 , n27938 , n27939 );
not ( n27941 , n27940 );
or ( n27942 , n27898 , n27941 );
or ( n27943 , n27940 , n27897 );
nand ( n27944 , n27942 , n27943 );
not ( n27945 , n12501 );
not ( n27946 , n27637 );
or ( n27947 , n27945 , n27946 );
not ( n27948 , n12501 );
nand ( n27949 , n27948 , n27638 );
nand ( n27950 , n27947 , n27949 );
and ( n27951 , n27950 , n15898 );
not ( n27952 , n27950 );
and ( n27953 , n27952 , n27645 );
nor ( n27954 , n27951 , n27953 );
not ( n27955 , n27954 );
not ( n27956 , n7172 );
not ( n27957 , n19805 );
or ( n27958 , n27956 , n27957 );
not ( n27959 , n7172 );
nand ( n27960 , n27959 , n25051 );
nand ( n27961 , n27958 , n27960 );
and ( n27962 , n27961 , n25778 );
not ( n27963 , n27961 );
and ( n27964 , n27963 , n25774 );
nor ( n27965 , n27962 , n27964 );
not ( n27966 , n27965 );
nand ( n27967 , n27955 , n27966 );
not ( n27968 , n27967 );
and ( n27969 , n19172 , n17692 );
not ( n27970 , n19172 );
and ( n27971 , n27970 , n13320 );
nor ( n27972 , n27969 , n27971 );
not ( n27973 , n17698 );
and ( n27974 , n27972 , n27973 );
not ( n27975 , n27972 );
and ( n27976 , n27975 , n17698 );
nor ( n27977 , n27974 , n27976 );
buf ( n27978 , n27977 );
not ( n27979 , n27978 );
and ( n27980 , n27968 , n27979 );
and ( n27981 , n27967 , n27978 );
nor ( n27982 , n27980 , n27981 );
and ( n27983 , n27944 , n27982 );
not ( n27984 , n27944 );
not ( n27985 , n27982 );
and ( n27986 , n27984 , n27985 );
nor ( n27987 , n27983 , n27986 );
and ( n27988 , n27857 , n27987 );
not ( n27989 , n27857 );
not ( n27990 , n27987 );
and ( n27991 , n27989 , n27990 );
nor ( n27992 , n27988 , n27991 );
not ( n27993 , n27992 );
not ( n27994 , n27993 );
not ( n27995 , n27994 );
or ( n27996 , n27794 , n27995 );
or ( n27997 , n27994 , n27793 );
nand ( n27998 , n27996 , n27997 );
xor ( n27999 , n17007 , n9221 );
xnor ( n28000 , n27999 , n9244 );
not ( n28001 , n12256 );
not ( n28002 , n9544 );
or ( n28003 , n28001 , n28002 );
not ( n28004 , n12256 );
nand ( n28005 , n28004 , n7207 );
nand ( n28006 , n28003 , n28005 );
and ( n28007 , n28006 , n12478 );
not ( n28008 , n28006 );
not ( n28009 , n7252 );
and ( n28010 , n28008 , n28009 );
nor ( n28011 , n28007 , n28010 );
nand ( n28012 , n28000 , n28011 );
not ( n28013 , n28012 );
not ( n28014 , n16092 );
not ( n28015 , n28014 );
not ( n28016 , n28015 );
not ( n28017 , n19374 );
not ( n28018 , n16098 );
or ( n28019 , n28017 , n28018 );
or ( n28020 , n16098 , n19374 );
nand ( n28021 , n28019 , n28020 );
not ( n28022 , n28021 );
or ( n28023 , n28016 , n28022 );
or ( n28024 , n28021 , n16093 );
nand ( n28025 , n28023 , n28024 );
not ( n28026 , n28025 );
and ( n28027 , n28013 , n28026 );
and ( n28028 , n28012 , n28025 );
nor ( n28029 , n28027 , n28028 );
not ( n28030 , n23272 );
buf ( n28031 , n12835 );
not ( n28032 , n28031 );
and ( n28033 , n28030 , n28032 );
and ( n28034 , n23272 , n28031 );
nor ( n28035 , n28033 , n28034 );
not ( n28036 , n12205 );
and ( n28037 , n28035 , n28036 );
not ( n28038 , n28035 );
and ( n28039 , n28038 , n12205 );
nor ( n28040 , n28037 , n28039 );
not ( n28041 , n28040 );
not ( n28042 , n13919 );
not ( n28043 , n24514 );
or ( n28044 , n28042 , n28043 );
or ( n28045 , n24514 , n13919 );
nand ( n28046 , n28044 , n28045 );
not ( n28047 , n28046 );
not ( n28048 , n24522 );
or ( n28049 , n28047 , n28048 );
or ( n28050 , n19889 , n28046 );
nand ( n28051 , n28049 , n28050 );
nand ( n28052 , n28041 , n28051 );
not ( n28053 , n6975 );
not ( n28054 , n9488 );
or ( n28055 , n28053 , n28054 );
or ( n28056 , n9488 , n6975 );
nand ( n28057 , n28055 , n28056 );
and ( n28058 , n28057 , n21214 );
not ( n28059 , n28057 );
and ( n28060 , n28059 , n9468 );
nor ( n28061 , n28058 , n28060 );
not ( n28062 , n28061 );
and ( n28063 , n28052 , n28062 );
not ( n28064 , n28052 );
not ( n28065 , n28062 );
and ( n28066 , n28064 , n28065 );
nor ( n28067 , n28063 , n28066 );
not ( n28068 , n28067 );
not ( n28069 , n28068 );
not ( n28070 , n15933 );
and ( n28071 , n8629 , n28070 );
not ( n28072 , n8629 );
and ( n28073 , n28072 , n15934 );
nor ( n28074 , n28071 , n28073 );
and ( n28075 , n28074 , n23988 );
not ( n28076 , n28074 );
buf ( n28077 , n23005 );
and ( n28078 , n28076 , n28077 );
nor ( n28079 , n28075 , n28078 );
not ( n28080 , n28079 );
xor ( n28081 , n23420 , n23439 );
buf ( n28082 , n23429 );
xnor ( n28083 , n28081 , n28082 );
buf ( n28084 , n28083 );
xor ( n28085 , n26513 , n28084 );
xnor ( n28086 , n28085 , n14970 );
nand ( n28087 , n28080 , n28086 );
not ( n28088 , n6591 );
not ( n28089 , n24323 );
or ( n28090 , n28088 , n28089 );
or ( n28091 , n24323 , n6591 );
nand ( n28092 , n28090 , n28091 );
and ( n28093 , n28092 , n18984 );
not ( n28094 , n28092 );
not ( n28095 , n18982 );
not ( n28096 , n28095 );
and ( n28097 , n28094 , n28096 );
nor ( n28098 , n28093 , n28097 );
and ( n28099 , n28087 , n28098 );
not ( n28100 , n28087 );
not ( n28101 , n28098 );
and ( n28102 , n28100 , n28101 );
nor ( n28103 , n28099 , n28102 );
not ( n28104 , n28103 );
not ( n28105 , n28104 );
or ( n28106 , n28069 , n28105 );
nand ( n28107 , n28103 , n28067 );
nand ( n28108 , n28106 , n28107 );
xor ( n28109 , n28029 , n28108 );
not ( n28110 , n24008 );
not ( n28111 , n28110 );
not ( n28112 , n18693 );
not ( n28113 , n20279 );
or ( n28114 , n28112 , n28113 );
or ( n28115 , n20279 , n18693 );
nand ( n28116 , n28114 , n28115 );
not ( n28117 , n28116 );
or ( n28118 , n28111 , n28117 );
or ( n28119 , n28116 , n28110 );
nand ( n28120 , n28118 , n28119 );
not ( n28121 , n28120 );
not ( n28122 , n8906 );
not ( n28123 , n18550 );
or ( n28124 , n28122 , n28123 );
or ( n28125 , n18550 , n8906 );
nand ( n28126 , n28124 , n28125 );
and ( n28127 , n28126 , n20632 );
not ( n28128 , n28126 );
and ( n28129 , n28128 , n25859 );
nor ( n28130 , n28127 , n28129 );
not ( n28131 , n28130 );
not ( n28132 , n12080 );
not ( n28133 , n17762 );
and ( n28134 , n28132 , n28133 );
and ( n28135 , n12080 , n17762 );
nor ( n28136 , n28134 , n28135 );
not ( n28137 , n28136 );
not ( n28138 , n12089 );
and ( n28139 , n28137 , n28138 );
and ( n28140 , n28136 , n12089 );
nor ( n28141 , n28139 , n28140 );
not ( n28142 , n28141 );
nand ( n28143 , n28131 , n28142 );
not ( n28144 , n28143 );
or ( n28145 , n28121 , n28144 );
or ( n28146 , n28143 , n28120 );
nand ( n28147 , n28145 , n28146 );
not ( n28148 , n28147 );
not ( n28149 , n14502 );
not ( n28150 , n12465 );
or ( n28151 , n28149 , n28150 );
or ( n28152 , n12465 , n14502 );
nand ( n28153 , n28151 , n28152 );
and ( n28154 , n28153 , n24762 );
not ( n28155 , n28153 );
and ( n28156 , n28155 , n24763 );
nor ( n28157 , n28154 , n28156 );
not ( n28158 , n28157 );
not ( n28159 , n14772 );
not ( n28160 , n9623 );
or ( n28161 , n28159 , n28160 );
not ( n28162 , n14772 );
nand ( n28163 , n28162 , n9629 );
nand ( n28164 , n28161 , n28163 );
and ( n28165 , n28164 , n14006 );
not ( n28166 , n28164 );
and ( n28167 , n28166 , n14007 );
nor ( n28168 , n28165 , n28167 );
not ( n28169 , n28168 );
nand ( n28170 , n28158 , n28169 );
not ( n28171 , n28170 );
not ( n28172 , n10237 );
not ( n28173 , n9658 );
not ( n28174 , n9343 );
or ( n28175 , n28173 , n28174 );
or ( n28176 , n9343 , n9658 );
nand ( n28177 , n28175 , n28176 );
not ( n28178 , n28177 );
or ( n28179 , n28172 , n28178 );
or ( n28180 , n10237 , n28177 );
nand ( n28181 , n28179 , n28180 );
not ( n28182 , n28181 );
and ( n28183 , n28171 , n28182 );
and ( n28184 , n28170 , n28181 );
nor ( n28185 , n28183 , n28184 );
not ( n28186 , n28185 );
or ( n28187 , n28148 , n28186 );
or ( n28188 , n28185 , n28147 );
nand ( n28189 , n28187 , n28188 );
xor ( n28190 , n28109 , n28189 );
buf ( n28191 , n28190 );
not ( n28192 , n28191 );
and ( n28193 , n27998 , n28192 );
not ( n28194 , n27998 );
and ( n28195 , n28194 , n28191 );
nor ( n28196 , n28193 , n28195 );
buf ( n28197 , n13744 );
nor ( n28198 , n28196 , n28197 );
not ( n28199 , n28198 );
or ( n28200 , n27759 , n28199 );
not ( n28201 , n28196 );
buf ( n28202 , n13745 );
not ( n28203 , n28202 );
nor ( n28204 , n28201 , n28203 );
nand ( n28205 , n27759 , n28204 );
buf ( n28206 , n13756 );
nand ( n28207 , n28206 , n21620 );
nand ( n28208 , n28200 , n28205 , n28207 );
buf ( n28209 , n28208 );
buf ( n28210 , n28209 );
not ( n28211 , n21193 );
not ( n28212 , n17170 );
not ( n28213 , n17039 );
or ( n28214 , n28212 , n28213 );
or ( n28215 , n17039 , n17170 );
nand ( n28216 , n28214 , n28215 );
not ( n28217 , n28216 );
or ( n28218 , n28211 , n28217 );
or ( n28219 , n28216 , n21194 );
nand ( n28220 , n28218 , n28219 );
not ( n28221 , n28220 );
xor ( n28222 , n12781 , n15743 );
xnor ( n28223 , n28222 , n14289 );
not ( n28224 , n16900 );
xor ( n28225 , n21860 , n9644 );
xnor ( n28226 , n28225 , n21871 );
buf ( n28227 , n28226 );
not ( n28228 , n28227 );
or ( n28229 , n28224 , n28228 );
or ( n28230 , n28227 , n16900 );
nand ( n28231 , n28229 , n28230 );
and ( n28232 , n28231 , n27767 );
not ( n28233 , n28231 );
and ( n28234 , n28233 , n19658 );
nor ( n28235 , n28232 , n28234 );
nand ( n28236 , n28223 , n28235 );
not ( n28237 , n28236 );
or ( n28238 , n28221 , n28237 );
not ( n28239 , n28236 );
not ( n28240 , n28220 );
nand ( n28241 , n28239 , n28240 );
nand ( n28242 , n28238 , n28241 );
not ( n28243 , n28242 );
not ( n28244 , n17949 );
not ( n28245 , n13546 );
or ( n28246 , n28244 , n28245 );
not ( n28247 , n17949 );
not ( n28248 , n13546 );
nand ( n28249 , n28247 , n28248 );
nand ( n28250 , n28246 , n28249 );
and ( n28251 , n28250 , n17003 );
not ( n28252 , n28250 );
and ( n28253 , n28252 , n17002 );
nor ( n28254 , n28251 , n28253 );
not ( n28255 , n28254 );
not ( n28256 , n28255 );
not ( n28257 , n18342 );
not ( n28258 , n17883 );
or ( n28259 , n28257 , n28258 );
or ( n28260 , n17883 , n18342 );
nand ( n28261 , n28259 , n28260 );
and ( n28262 , n9624 , n28261 );
not ( n28263 , n9624 );
not ( n28264 , n28261 );
and ( n28265 , n28263 , n28264 );
nor ( n28266 , n28262 , n28265 );
not ( n28267 , n28266 );
not ( n28268 , n22198 );
not ( n28269 , n13390 );
or ( n28270 , n28268 , n28269 );
not ( n28271 , n22198 );
not ( n28272 , n13390 );
nand ( n28273 , n28271 , n28272 );
nand ( n28274 , n28270 , n28273 );
and ( n28275 , n28274 , n13403 );
not ( n28276 , n28274 );
and ( n28277 , n28276 , n13399 );
nor ( n28278 , n28275 , n28277 );
nand ( n28279 , n28267 , n28278 );
not ( n28280 , n28279 );
or ( n28281 , n28256 , n28280 );
or ( n28282 , n28279 , n28255 );
nand ( n28283 , n28281 , n28282 );
not ( n28284 , n28283 );
not ( n28285 , n6739 );
not ( n28286 , n11777 );
or ( n28287 , n28285 , n28286 );
not ( n28288 , n6739 );
nand ( n28289 , n28288 , n14060 );
nand ( n28290 , n28287 , n28289 );
not ( n28291 , n11756 );
and ( n28292 , n28290 , n28291 );
not ( n28293 , n28290 );
and ( n28294 , n28293 , n9127 );
nor ( n28295 , n28292 , n28294 );
not ( n28296 , n12706 );
not ( n28297 , n7377 );
or ( n28298 , n28296 , n28297 );
not ( n28299 , n12706 );
xor ( n28300 , n7355 , n7375 );
not ( n28301 , n7365 );
xnor ( n28302 , n28300 , n28301 );
nand ( n28303 , n28299 , n28302 );
nand ( n28304 , n28298 , n28303 );
not ( n28305 , n19703 );
not ( n28306 , n16731 );
or ( n28307 , n28305 , n28306 );
not ( n28308 , n19702 );
nand ( n28309 , n28308 , n16727 );
nand ( n28310 , n28307 , n28309 );
not ( n28311 , n25089 );
and ( n28312 , n28310 , n28311 );
not ( n28313 , n28310 );
and ( n28314 , n28313 , n25090 );
nor ( n28315 , n28312 , n28314 );
buf ( n28316 , n6578 );
nand ( n28317 , n7412 , n28316 );
buf ( n28318 , n6579 );
buf ( n28319 , n28318 );
and ( n28320 , n28317 , n28319 );
not ( n28321 , n28317 );
not ( n28322 , n28318 );
and ( n28323 , n28321 , n28322 );
nor ( n28324 , n28320 , n28323 );
xor ( n28325 , n28315 , n28324 );
xnor ( n28326 , n28325 , n11941 );
buf ( n28327 , n28326 );
not ( n28328 , n28327 );
and ( n28329 , n28304 , n28328 );
not ( n28330 , n28304 );
and ( n28331 , n28330 , n28326 );
nor ( n28332 , n28329 , n28331 );
nand ( n28333 , n28295 , n28332 );
not ( n28334 , n28333 );
not ( n28335 , n21728 );
not ( n28336 , n10994 );
or ( n28337 , n28335 , n28336 );
not ( n28338 , n21728 );
nand ( n28339 , n28338 , n11007 );
nand ( n28340 , n28337 , n28339 );
and ( n28341 , n28340 , n10018 );
not ( n28342 , n28340 );
not ( n28343 , n10018 );
and ( n28344 , n28342 , n28343 );
nor ( n28345 , n28341 , n28344 );
not ( n28346 , n28345 );
not ( n28347 , n28346 );
and ( n28348 , n28334 , n28347 );
and ( n28349 , n28333 , n28346 );
nor ( n28350 , n28348 , n28349 );
not ( n28351 , n28350 );
or ( n28352 , n28284 , n28351 );
or ( n28353 , n28350 , n28283 );
nand ( n28354 , n28352 , n28353 );
not ( n28355 , n28354 );
not ( n28356 , n28355 );
not ( n28357 , n28223 );
nand ( n28358 , n28357 , n28240 );
not ( n28359 , n28358 );
and ( n28360 , n15472 , n7334 );
not ( n28361 , n15472 );
and ( n28362 , n28361 , n7335 );
or ( n28363 , n28360 , n28362 );
not ( n28364 , n22564 );
xnor ( n28365 , n28363 , n28364 );
not ( n28366 , n28365 );
not ( n28367 , n28366 );
and ( n28368 , n28359 , n28367 );
and ( n28369 , n28358 , n28366 );
nor ( n28370 , n28368 , n28369 );
not ( n28371 , n28370 );
not ( n28372 , n28371 );
or ( n28373 , n28356 , n28372 );
nand ( n28374 , n28370 , n28354 );
nand ( n28375 , n28373 , n28374 );
not ( n28376 , n11651 );
not ( n28377 , n22920 );
or ( n28378 , n28376 , n28377 );
not ( n28379 , n11651 );
nand ( n28380 , n28379 , n22919 );
nand ( n28381 , n28378 , n28380 );
and ( n28382 , n28381 , n10377 );
not ( n28383 , n28381 );
and ( n28384 , n28383 , n14494 );
nor ( n28385 , n28382 , n28384 );
not ( n28386 , n28385 );
not ( n28387 , n28386 );
not ( n28388 , n28387 );
not ( n28389 , n20758 );
not ( n28390 , n21688 );
or ( n28391 , n28389 , n28390 );
or ( n28392 , n20758 , n21688 );
nand ( n28393 , n28391 , n28392 );
and ( n28394 , n28393 , n23311 );
not ( n28395 , n28393 );
and ( n28396 , n28395 , n23314 );
nor ( n28397 , n28394 , n28396 );
not ( n28398 , n28397 );
not ( n28399 , n11130 );
not ( n28400 , n20477 );
not ( n28401 , n11104 );
or ( n28402 , n28400 , n28401 );
or ( n28403 , n11104 , n20477 );
nand ( n28404 , n28402 , n28403 );
not ( n28405 , n28404 );
and ( n28406 , n28399 , n28405 );
and ( n28407 , n11130 , n28404 );
nor ( n28408 , n28406 , n28407 );
not ( n28409 , n28408 );
nand ( n28410 , n28398 , n28409 );
not ( n28411 , n28410 );
or ( n28412 , n28388 , n28411 );
or ( n28413 , n28410 , n28387 );
nand ( n28414 , n28412 , n28413 );
not ( n28415 , n28414 );
not ( n28416 , n28415 );
not ( n28417 , n23346 );
not ( n28418 , n26515 );
or ( n28419 , n28417 , n28418 );
not ( n28420 , n23346 );
nand ( n28421 , n28420 , n7520 );
nand ( n28422 , n28419 , n28421 );
and ( n28423 , n28422 , n18550 );
not ( n28424 , n28422 );
and ( n28425 , n28424 , n26520 );
nor ( n28426 , n28423 , n28425 );
not ( n28427 , n28426 );
buf ( n28428 , n11147 );
not ( n28429 , n28428 );
not ( n28430 , n22141 );
or ( n28431 , n28429 , n28430 );
not ( n28432 , n28428 );
nand ( n28433 , n28432 , n22145 );
nand ( n28434 , n28431 , n28433 );
and ( n28435 , n28434 , n22189 );
not ( n28436 , n28434 );
and ( n28437 , n28436 , n22185 );
nor ( n28438 , n28435 , n28437 );
nand ( n28439 , n28427 , n28438 );
not ( n28440 , n28439 );
not ( n28441 , n8636 );
not ( n28442 , n15934 );
or ( n28443 , n28441 , n28442 );
or ( n28444 , n15934 , n8636 );
nand ( n28445 , n28443 , n28444 );
and ( n28446 , n28445 , n28077 );
not ( n28447 , n28445 );
and ( n28448 , n28447 , n23988 );
nor ( n28449 , n28446 , n28448 );
not ( n28450 , n28449 );
not ( n28451 , n28450 );
and ( n28452 , n28440 , n28451 );
and ( n28453 , n28439 , n28450 );
nor ( n28454 , n28452 , n28453 );
not ( n28455 , n28454 );
not ( n28456 , n28455 );
or ( n28457 , n28416 , n28456 );
nand ( n28458 , n28454 , n28414 );
nand ( n28459 , n28457 , n28458 );
and ( n28460 , n28375 , n28459 );
not ( n28461 , n28375 );
not ( n28462 , n28459 );
and ( n28463 , n28461 , n28462 );
nor ( n28464 , n28460 , n28463 );
not ( n28465 , n28464 );
not ( n28466 , n28465 );
or ( n28467 , n28243 , n28466 );
and ( n28468 , n28375 , n28459 );
not ( n28469 , n28375 );
and ( n28470 , n28469 , n28462 );
nor ( n28471 , n28468 , n28470 );
not ( n28472 , n28471 );
or ( n28473 , n28472 , n28242 );
nand ( n28474 , n28467 , n28473 );
not ( n28475 , n28474 );
buf ( n28476 , n15587 );
nor ( n28477 , n17666 , n28476 );
not ( n28478 , n28477 );
nand ( n28479 , n17666 , n28476 );
nand ( n28480 , n28478 , n28479 );
not ( n28481 , n28480 );
not ( n28482 , n19727 );
and ( n28483 , n28481 , n28482 );
not ( n28484 , n13618 );
and ( n28485 , n28480 , n28484 );
nor ( n28486 , n28483 , n28485 );
not ( n28487 , n28486 );
not ( n28488 , n28487 );
xor ( n28489 , n24379 , n16781 );
xnor ( n28490 , n28489 , n12730 );
not ( n28491 , n28490 );
not ( n28492 , n17198 );
not ( n28493 , n17037 );
or ( n28494 , n28492 , n28493 );
not ( n28495 , n17198 );
nand ( n28496 , n28495 , n17043 );
nand ( n28497 , n28494 , n28496 );
and ( n28498 , n28497 , n21191 );
not ( n28499 , n28497 );
and ( n28500 , n28499 , n21176 );
nor ( n28501 , n28498 , n28500 );
not ( n28502 , n28501 );
nand ( n28503 , n28491 , n28502 );
not ( n28504 , n28503 );
or ( n28505 , n28488 , n28504 );
not ( n28506 , n28501 );
nand ( n28507 , n28506 , n28491 );
or ( n28508 , n28507 , n28487 );
nand ( n28509 , n28505 , n28508 );
not ( n28510 , n28509 );
not ( n28511 , n10237 );
not ( n28512 , n9686 );
not ( n28513 , n9342 );
or ( n28514 , n28512 , n28513 );
or ( n28515 , n9342 , n9686 );
nand ( n28516 , n28514 , n28515 );
not ( n28517 , n28516 );
or ( n28518 , n28511 , n28517 );
not ( n28519 , n28516 );
nand ( n28520 , n28519 , n27534 );
nand ( n28521 , n28518 , n28520 );
not ( n28522 , n28521 );
not ( n28523 , n14801 );
not ( n28524 , n24702 );
not ( n28525 , n18369 );
or ( n28526 , n28524 , n28525 );
or ( n28527 , n18369 , n24702 );
nand ( n28528 , n28526 , n28527 );
not ( n28529 , n28528 );
or ( n28530 , n28523 , n28529 );
buf ( n28531 , n14797 );
or ( n28532 , n28528 , n28531 );
nand ( n28533 , n28530 , n28532 );
nand ( n28534 , n28522 , n28533 );
not ( n28535 , n28534 );
not ( n28536 , n14206 );
not ( n28537 , n18263 );
not ( n28538 , n14160 );
or ( n28539 , n28537 , n28538 );
or ( n28540 , n14160 , n18263 );
nand ( n28541 , n28539 , n28540 );
not ( n28542 , n28541 );
or ( n28543 , n28536 , n28542 );
or ( n28544 , n28541 , n14208 );
nand ( n28545 , n28543 , n28544 );
not ( n28546 , n28545 );
and ( n28547 , n28535 , n28546 );
and ( n28548 , n28534 , n28545 );
nor ( n28549 , n28547 , n28548 );
not ( n28550 , n28549 );
or ( n28551 , n28510 , n28550 );
or ( n28552 , n28549 , n28509 );
nand ( n28553 , n28551 , n28552 );
not ( n28554 , n21466 );
not ( n28555 , n7795 );
or ( n28556 , n28554 , n28555 );
not ( n28557 , n21466 );
nand ( n28558 , n28557 , n20016 );
nand ( n28559 , n28556 , n28558 );
and ( n28560 , n28559 , n20064 );
not ( n28561 , n28559 );
not ( n28562 , n20058 );
and ( n28563 , n28561 , n28562 );
nor ( n28564 , n28560 , n28563 );
not ( n28565 , n28564 );
not ( n28566 , n11130 );
not ( n28567 , n24617 );
nor ( n28568 , n11109 , n28567 );
not ( n28569 , n28568 );
nand ( n28570 , n11109 , n28567 );
nand ( n28571 , n28569 , n28570 );
not ( n28572 , n28571 );
and ( n28573 , n28566 , n28572 );
and ( n28574 , n11130 , n28571 );
nor ( n28575 , n28573 , n28574 );
not ( n28576 , n28575 );
nand ( n28577 , n28565 , n28576 );
not ( n28578 , n9923 );
not ( n28579 , n15503 );
or ( n28580 , n28578 , n28579 );
nand ( n28581 , n20981 , n9926 );
nand ( n28582 , n28580 , n28581 );
not ( n28583 , n28582 );
not ( n28584 , n15550 );
and ( n28585 , n28583 , n28584 );
and ( n28586 , n28582 , n15550 );
nor ( n28587 , n28585 , n28586 );
and ( n28588 , n28577 , n28587 );
not ( n28589 , n28577 );
not ( n28590 , n28587 );
and ( n28591 , n28589 , n28590 );
nor ( n28592 , n28588 , n28591 );
not ( n28593 , n28592 );
and ( n28594 , n28553 , n28593 );
not ( n28595 , n28553 );
and ( n28596 , n28595 , n28592 );
nor ( n28597 , n28594 , n28596 );
not ( n28598 , n28597 );
buf ( n28599 , n7239 );
not ( n28600 , n28599 );
not ( n28601 , n28600 );
not ( n28602 , n25060 );
not ( n28603 , n28602 );
or ( n28604 , n28601 , n28603 );
nand ( n28605 , n25777 , n28599 );
nand ( n28606 , n28604 , n28605 );
not ( n28607 , n27673 );
and ( n28608 , n28606 , n28607 );
not ( n28609 , n28606 );
not ( n28610 , n27676 );
and ( n28611 , n28609 , n28610 );
nor ( n28612 , n28608 , n28611 );
not ( n28613 , n12718 );
not ( n28614 , n7378 );
or ( n28615 , n28613 , n28614 );
not ( n28616 , n12718 );
nand ( n28617 , n28616 , n7435 );
nand ( n28618 , n28615 , n28617 );
not ( n28619 , n28618 );
not ( n28620 , n28327 );
and ( n28621 , n28619 , n28620 );
and ( n28622 , n28618 , n28327 );
nor ( n28623 , n28621 , n28622 );
nand ( n28624 , n28612 , n28623 );
not ( n28625 , n28624 );
not ( n28626 , n18334 );
xor ( n28627 , n23418 , n28626 );
xnor ( n28628 , n28627 , n20113 );
not ( n28629 , n28628 );
not ( n28630 , n28629 );
or ( n28631 , n28625 , n28630 );
or ( n28632 , n28629 , n28624 );
nand ( n28633 , n28631 , n28632 );
not ( n28634 , n28633 );
not ( n28635 , n28634 );
buf ( n28636 , n20329 );
buf ( n28637 , n17717 );
xor ( n28638 , n28636 , n28637 );
xnor ( n28639 , n28638 , n14664 );
buf ( n28640 , n12893 );
not ( n28641 , n28640 );
not ( n28642 , n28641 );
not ( n28643 , n16902 );
or ( n28644 , n28642 , n28643 );
nand ( n28645 , n16905 , n28640 );
nand ( n28646 , n28644 , n28645 );
and ( n28647 , n28646 , n14533 );
not ( n28648 , n28646 );
and ( n28649 , n28648 , n14534 );
nor ( n28650 , n28647 , n28649 );
not ( n28651 , n28650 );
nand ( n28652 , n28639 , n28651 );
not ( n28653 , n28652 );
not ( n28654 , n10091 );
not ( n28655 , n24239 );
or ( n28656 , n28654 , n28655 );
or ( n28657 , n24239 , n10091 );
nand ( n28658 , n28656 , n28657 );
and ( n28659 , n28658 , n18084 );
not ( n28660 , n28658 );
buf ( n28661 , n18070 );
xor ( n28662 , n28661 , n18078 );
xnor ( n28663 , n28662 , n18082 );
buf ( n28664 , n28663 );
and ( n28665 , n28660 , n28664 );
nor ( n28666 , n28659 , n28665 );
not ( n28667 , n28666 );
not ( n28668 , n28667 );
and ( n28669 , n28653 , n28668 );
nand ( n28670 , n28639 , n28651 );
and ( n28671 , n28670 , n28667 );
nor ( n28672 , n28669 , n28671 );
not ( n28673 , n28672 );
not ( n28674 , n28673 );
or ( n28675 , n28635 , n28674 );
nand ( n28676 , n28672 , n28633 );
nand ( n28677 , n28675 , n28676 );
not ( n28678 , n28677 );
and ( n28679 , n28598 , n28678 );
and ( n28680 , n28677 , n28597 );
nor ( n28681 , n28679 , n28680 );
buf ( n28682 , n28681 );
not ( n28683 , n28682 );
and ( n28684 , n28475 , n28683 );
and ( n28685 , n28474 , n28682 );
nor ( n28686 , n28684 , n28685 );
not ( n28687 , n28197 );
nand ( n28688 , n28686 , n28687 );
nand ( n28689 , n24543 , n27410 );
not ( n28690 , n28689 );
not ( n28691 , n27405 );
and ( n28692 , n28690 , n28691 );
and ( n28693 , n28689 , n27405 );
nor ( n28694 , n28692 , n28693 );
not ( n28695 , n28694 );
not ( n28696 , n28695 );
not ( n28697 , n27447 );
not ( n28698 , n28697 );
or ( n28699 , n28696 , n28698 );
not ( n28700 , n28695 );
nand ( n28701 , n28700 , n27447 );
nand ( n28702 , n28699 , n28701 );
buf ( n28703 , n19576 );
and ( n28704 , n28702 , n28703 );
not ( n28705 , n28702 );
not ( n28706 , n19584 );
not ( n28707 , n28706 );
and ( n28708 , n28705 , n28707 );
nor ( n28709 , n28704 , n28708 );
not ( n28710 , n28709 );
buf ( n28711 , n11948 );
xor ( n28712 , n7350 , n28711 );
not ( n28713 , n9974 );
xnor ( n28714 , n28712 , n28713 );
not ( n28715 , n28714 );
not ( n28716 , n28715 );
not ( n28717 , n12862 );
not ( n28718 , n23272 );
or ( n28719 , n28717 , n28718 );
not ( n28720 , n12862 );
nand ( n28721 , n28720 , n23268 );
nand ( n28722 , n28719 , n28721 );
and ( n28723 , n28722 , n12205 );
not ( n28724 , n28722 );
not ( n28725 , n12205 );
and ( n28726 , n28724 , n28725 );
nor ( n28727 , n28723 , n28726 );
not ( n28728 , n28727 );
not ( n28729 , n19826 );
buf ( n28730 , n20180 );
xor ( n28731 , n28729 , n28730 );
buf ( n28732 , n20218 );
xnor ( n28733 , n28731 , n28732 );
not ( n28734 , n28733 );
nand ( n28735 , n28728 , n28734 );
not ( n28736 , n28735 );
or ( n28737 , n28716 , n28736 );
not ( n28738 , n28727 );
nand ( n28739 , n28738 , n28734 );
or ( n28740 , n28739 , n28715 );
nand ( n28741 , n28737 , n28740 );
not ( n28742 , n28741 );
not ( n28743 , n12463 );
not ( n28744 , n19411 );
or ( n28745 , n28743 , n28744 );
not ( n28746 , n12463 );
not ( n28747 , n19411 );
nand ( n28748 , n28746 , n28747 );
nand ( n28749 , n28745 , n28748 );
not ( n28750 , n15395 );
and ( n28751 , n28749 , n28750 );
not ( n28752 , n28749 );
and ( n28753 , n28752 , n19416 );
nor ( n28754 , n28751 , n28753 );
not ( n28755 , n28754 );
not ( n28756 , n16600 );
not ( n28757 , n17191 );
or ( n28758 , n28756 , n28757 );
not ( n28759 , n16600 );
nand ( n28760 , n28759 , n17199 );
nand ( n28761 , n28758 , n28760 );
and ( n28762 , n28761 , n17203 );
not ( n28763 , n28761 );
and ( n28764 , n28763 , n17209 );
nor ( n28765 , n28762 , n28764 );
not ( n28766 , n28765 );
nand ( n28767 , n28755 , n28766 );
not ( n28768 , n28767 );
not ( n28769 , n8238 );
not ( n28770 , n15803 );
not ( n28771 , n8280 );
or ( n28772 , n28770 , n28771 );
nand ( n28773 , n8279 , n15799 );
nand ( n28774 , n28772 , n28773 );
not ( n28775 , n28774 );
and ( n28776 , n28769 , n28775 );
and ( n28777 , n24898 , n28774 );
nor ( n28778 , n28776 , n28777 );
not ( n28779 , n28778 );
not ( n28780 , n28779 );
and ( n28781 , n28768 , n28780 );
nand ( n28782 , n28755 , n28766 );
and ( n28783 , n28782 , n28779 );
nor ( n28784 , n28781 , n28783 );
not ( n28785 , n28784 );
buf ( n28786 , n15316 );
not ( n28787 , n28786 );
not ( n28788 , n6677 );
or ( n28789 , n28787 , n28788 );
not ( n28790 , n28786 );
nand ( n28791 , n28790 , n6676 );
nand ( n28792 , n28789 , n28791 );
and ( n28793 , n28792 , n17232 );
not ( n28794 , n28792 );
and ( n28795 , n28794 , n17229 );
nor ( n28796 , n28793 , n28795 );
not ( n28797 , n7733 );
not ( n28798 , n15743 );
or ( n28799 , n28797 , n28798 );
not ( n28800 , n7733 );
nand ( n28801 , n28800 , n15738 );
nand ( n28802 , n28799 , n28801 );
and ( n28803 , n28802 , n24026 );
not ( n28804 , n28802 );
and ( n28805 , n28804 , n15696 );
nor ( n28806 , n28803 , n28805 );
nand ( n28807 , n28796 , n28806 );
not ( n28808 , n19804 );
and ( n28809 , n9495 , n21103 );
not ( n28810 , n9495 );
and ( n28811 , n28810 , n21096 );
nor ( n28812 , n28809 , n28811 );
xnor ( n28813 , n28808 , n28812 );
and ( n28814 , n28807 , n28813 );
not ( n28815 , n28807 );
not ( n28816 , n28813 );
and ( n28817 , n28815 , n28816 );
nor ( n28818 , n28814 , n28817 );
not ( n28819 , n28818 );
or ( n28820 , n28785 , n28819 );
or ( n28821 , n28818 , n28784 );
nand ( n28822 , n28820 , n28821 );
not ( n28823 , n11033 );
not ( n28824 , n18903 );
or ( n28825 , n28823 , n28824 );
nand ( n28826 , n18906 , n11036 );
nand ( n28827 , n28825 , n28826 );
and ( n28828 , n28827 , n7932 );
not ( n28829 , n28827 );
and ( n28830 , n28829 , n13015 );
nor ( n28831 , n28828 , n28830 );
not ( n28832 , n28831 );
not ( n28833 , n21174 );
not ( n28834 , n10854 );
or ( n28835 , n28833 , n28834 );
nand ( n28836 , n9220 , n21175 );
nand ( n28837 , n28835 , n28836 );
not ( n28838 , n28837 );
not ( n28839 , n10896 );
and ( n28840 , n28838 , n28839 );
and ( n28841 , n28837 , n18021 );
nor ( n28842 , n28840 , n28841 );
not ( n28843 , n28842 );
nand ( n28844 , n28832 , n28843 );
not ( n28845 , n28844 );
xor ( n28846 , n24838 , n15120 );
xnor ( n28847 , n28846 , n23791 );
not ( n28848 , n28847 );
not ( n28849 , n28848 );
or ( n28850 , n28845 , n28849 );
or ( n28851 , n28848 , n28844 );
nand ( n28852 , n28850 , n28851 );
xor ( n28853 , n28822 , n28852 );
not ( n28854 , n28853 );
not ( n28855 , n21439 );
not ( n28856 , n7796 );
or ( n28857 , n28855 , n28856 );
or ( n28858 , n7796 , n21439 );
nand ( n28859 , n28857 , n28858 );
and ( n28860 , n28859 , n20065 );
not ( n28861 , n28859 );
and ( n28862 , n28861 , n20059 );
nor ( n28863 , n28860 , n28862 );
not ( n28864 , n28863 );
not ( n28865 , n28864 );
not ( n28866 , n6703 );
not ( n28867 , n26633 );
or ( n28868 , n28866 , n28867 );
or ( n28869 , n26636 , n6703 );
nand ( n28870 , n28868 , n28869 );
and ( n28871 , n28870 , n11778 );
not ( n28872 , n28870 );
and ( n28873 , n28872 , n14061 );
nor ( n28874 , n28871 , n28873 );
not ( n28875 , n28874 );
buf ( n28876 , n20561 );
not ( n28877 , n28876 );
not ( n28878 , n20558 );
and ( n28879 , n28877 , n28878 );
and ( n28880 , n28876 , n20558 );
nor ( n28881 , n28879 , n28880 );
xor ( n28882 , n28881 , n11717 );
and ( n28883 , n28882 , n21834 );
not ( n28884 , n28882 );
and ( n28885 , n28884 , n21828 );
nor ( n28886 , n28883 , n28885 );
nand ( n28887 , n28875 , n28886 );
not ( n28888 , n28887 );
or ( n28889 , n28865 , n28888 );
or ( n28890 , n28887 , n28864 );
nand ( n28891 , n28889 , n28890 );
nand ( n28892 , n28714 , n28727 );
not ( n28893 , n28892 );
not ( n28894 , n8770 );
buf ( n28895 , n24618 );
not ( n28896 , n28895 );
or ( n28897 , n28894 , n28896 );
or ( n28898 , n24620 , n8770 );
nand ( n28899 , n28897 , n28898 );
and ( n28900 , n28899 , n24186 );
not ( n28901 , n28899 );
and ( n28902 , n28901 , n24187 );
nor ( n28903 , n28900 , n28902 );
not ( n28904 , n28903 );
not ( n28905 , n28904 );
and ( n28906 , n28893 , n28905 );
and ( n28907 , n28892 , n28904 );
nor ( n28908 , n28906 , n28907 );
and ( n28909 , n28891 , n28908 );
not ( n28910 , n28891 );
not ( n28911 , n28908 );
and ( n28912 , n28910 , n28911 );
nor ( n28913 , n28909 , n28912 );
not ( n28914 , n28913 );
and ( n28915 , n28854 , n28914 );
not ( n28916 , n28854 );
and ( n28917 , n28916 , n28913 );
nor ( n28918 , n28915 , n28917 );
not ( n28919 , n28918 );
or ( n28920 , n28742 , n28919 );
not ( n28921 , n28741 );
not ( n28922 , n28913 );
not ( n28923 , n28853 );
or ( n28924 , n28922 , n28923 );
nand ( n28925 , n28854 , n28914 );
nand ( n28926 , n28924 , n28925 );
nand ( n28927 , n28921 , n28926 );
nand ( n28928 , n28920 , n28927 );
buf ( n28929 , n24991 );
and ( n28930 , n28928 , n28929 );
not ( n28931 , n28928 );
buf ( n28932 , n24985 );
and ( n28933 , n28931 , n28932 );
nor ( n28934 , n28930 , n28933 );
nand ( n28935 , n28710 , n28934 );
or ( n28936 , n28688 , n28935 );
buf ( n28937 , n13745 );
not ( n28938 , n28937 );
nor ( n28939 , n28686 , n28938 );
nand ( n28940 , n28939 , n28935 );
buf ( n28941 , n28206 );
buf ( n28942 , n10396 );
nand ( n28943 , n28941 , n28942 );
nand ( n28944 , n28936 , n28940 , n28943 );
buf ( n28945 , n28944 );
buf ( n28946 , n28945 );
endmodule

