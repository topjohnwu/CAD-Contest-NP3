//
// Conformal-LEC Version 16.10-d005 ( 21-Apr-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 ;
output n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 ;

wire n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
     n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
     n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , 
     n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , 
     n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , 
     n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , 
     n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , 
     n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
     n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
     n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
     n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
     n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
     n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
     n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
     n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
     n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
     n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
     n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
     n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
     n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
     n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
     n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
     n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
     n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
     n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
     n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
     n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
     n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
     n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
     n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
     n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
     n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , 
     n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , 
     n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
     n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , 
     n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
     n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , 
     n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
     n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
     n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
     n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , 
     n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
     n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
     n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
     n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
     n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
     n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
     n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
     n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
     n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
     n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
     n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
     n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
     n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , 
     n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , 
     n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , 
     n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , 
     n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , 
     n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , 
     n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , 
     n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
     n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , 
     n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , 
     n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , 
     n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , 
     n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , 
     n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , 
     n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , 
     n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , 
     n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , 
     n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , 
     n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , 
     n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , 
     n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , 
     n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , 
     n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
     n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
     n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
     n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
     n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
     n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
     n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
     n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
     n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
     n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
     n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
     n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
     n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
     n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
     n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , 
     n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , 
     n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
     n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , 
     n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , 
     n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , 
     n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , 
     n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , 
     n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , 
     n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , 
     n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , 
     n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
     n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , 
     n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , 
     n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , 
     n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
     n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , 
     n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , 
     n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
     n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , 
     n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , 
     n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , 
     n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , 
     n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , 
     n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , 
     n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , 
     n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , 
     n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , 
     n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , 
     n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , 
     n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , 
     n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , 
     n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , 
     n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , 
     n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , 
     n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , 
     n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , 
     n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
     n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , 
     n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , 
     n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , 
     n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , 
     n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , 
     n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , 
     n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , 
     n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , 
     n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , 
     n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , 
     n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , 
     n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , 
     n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , 
     n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , 
     n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , 
     n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , 
     n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , 
     n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , 
     n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , 
     n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , 
     n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , 
     n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , 
     n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , 
     n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , 
     n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , 
     n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , 
     n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , 
     n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , 
     n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , 
     n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , 
     n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , 
     n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , 
     n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , 
     n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , 
     n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , 
     n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , 
     n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , 
     n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , 
     n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , 
     n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , 
     n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , 
     n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , 
     n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , 
     n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , 
     n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , 
     n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , 
     n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , 
     n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , 
     n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , 
     n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , 
     n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , 
     n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , 
     n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , 
     n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , 
     n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , 
     n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , 
     n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , 
     n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , 
     n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , 
     n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , 
     n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , 
     n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , 
     n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , 
     n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , 
     n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , 
     n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , 
     n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , 
     n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , 
     n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , 
     n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , 
     n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , 
     n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , 
     n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , 
     n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , 
     n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , 
     n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , 
     n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , 
     n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , 
     n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , 
     n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , 
     n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , 
     n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , 
     n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , 
     n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , 
     n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , 
     n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , 
     n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , 
     n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , 
     n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , 
     n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , 
     n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , 
     n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , 
     n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , 
     n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , 
     n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , 
     n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , 
     n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , 
     n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , 
     n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , 
     n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , 
     n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , 
     n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , 
     n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , 
     n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , 
     n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , 
     n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , 
     n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , 
     n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , 
     n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , 
     n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , 
     n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , 
     n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , 
     n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , 
     n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , 
     n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , 
     n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , 
     n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , 
     n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , 
     n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , 
     n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , 
     n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , 
     n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , 
     n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , 
     n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , 
     n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , 
     n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , 
     n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , 
     n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , 
     n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , 
     n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , 
     n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , 
     n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , 
     n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , 
     n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , 
     n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , 
     n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , 
     n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , 
     n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , 
     n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , 
     n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , 
     n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , 
     n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , 
     n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , 
     n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , 
     n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , 
     n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , 
     n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , 
     n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , 
     n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , 
     n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , 
     n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , 
     n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , 
     n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , 
     n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , 
     n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , 
     n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , 
     n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , 
     n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , 
     n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , 
     n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , 
     n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , 
     n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , 
     n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , 
     n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , 
     n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , 
     n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , 
     n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , 
     n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , 
     n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , 
     n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , 
     n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , 
     n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , 
     n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , 
     n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , 
     n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , 
     n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , 
     n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , 
     n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , 
     n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , 
     n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , 
     n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , 
     n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , 
     n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , 
     n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , 
     n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , 
     n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , 
     n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , 
     n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , 
     n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , 
     n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , 
     n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , 
     n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , 
     n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , 
     n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , 
     n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , 
     n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , 
     n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , 
     n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , 
     n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , 
     n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , 
     n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , 
     n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , 
     n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , 
     n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , 
     n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , 
     n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , 
     n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , 
     n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , 
     n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , 
     n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , 
     n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , 
     n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , 
     n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , 
     n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , 
     n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , 
     n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , 
     n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , 
     n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , 
     n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , 
     n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , 
     n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , 
     n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , 
     n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , 
     n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , 
     n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , 
     n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , 
     n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , 
     n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , 
     n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , 
     n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , 
     n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , 
     n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , 
     n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , 
     n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , 
     n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , 
     n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , 
     n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , 
     n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , 
     n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , 
     n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , 
     n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , 
     n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , 
     n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , 
     n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , 
     n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , 
     n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , 
     n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , 
     n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , 
     n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , 
     n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , 
     n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , 
     n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , 
     n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , 
     n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , 
     n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , 
     n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , 
     n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , 
     n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , 
     n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , 
     n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , 
     n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , 
     n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , 
     n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , 
     n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , 
     n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , 
     n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , 
     n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , 
     n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , 
     n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , 
     n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , 
     n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , 
     n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , 
     n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , 
     n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , 
     n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , 
     n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , 
     n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , 
     n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , 
     n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , 
     n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , 
     n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , 
     n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , 
     n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , 
     n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , 
     n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , 
     n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , 
     n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , 
     n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , 
     n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , 
     n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , 
     n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , 
     n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , 
     n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , 
     n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , 
     n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , 
     n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , 
     n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , 
     n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , 
     n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , 
     n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , 
     n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , 
     n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , 
     n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , 
     n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , 
     n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , 
     n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , 
     n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , 
     n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , 
     n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , 
     n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , 
     n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , 
     n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , 
     n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , 
     n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , 
     n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , 
     n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , 
     n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , 
     n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , 
     n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , 
     n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , 
     n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , 
     n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , 
     n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , 
     n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , 
     n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , 
     n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , 
     n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , 
     n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , 
     n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , 
     n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , 
     n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , 
     n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , 
     n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , 
     n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , 
     n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , 
     n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , 
     n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , 
     n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , 
     n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , 
     n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , 
     n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , 
     n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , 
     n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , 
     n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , 
     n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , 
     n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , 
     n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , 
     n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , 
     n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , 
     n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , 
     n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , 
     n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , 
     n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , 
     n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , 
     n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , 
     n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , 
     n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , 
     n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , 
     n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , 
     n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , 
     n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , 
     n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , 
     n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , 
     n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , 
     n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , 
     n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , 
     n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , 
     n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , 
     n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , 
     n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , 
     n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , 
     n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , 
     n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , 
     n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , 
     n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , 
     n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , 
     n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , 
     n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , 
     n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , 
     n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , 
     n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , 
     n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , 
     n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , 
     n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , 
     n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , 
     n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , 
     n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , 
     n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , 
     n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , 
     n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , 
     n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , 
     n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , 
     n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , 
     n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , 
     n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , 
     n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , 
     n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , 
     n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , 
     n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , 
     n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , 
     n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , 
     n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , 
     n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , 
     n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , 
     n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , 
     n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , 
     n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , 
     n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , 
     n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , 
     n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , 
     n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , 
     n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , 
     n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , 
     n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , 
     n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , 
     n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , 
     n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , 
     n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , 
     n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , 
     n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , 
     n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , 
     n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , 
     n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , 
     n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , 
     n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , 
     n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , 
     n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , 
     n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , 
     n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , 
     n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , 
     n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , 
     n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , 
     n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , 
     n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , 
     n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , 
     n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , 
     n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , 
     n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , 
     n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , 
     n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , 
     n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , 
     n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , 
     n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , 
     n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , 
     n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , 
     n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , 
     n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , 
     n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , 
     n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , 
     n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , 
     n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , 
     n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , 
     n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , 
     n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , 
     n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , 
     n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , 
     n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , 
     n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , 
     n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , 
     n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , 
     n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , 
     n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , 
     n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , 
     n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , 
     n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , 
     n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , 
     n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , 
     n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , 
     n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , 
     n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , 
     n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , 
     n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , 
     n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , 
     n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , 
     n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , 
     n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , 
     n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , 
     n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , 
     n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , 
     n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , 
     n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , 
     n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , 
     n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , 
     n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , 
     n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , 
     n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , 
     n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , 
     n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , 
     n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , 
     n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , 
     n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , 
     n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , 
     n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , 
     n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , 
     n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , 
     n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , 
     n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , 
     n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , 
     n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , 
     n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , 
     n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , 
     n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , 
     n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , 
     n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , 
     n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , 
     n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , 
     n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , 
     n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , 
     n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , 
     n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , 
     n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , 
     n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , 
     n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , 
     n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , 
     n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , 
     n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , 
     n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , 
     n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , 
     n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , 
     n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , 
     n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , 
     n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , 
     n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , 
     n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , 
     n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , 
     n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , 
     n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , 
     n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , 
     n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , 
     n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , 
     n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , 
     n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , 
     n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , 
     n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , 
     n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , 
     n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , 
     n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , 
     n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , 
     n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , 
     n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , 
     n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , 
     n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , 
     n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , 
     n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , 
     n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , 
     n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , 
     n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , 
     n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , 
     n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , 
     n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , 
     n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , 
     n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , 
     n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , 
     n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , 
     n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , 
     n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , 
     n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , 
     n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , 
     n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , 
     n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , 
     n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , 
     n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , 
     n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , 
     n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , 
     n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , 
     n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , 
     n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , 
     n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , 
     n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , 
     n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , 
     n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , 
     n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , 
     n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , 
     n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , 
     n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , 
     n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , 
     n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , 
     n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , 
     n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , 
     n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , 
     n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , 
     n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , 
     n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , 
     n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , 
     n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , 
     n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , 
     n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , 
     n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , 
     n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , 
     n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , 
     n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , 
     n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , 
     n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , 
     n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , 
     n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , 
     n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , 
     n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , 
     n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , 
     n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , 
     n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , 
     n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , 
     n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , 
     n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , 
     n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , 
     n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , 
     n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , 
     n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , 
     n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , 
     n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , 
     n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , 
     n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , 
     n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , 
     n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , 
     n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , 
     n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , 
     n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , 
     n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , 
     n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , 
     n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , 
     n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , 
     n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , 
     n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , 
     n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , 
     n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , 
     n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , 
     n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , 
     n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , 
     n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , 
     n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , 
     n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , 
     n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , 
     n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , 
     n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , 
     n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , 
     n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , 
     n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , 
     n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , 
     n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , 
     n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , 
     n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , 
     n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , 
     n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , 
     n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , 
     n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , 
     n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , 
     n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , 
     n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , 
     n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , 
     n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , 
     n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , 
     n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , 
     n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , 
     n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , 
     n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , 
     n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , 
     n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , 
     n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , 
     n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , 
     n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , 
     n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , 
     n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , 
     n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , 
     n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , 
     n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , 
     n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , 
     n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , 
     n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , 
     n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , 
     n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , 
     n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , 
     n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , 
     n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , 
     n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , 
     n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , 
     n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , 
     n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , 
     n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , 
     n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , 
     n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , 
     n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , 
     n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , 
     n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , 
     n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , 
     n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , 
     n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , 
     n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , 
     n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , 
     n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , 
     n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , 
     n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , 
     n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , 
     n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , 
     n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , 
     n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , 
     n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , 
     n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , 
     n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , 
     n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , 
     n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , 
     n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , 
     n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , 
     n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , 
     n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , 
     n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , 
     n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , 
     n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , 
     n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , 
     n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , 
     n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , 
     n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , 
     n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , 
     n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , 
     n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , 
     n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , 
     n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , 
     n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , 
     n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , 
     n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , 
     n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , 
     n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , 
     n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , 
     n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , 
     n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , 
     n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , 
     n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , 
     n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , 
     n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , 
     n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , 
     n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , 
     n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , 
     n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , 
     n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , 
     n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , 
     n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , 
     n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , 
     n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , 
     n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , 
     n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , 
     n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , 
     n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , 
     n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , 
     n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , 
     n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , 
     n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , 
     n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , 
     n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , 
     n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , 
     n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , 
     n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , 
     n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , 
     n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , 
     n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , 
     n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , 
     n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , 
     n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , 
     n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , 
     n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , 
     n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , 
     n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , 
     n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , 
     n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , 
     n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , 
     n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , 
     n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , 
     n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , 
     n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , 
     n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , 
     n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , 
     n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , 
     n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , 
     n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , 
     n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , 
     n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , 
     n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , 
     n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , 
     n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , 
     n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , 
     n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , 
     n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , 
     n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , 
     n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , 
     n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , 
     n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , 
     n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , 
     n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , 
     n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , 
     n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , 
     n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , 
     n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , 
     n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , 
     n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , 
     n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , 
     n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , 
     n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , 
     n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , 
     n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , 
     n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , 
     n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , 
     n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , 
     n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , 
     n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , 
     n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , 
     n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , 
     n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , 
     n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , 
     n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , 
     n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , 
     n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , 
     n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , 
     n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , 
     n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , 
     n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , 
     n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , 
     n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , 
     n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , 
     n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , 
     n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , 
     n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , 
     n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , 
     n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , 
     n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , 
     n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , 
     n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , 
     n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , 
     n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , 
     n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , 
     n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , 
     n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , 
     n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , 
     n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , 
     n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , 
     n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , 
     n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , 
     n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , 
     n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , 
     n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , 
     n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , 
     n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , 
     n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , 
     n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , 
     n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , 
     n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , 
     n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , 
     n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , 
     n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , 
     n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , 
     n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , 
     n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , 
     n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , 
     n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , 
     n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , 
     n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , 
     n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , 
     n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , 
     n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , 
     n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , 
     n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , 
     n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , 
     n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , 
     n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , 
     n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , 
     n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , 
     n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , 
     n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , 
     n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , 
     n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , 
     n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , 
     n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , 
     n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , 
     n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , 
     n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , 
     n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , 
     n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , 
     n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , 
     n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , 
     n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , 
     n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , 
     n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , 
     n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , 
     n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , 
     n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , 
     n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , 
     n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , 
     n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , 
     n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , 
     n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , 
     n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , 
     n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , 
     n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , 
     n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , 
     n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , 
     n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , 
     n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , 
     n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , 
     n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , 
     n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , 
     n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , 
     n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , 
     n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , 
     n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , 
     n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , 
     n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , 
     n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , 
     n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , 
     n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , 
     n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , 
     n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , 
     n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , 
     n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , 
     n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , 
     n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , 
     n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , 
     n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , 
     n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , 
     n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , 
     n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , 
     n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , 
     n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , 
     n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , 
     n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , 
     n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , 
     n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , 
     n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , 
     n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , 
     n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , 
     n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , 
     n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , 
     n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , 
     n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , 
     n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , 
     n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , 
     n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , 
     n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , 
     n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , 
     n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , 
     n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , 
     n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , 
     n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , 
     n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , 
     n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , 
     n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , 
     n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , 
     n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , 
     n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , 
     n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , 
     n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , 
     n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , 
     n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , 
     n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , 
     n15081 , n15082 , n15083 ;
buf ( n2155 , n9744 );
buf ( n2160 , n11669 );
buf ( n2153 , n12927 );
buf ( n2156 , n13169 );
buf ( n2154 , n13618 );
buf ( n2158 , n14141 );
buf ( n2159 , n14428 );
buf ( n2151 , n14703 );
buf ( n2157 , n14855 );
buf ( n2152 , n15083 );
buf ( n4324 , n1942 );
buf ( n4325 , n855 );
buf ( n4326 , n1824 );
buf ( n4327 , n1443 );
buf ( n4328 , n1926 );
buf ( n4329 , n862 );
buf ( n4330 , n2088 );
buf ( n4331 , n150 );
buf ( n4332 , n1589 );
buf ( n4333 , n1827 );
buf ( n4334 , n617 );
buf ( n4335 , n478 );
buf ( n4336 , n1159 );
buf ( n4337 , n1856 );
buf ( n4338 , n1828 );
buf ( n4339 , n2015 );
buf ( n4340 , n2119 );
buf ( n4341 , n1660 );
buf ( n4342 , n2049 );
buf ( n4343 , n1934 );
buf ( n4344 , n808 );
buf ( n4345 , n405 );
buf ( n4346 , n446 );
buf ( n4347 , n504 );
buf ( n4348 , n335 );
buf ( n4349 , n462 );
buf ( n4350 , n1885 );
buf ( n4351 , n1102 );
buf ( n4352 , n540 );
buf ( n4353 , n299 );
buf ( n4354 , n1456 );
buf ( n4355 , n112 );
buf ( n4356 , n433 );
buf ( n4357 , n1171 );
buf ( n4358 , n1149 );
buf ( n4359 , n1860 );
buf ( n4360 , n53 );
buf ( n4361 , n1490 );
buf ( n4362 , n709 );
buf ( n4363 , n612 );
buf ( n4364 , n788 );
buf ( n4365 , n710 );
buf ( n4366 , n1773 );
buf ( n4367 , n1557 );
buf ( n4368 , n323 );
buf ( n4369 , n2130 );
buf ( n4370 , n332 );
buf ( n4371 , n2122 );
buf ( n4372 , n86 );
buf ( n4373 , n1536 );
buf ( n4374 , n261 );
buf ( n4375 , n960 );
buf ( n4376 , n85 );
buf ( n4377 , n2114 );
buf ( n4378 , n1616 );
buf ( n4379 , n1030 );
buf ( n4380 , n354 );
buf ( n4381 , n2012 );
buf ( n4382 , n977 );
buf ( n4383 , n1800 );
buf ( n4384 , n1894 );
buf ( n4385 , n1965 );
buf ( n4386 , n1432 );
buf ( n4387 , n1895 );
buf ( n4388 , n794 );
buf ( n4389 , n362 );
buf ( n4390 , n1685 );
buf ( n4391 , n1447 );
buf ( n4392 , n281 );
buf ( n4393 , n227 );
buf ( n4394 , n1903 );
buf ( n4395 , n1297 );
buf ( n4396 , n539 );
buf ( n4397 , n1199 );
buf ( n4398 , n1110 );
buf ( n4399 , n1591 );
buf ( n4400 , n1901 );
buf ( n4401 , n1809 );
buf ( n4402 , n1052 );
buf ( n4403 , n1700 );
buf ( n4404 , n1542 );
buf ( n4405 , n145 );
buf ( n4406 , n57 );
buf ( n4407 , n1155 );
buf ( n4408 , n853 );
buf ( n4409 , n1442 );
buf ( n4410 , n2070 );
buf ( n4411 , n1461 );
buf ( n4412 , n1971 );
buf ( n4413 , n1944 );
buf ( n4414 , n2065 );
buf ( n4415 , n886 );
buf ( n4416 , n1091 );
buf ( n4417 , n458 );
buf ( n4418 , n910 );
buf ( n4419 , n1884 );
buf ( n4420 , n1933 );
buf ( n4421 , n185 );
buf ( n4422 , n1917 );
buf ( n4423 , n1517 );
buf ( n4424 , n1981 );
buf ( n4425 , n1318 );
buf ( n4426 , n1814 );
buf ( n4427 , n743 );
buf ( n4428 , n270 );
buf ( n4429 , n682 );
buf ( n4430 , n2019 );
buf ( n4431 , n1729 );
buf ( n4432 , n334 );
buf ( n4433 , n1434 );
buf ( n4434 , n1332 );
buf ( n4435 , n1435 );
buf ( n4436 , n1397 );
buf ( n4437 , n1522 );
buf ( n4438 , n2043 );
buf ( n4439 , n1538 );
buf ( n4440 , n298 );
buf ( n4441 , n1646 );
buf ( n4442 , n1859 );
buf ( n4443 , n1280 );
buf ( n4444 , n1873 );
buf ( n4445 , n1380 );
buf ( n4446 , n83 );
buf ( n4447 , n938 );
buf ( n4448 , n649 );
buf ( n4449 , n1484 );
buf ( n4450 , n418 );
buf ( n4451 , n1419 );
buf ( n4452 , n651 );
buf ( n4453 , n94 );
buf ( n4454 , n292 );
buf ( n4455 , n211 );
buf ( n4456 , n833 );
buf ( n4457 , n1485 );
buf ( n4458 , n614 );
buf ( n4459 , n1483 );
buf ( n4460 , n1682 );
buf ( n4461 , n878 );
buf ( n4462 , n1277 );
buf ( n4463 , n1364 );
buf ( n4464 , n1546 );
buf ( n4465 , n1830 );
buf ( n4466 , n560 );
buf ( n4467 , n1357 );
buf ( n4468 , n1541 );
buf ( n4469 , n728 );
buf ( n4470 , n1991 );
buf ( n4471 , n570 );
buf ( n4472 , n1486 );
buf ( n4473 , n1999 );
buf ( n4474 , n454 );
buf ( n4475 , n267 );
buf ( n4476 , n2041 );
buf ( n4477 , n2031 );
buf ( n4478 , n180 );
buf ( n4479 , n136 );
buf ( n4480 , n857 );
buf ( n4481 , n719 );
buf ( n4482 , n983 );
buf ( n4483 , n2146 );
buf ( n4484 , n1068 );
buf ( n4485 , n1939 );
buf ( n4486 , n965 );
buf ( n4487 , n1197 );
buf ( n4488 , n1387 );
buf ( n4489 , n1709 );
buf ( n4490 , n1014 );
buf ( n4491 , n927 );
buf ( n4492 , n1531 );
buf ( n4493 , n301 );
buf ( n4494 , n222 );
buf ( n4495 , n1561 );
buf ( n4496 , n1931 );
buf ( n4497 , n242 );
buf ( n4498 , n1703 );
buf ( n4499 , n1889 );
buf ( n4500 , n732 );
buf ( n4501 , n1785 );
buf ( n4502 , n16 );
buf ( n4503 , n966 );
buf ( n4504 , n133 );
buf ( n4505 , n2028 );
buf ( n4506 , n946 );
buf ( n4507 , n375 );
buf ( n4508 , n8 );
buf ( n4509 , n1993 );
buf ( n4510 , n588 );
buf ( n4511 , n1691 );
buf ( n4512 , n1601 );
buf ( n4513 , n1044 );
buf ( n4514 , n703 );
buf ( n4515 , n825 );
buf ( n4516 , n976 );
buf ( n4517 , n1563 );
buf ( n4518 , n1831 );
buf ( n4519 , n403 );
buf ( n4520 , n643 );
buf ( n4521 , n579 );
buf ( n4522 , n1867 );
buf ( n4523 , n1912 );
buf ( n4524 , n998 );
buf ( n4525 , n1481 );
buf ( n4526 , n291 );
buf ( n4527 , n1697 );
buf ( n4528 , n1169 );
buf ( n4529 , n2080 );
buf ( n4530 , n1739 );
buf ( n4531 , n727 );
buf ( n4532 , n131 );
buf ( n4533 , n1238 );
buf ( n4534 , n1845 );
buf ( n4535 , n737 );
buf ( n4536 , n1244 );
buf ( n4537 , n1569 );
buf ( n4538 , n1018 );
buf ( n4539 , n1515 );
buf ( n4540 , n188 );
buf ( n4541 , n1115 );
buf ( n4542 , n2023 );
buf ( n4543 , n598 );
buf ( n4544 , n807 );
buf ( n4545 , n1241 );
buf ( n4546 , n1263 );
buf ( n4547 , n77 );
buf ( n4548 , n1207 );
buf ( n4549 , n1130 );
buf ( n4550 , n892 );
buf ( n4551 , n2045 );
buf ( n4552 , n979 );
buf ( n4553 , n169 );
buf ( n4554 , n1 );
buf ( n4555 , n1790 );
buf ( n4556 , n245 );
buf ( n4557 , n1202 );
buf ( n4558 , n1426 );
buf ( n4559 , n536 );
buf ( n4560 , n990 );
buf ( n4561 , n1161 );
buf ( n4562 , n722 );
buf ( n4563 , n30 );
buf ( n4564 , n2069 );
buf ( n4565 , n1943 );
buf ( n4566 , n609 );
buf ( n4567 , n1659 );
buf ( n4568 , n1356 );
buf ( n4569 , n1324 );
buf ( n4570 , n929 );
buf ( n4571 , n1510 );
buf ( n4572 , n1065 );
buf ( n4573 , n895 );
buf ( n4574 , n1609 );
buf ( n4575 , n1008 );
buf ( n4576 , n1424 );
buf ( n4577 , n82 );
buf ( n4578 , n618 );
buf ( n4579 , n1249 );
buf ( n4580 , n922 );
buf ( n4581 , n1182 );
buf ( n4582 , n681 );
buf ( n4583 , n184 );
buf ( n4584 , n528 );
buf ( n4585 , n535 );
buf ( n4586 , n1898 );
buf ( n4587 , n489 );
buf ( n4588 , n353 );
buf ( n4589 , n1163 );
buf ( n4590 , n899 );
buf ( n4591 , n1540 );
buf ( n4592 , n2058 );
buf ( n4593 , n129 );
buf ( n4594 , n1526 );
buf ( n4595 , n532 );
buf ( n4596 , n1454 );
buf ( n4597 , n974 );
buf ( n4598 , n1920 );
buf ( n4599 , n805 );
buf ( n4600 , n507 );
buf ( n4601 , n39 );
buf ( n4602 , n165 );
buf ( n4603 , n193 );
buf ( n4604 , n343 );
buf ( n4605 , n2135 );
buf ( n4606 , n1472 );
buf ( n4607 , n2044 );
buf ( n4608 , n600 );
buf ( n4609 , n2020 );
buf ( n4610 , n1690 );
buf ( n4611 , n199 );
buf ( n4612 , n1204 );
buf ( n4613 , n662 );
buf ( n4614 , n1096 );
buf ( n4615 , n360 );
buf ( n4616 , n881 );
buf ( n4617 , n395 );
buf ( n4618 , n1922 );
buf ( n4619 , n1964 );
buf ( n4620 , n1608 );
buf ( n4621 , n1452 );
buf ( n4622 , n1752 );
buf ( n4623 , n1640 );
buf ( n4624 , n1787 );
buf ( n4625 , n621 );
buf ( n4626 , n1172 );
buf ( n4627 , n1404 );
buf ( n4628 , n993 );
buf ( n4629 , n1594 );
buf ( n4630 , n1248 );
buf ( n4631 , n209 );
buf ( n4632 , n1467 );
buf ( n4633 , n501 );
buf ( n4634 , n1832 );
buf ( n4635 , n1675 );
buf ( n4636 , n2016 );
buf ( n4637 , n2120 );
buf ( n4638 , n1529 );
buf ( n4639 , n1413 );
buf ( n4640 , n1862 );
buf ( n4641 , n386 );
buf ( n4642 , n1665 );
buf ( n4643 , n970 );
buf ( n4644 , n1041 );
buf ( n4645 , n1039 );
buf ( n4646 , n942 );
buf ( n4647 , n823 );
buf ( n4648 , n260 );
buf ( n4649 , n711 );
buf ( n4650 , n1144 );
buf ( n4651 , n1004 );
buf ( n4652 , n764 );
buf ( n4653 , n293 );
buf ( n4654 , n1812 );
buf ( n4655 , n288 );
buf ( n4656 , n918 );
buf ( n4657 , n11 );
buf ( n4658 , n1639 );
buf ( n4659 , n1308 );
buf ( n4660 , n356 );
buf ( n4661 , n198 );
buf ( n4662 , n747 );
buf ( n4663 , n48 );
buf ( n4664 , n376 );
buf ( n4665 , n465 );
buf ( n4666 , n445 );
buf ( n4667 , n1469 );
buf ( n4668 , n1389 );
buf ( n4669 , n1525 );
buf ( n4670 , n1181 );
buf ( n4671 , n510 );
buf ( n4672 , n880 );
buf ( n4673 , n1474 );
buf ( n4674 , n278 );
buf ( n4675 , n1829 );
buf ( n4676 , n1326 );
buf ( n4677 , n1506 );
buf ( n4678 , n2053 );
buf ( n4679 , n1875 );
buf ( n4680 , n443 );
buf ( n4681 , n940 );
buf ( n4682 , n246 );
buf ( n4683 , n240 );
buf ( n4684 , n1037 );
buf ( n4685 , n144 );
buf ( n4686 , n992 );
buf ( n4687 , n296 );
buf ( n4688 , n42 );
buf ( n4689 , n1650 );
buf ( n4690 , n1187 );
buf ( n4691 , n1183 );
buf ( n4692 , n306 );
buf ( n4693 , n2017 );
buf ( n4694 , n1232 );
buf ( n4695 , n453 );
buf ( n4696 , n1710 );
buf ( n4697 , n1198 );
buf ( n4698 , n1794 );
buf ( n4699 , n1567 );
buf ( n4700 , n64 );
buf ( n4701 , n1251 );
buf ( n4702 , n1261 );
buf ( n4703 , n1027 );
buf ( n4704 , n784 );
buf ( n4705 , n388 );
buf ( n4706 , n754 );
buf ( n4707 , n619 );
buf ( n4708 , n2022 );
buf ( n4709 , n801 );
buf ( n4710 , n1975 );
buf ( n4711 , n1177 );
buf ( n4712 , n2084 );
buf ( n4713 , n1491 );
buf ( n4714 , n900 );
buf ( n4715 , n790 );
buf ( n4716 , n1784 );
buf ( n4717 , n1861 );
buf ( n4718 , n2033 );
buf ( n4719 , n2047 );
buf ( n4720 , n1976 );
buf ( n4721 , n533 );
buf ( n4722 , n1103 );
buf ( n4723 , n1393 );
buf ( n4724 , n1410 );
buf ( n4725 , n2060 );
buf ( n4726 , n1225 );
buf ( n4727 , n1841 );
buf ( n4728 , n1222 );
buf ( n4729 , n1322 );
buf ( n4730 , n1825 );
buf ( n4731 , n487 );
buf ( n4732 , n497 );
buf ( n4733 , n836 );
buf ( n4734 , n1977 );
buf ( n4735 , n1568 );
buf ( n4736 , n1153 );
buf ( n4737 , n1124 );
buf ( n4738 , n2112 );
buf ( n4739 , n2026 );
buf ( n4740 , n714 );
buf ( n4741 , n5 );
buf ( n4742 , n1108 );
buf ( n4743 , n1267 );
buf ( n4744 , n2089 );
buf ( n4745 , n68 );
buf ( n4746 , n2004 );
buf ( n4747 , n1087 );
buf ( n4748 , n997 );
buf ( n4749 , n21 );
buf ( n4750 , n680 );
buf ( n4751 , n1116 );
buf ( n4752 , n340 );
buf ( n4753 , n1822 );
buf ( n4754 , n1274 );
buf ( n4755 , n771 );
buf ( n4756 , n2024 );
buf ( n4757 , n2066 );
buf ( n4758 , n1462 );
buf ( n4759 , n1985 );
buf ( n4760 , n913 );
buf ( n4761 , n787 );
buf ( n4762 , n1978 );
buf ( n4763 , n1123 );
buf ( n4764 , n415 );
buf ( n4765 , n1063 );
buf ( n4766 , n995 );
buf ( n4767 , n370 );
buf ( n4768 , n544 );
buf ( n4769 , n1119 );
buf ( n4770 , n1492 );
buf ( n4771 , n636 );
buf ( n4772 , n172 );
buf ( n4773 , n1450 );
buf ( n4774 , n26 );
buf ( n4775 , n2123 );
buf ( n4776 , n18 );
buf ( n4777 , n838 );
buf ( n4778 , n146 );
buf ( n4779 , n123 );
buf ( n4780 , n1910 );
buf ( n4781 , n441 );
buf ( n4782 , n700 );
buf ( n4783 , n194 );
buf ( n4784 , n1127 );
buf ( n4785 , n872 );
buf ( n4786 , n1239 );
buf ( n4787 , n848 );
buf ( n4788 , n765 );
buf ( n4789 , n1580 );
buf ( n4790 , n751 );
buf ( n4791 , n1560 );
buf ( n4792 , n920 );
buf ( n4793 , n318 );
buf ( n4794 , n1819 );
buf ( n4795 , n206 );
buf ( n4796 , n1145 );
buf ( n4797 , n1562 );
buf ( n4798 , n1651 );
buf ( n4799 , n2064 );
buf ( n4800 , n1464 );
buf ( n4801 , n1367 );
buf ( n4802 , n1950 );
buf ( n4803 , n1994 );
buf ( n4804 , n1487 );
buf ( n4805 , n1081 );
buf ( n4806 , n1575 );
buf ( n4807 , n2082 );
buf ( n4808 , n338 );
buf ( n4809 , n592 );
buf ( n4810 , n961 );
buf ( n4811 , n546 );
buf ( n4812 , n1801 );
buf ( n4813 , n119 );
buf ( n4814 , n1283 );
buf ( n4815 , n1743 );
buf ( n4816 , n1792 );
buf ( n4817 , n432 );
buf ( n4818 , n1770 );
buf ( n4819 , n821 );
buf ( n4820 , n1547 );
buf ( n4821 , n2042 );
buf ( n4822 , n1293 );
buf ( n4823 , n557 );
buf ( n4824 , n1657 );
buf ( n4825 , n173 );
buf ( n4826 , n1047 );
buf ( n4827 , n1771 );
buf ( n4828 , n156 );
buf ( n4829 , n1558 );
buf ( n4830 , n1803 );
buf ( n4831 , n1602 );
buf ( n4832 , n740 );
buf ( n4833 , n1804 );
buf ( n4834 , n191 );
buf ( n4835 , n1001 );
buf ( n4836 , n605 );
buf ( n4837 , n777 );
buf ( n4838 , n1275 );
buf ( n4839 , n226 );
buf ( n4840 , n1671 );
buf ( n4841 , n1628 );
buf ( n4842 , n803 );
buf ( n4843 , n502 );
buf ( n4844 , n361 );
buf ( n4845 , n1365 );
buf ( n4846 , n516 );
buf ( n4847 , n111 );
buf ( n4848 , n475 );
buf ( n4849 , n98 );
buf ( n4850 , n2054 );
buf ( n4851 , n1963 );
buf ( n4852 , n1019 );
buf ( n4853 , n843 );
buf ( n4854 , n1016 );
buf ( n4855 , n1125 );
buf ( n4856 , n1706 );
buf ( n4857 , n574 );
buf ( n4858 , n2098 );
buf ( n4859 , n1255 );
buf ( n4860 , n2108 );
buf ( n4861 , n2046 );
buf ( n4862 , n873 );
buf ( n4863 , n639 );
buf ( n4864 , n1677 );
buf ( n4865 , n1061 );
buf ( n4866 , n964 );
buf ( n4867 , n1220 );
buf ( n4868 , n904 );
buf ( n4869 , n108 );
buf ( n4870 , n683 );
buf ( n4871 , n554 );
buf ( n4872 , n1478 );
buf ( n4873 , n394 );
buf ( n4874 , n1708 );
buf ( n4875 , n1618 );
buf ( n4876 , n1279 );
buf ( n4877 , n328 );
buf ( n4878 , n1042 );
buf ( n4879 , n1699 );
buf ( n4880 , n1190 );
buf ( n4881 , n40 );
buf ( n4882 , n2150 );
buf ( n4883 , n1023 );
buf ( n4884 , n371 );
buf ( n4885 , n2145 );
buf ( n4886 , n1216 );
buf ( n4887 , n1635 );
buf ( n4888 , n1218 );
buf ( n4889 , n551 );
buf ( n4890 , n1806 );
buf ( n4891 , n320 );
buf ( n4892 , n494 );
buf ( n4893 , n827 );
buf ( n4894 , n1865 );
buf ( n4895 , n1139 );
buf ( n4896 , n23 );
buf ( n4897 , n1412 );
buf ( n4898 , n324 );
buf ( n4899 , n495 );
buf ( n4900 , n778 );
buf ( n4901 , n792 );
buf ( n4902 , n654 );
buf ( n4903 , n312 );
buf ( n4904 , n383 );
buf ( n4905 , n1347 );
buf ( n4906 , n520 );
buf ( n4907 , n816 );
buf ( n4908 , n1749 );
buf ( n4909 , n20 );
buf ( n4910 , n103 );
buf ( n4911 , n263 );
buf ( n4912 , n1128 );
buf ( n4913 , n2009 );
buf ( n4914 , n1284 );
buf ( n4915 , n891 );
buf ( n4916 , n1737 );
buf ( n4917 , n679 );
buf ( n4918 , n1282 );
buf ( n4919 , n425 );
buf ( n4920 , n1644 );
buf ( n4921 , n1610 );
buf ( n4922 , n33 );
buf ( n4923 , n2137 );
buf ( n4924 , n1906 );
buf ( n4925 , n1196 );
buf ( n4926 , n1619 );
buf ( n4927 , n1430 );
buf ( n4928 , n1213 );
buf ( n4929 , n170 );
buf ( n4930 , n1031 );
buf ( n4931 , n686 );
buf ( n4932 , n234 );
buf ( n4933 , n480 );
buf ( n4934 , n1359 );
buf ( n4935 , n1681 );
buf ( n4936 , n1720 );
buf ( n4937 , n9 );
buf ( n4938 , n1571 );
buf ( n4939 , n943 );
buf ( n4940 , n645 );
buf ( n4941 , n1329 );
buf ( n4942 , n1390 );
buf ( n4943 , n1496 );
buf ( n4944 , n907 );
buf ( n4945 , n1338 );
buf ( n4946 , n933 );
buf ( n4947 , n1111 );
buf ( n4948 , n810 );
buf ( n4949 , n569 );
buf ( n4950 , n517 );
buf ( n4951 , n916 );
buf ( n4952 , n1998 );
buf ( n4953 , n1319 );
buf ( n4954 , n1961 );
buf ( n4955 , n587 );
buf ( n4956 , n1438 );
buf ( n4957 , n1925 );
buf ( n4958 , n715 );
buf ( n4959 , n1764 );
buf ( n4960 , n1033 );
buf ( n4961 , n1995 );
buf ( n4962 , n461 );
buf ( n4963 , n1075 );
buf ( n4964 , n661 );
buf ( n4965 , n344 );
buf ( n4966 , n2149 );
buf ( n4967 , n1882 );
buf ( n4968 , n1872 );
buf ( n4969 , n2013 );
buf ( n4970 , n1291 );
buf ( n4971 , n1695 );
buf ( n4972 , n746 );
buf ( n4973 , n2105 );
buf ( n4974 , n1757 );
buf ( n4975 , n748 );
buf ( n4976 , n2115 );
buf ( n4977 , n1339 );
buf ( n4978 , n1721 );
buf ( n4979 , n841 );
buf ( n4980 , n1946 );
buf ( n4981 , n1970 );
buf ( n4982 , n1897 );
buf ( n4983 , n444 );
buf ( n4984 , n92 );
buf ( n4985 , n266 );
buf ( n4986 , n834 );
buf ( n4987 , n814 );
buf ( n4988 , n1024 );
buf ( n4989 , n1473 );
buf ( n4990 , n1226 );
buf ( n4991 , n1554 );
buf ( n4992 , n628 );
buf ( n4993 , n1133 );
buf ( n4994 , n471 );
buf ( n4995 , n1323 );
buf ( n4996 , n1109 );
buf ( n4997 , n317 );
buf ( n4998 , n730 );
buf ( n4999 , n236 );
buf ( n5000 , n753 );
buf ( n5001 , n1870 );
buf ( n5002 , n513 );
buf ( n5003 , n1751 );
buf ( n5004 , n1394 );
buf ( n5005 , n158 );
buf ( n5006 , n249 );
buf ( n5007 , n248 );
buf ( n5008 , n572 );
buf ( n5009 , n190 );
buf ( n5010 , n421 );
buf ( n5011 , n1600 );
buf ( n5012 , n1564 );
buf ( n5013 , n247 );
buf ( n5014 , n1361 );
buf ( n5015 , n1871 );
buf ( n5016 , n1100 );
buf ( n5017 , n956 );
buf ( n5018 , n2079 );
buf ( n5019 , n1195 );
buf ( n5020 , n1980 );
buf ( n5021 , n692 );
buf ( n5022 , n1876 );
buf ( n5023 , n382 );
buf ( n5024 , n1437 );
buf ( n5025 , n869 );
buf ( n5026 , n1919 );
buf ( n5027 , n1632 );
buf ( n5028 , n45 );
buf ( n5029 , n2068 );
buf ( n5030 , n1669 );
buf ( n5031 , n391 );
buf ( n5032 , n1223 );
buf ( n5033 , n1736 );
buf ( n5034 , n349 );
buf ( n5035 , n476 );
buf ( n5036 , n1893 );
buf ( n5037 , n1193 );
buf ( n5038 , n1949 );
buf ( n5039 , n2067 );
buf ( n5040 , n731 );
buf ( n5041 , n315 );
buf ( n5042 , n1234 );
buf ( n5043 , n1070 );
buf ( n5044 , n1458 );
buf ( n5045 , n1505 );
buf ( n5046 , n1034 );
buf ( n5047 , n1900 );
buf ( n5048 , n2093 );
buf ( n5049 , n739 );
buf ( n5050 , n538 );
buf ( n5051 , n19 );
buf ( n5052 , n1664 );
buf ( n5053 , n758 );
buf ( n5054 , n1088 );
buf ( n5055 , n287 );
buf ( n5056 , n789 );
buf ( n5057 , n34 );
buf ( n5058 , n791 );
buf ( n5059 , n717 );
buf ( n5060 , n1840 );
buf ( n5061 , n697 );
buf ( n5062 , n1170 );
buf ( n5063 , n1537 );
buf ( n5064 , n1683 );
buf ( n5065 , n999 );
buf ( n5066 , n367 );
buf ( n5067 , n393 );
buf ( n5068 , n1559 );
buf ( n5069 , n1599 );
buf ( n5070 , n1342 );
buf ( n5071 , n2078 );
buf ( n5072 , n1050 );
buf ( n5073 , n243 );
buf ( n5074 , n2144 );
buf ( n5075 , n1266 );
buf ( n5076 , n1298 );
buf ( n5077 , n1301 );
buf ( n5078 , n1962 );
buf ( n5079 , n812 );
buf ( n5080 , n583 );
buf ( n5081 , n27 );
buf ( n5082 , n87 );
buf ( n5083 , n1415 );
buf ( n5084 , n201 );
buf ( n5085 , n1497 );
buf ( n5086 , n1808 );
buf ( n5087 , n1570 );
buf ( n5088 , n327 );
buf ( n5089 , n2086 );
buf ( n5090 , n1448 );
buf ( n5091 , n414 );
buf ( n5092 , n1320 );
buf ( n5093 , n775 );
buf ( n5094 , n760 );
buf ( n5095 , n1307 );
buf ( n5096 , n2036 );
buf ( n5097 , n404 );
buf ( n5098 , n1519 );
buf ( n5099 , n254 );
buf ( n5100 , n1548 );
buf ( n5101 , n647 );
buf ( n5102 , n1908 );
buf ( n5103 , n1979 );
buf ( n5104 , n1890 );
buf ( n5105 , n1136 );
buf ( n5106 , n276 );
buf ( n5107 , n67 );
buf ( n5108 , n988 );
buf ( n5109 , n1603 );
buf ( n5110 , n274 );
buf ( n5111 , n231 );
buf ( n5112 , n625 );
buf ( n5113 , n366 );
buf ( n5114 , n413 );
buf ( n5115 , n428 );
buf ( n5116 , n381 );
buf ( n5117 , n1230 );
buf ( n5118 , n1772 );
buf ( n5119 , n179 );
buf ( n5120 , n978 );
buf ( n5121 , n147 );
buf ( n5122 , n1987 );
buf ( n5123 , n177 );
buf ( n5124 , n1252 );
buf ( n5125 , n1309 );
buf ( n5126 , n1673 );
buf ( n5127 , n1160 );
buf ( n5128 , n914 );
buf ( n5129 , n811 );
buf ( n5130 , n498 );
buf ( n5131 , n725 );
buf ( n5132 , n1625 );
buf ( n5133 , n79 );
buf ( n5134 , n2103 );
buf ( n5135 , n503 );
buf ( n5136 , n1140 );
buf ( n5137 , n1762 );
buf ( n5138 , n1362 );
buf ( n5139 , n842 );
buf ( n5140 , n1643 );
buf ( n5141 , n1045 );
buf ( n5142 , n809 );
buf ( n5143 , n1718 );
buf ( n5144 , n303 );
buf ( n5145 , n2096 );
buf ( n5146 , n1730 );
buf ( n5147 , n1530 );
buf ( n5148 , n157 );
buf ( n5149 , n32 );
buf ( n5150 , n1494 );
buf ( n5151 , n1208 );
buf ( n5152 , n1094 );
buf ( n5153 , n580 );
buf ( n5154 , n2021 );
buf ( n5155 , n599 );
buf ( n5156 , n1314 );
buf ( n5157 , n1224 );
buf ( n5158 , n1378 );
buf ( n5159 , n1959 );
buf ( n5160 , n212 );
buf ( n5161 , n1117 );
buf ( n5162 , n1966 );
buf ( n5163 , n930 );
buf ( n5164 , n1731 );
buf ( n5165 , n1214 );
buf ( n5166 , n59 );
buf ( n5167 , n275 );
buf ( n5168 , n901 );
buf ( n5169 , n694 );
buf ( n5170 , n1395 );
buf ( n5171 , n529 );
buf ( n5172 , n1521 );
buf ( n5173 , n543 );
buf ( n5174 , n1465 );
buf ( n5175 , n1436 );
buf ( n5176 , n219 );
buf ( n5177 , n396 );
buf ( n5178 , n1194 );
buf ( n5179 , n104 );
buf ( n5180 , n1015 );
buf ( n5181 , n1092 );
buf ( n5182 , n1089 );
buf ( n5183 , n1909 );
buf ( n5184 , n481 );
buf ( n5185 , n925 );
buf ( n5186 , n1672 );
buf ( n5187 , n38 );
buf ( n5188 , n646 );
buf ( n5189 , n1622 );
buf ( n5190 , n490 );
buf ( n5191 , n250 );
buf ( n5192 , n436 );
buf ( n5193 , n1209 );
buf ( n5194 , n1414 );
buf ( n5195 , n218 );
buf ( n5196 , n1341 );
buf ( n5197 , n400 );
buf ( n5198 , n594 );
buf ( n5199 , n1340 );
buf ( n5200 , n1440 );
buf ( n5201 , n795 );
buf ( n5202 , n1688 );
buf ( n5203 , n813 );
buf ( n5204 , n768 );
buf ( n5205 , n1837 );
buf ( n5206 , n4 );
buf ( n5207 , n1250 );
buf ( n5208 , n449 );
buf ( n5209 , n1888 );
buf ( n5210 , n74 );
buf ( n5211 , n106 );
buf ( n5212 , n534 );
buf ( n5213 , n1711 );
buf ( n5214 , n500 );
buf ( n5215 , n1881 );
buf ( n5216 , n766 );
buf ( n5217 , n66 );
buf ( n5218 , n849 );
buf ( n5219 , n470 );
buf ( n5220 , n620 );
buf ( n5221 , n1797 );
buf ( n5222 , n460 );
buf ( n5223 , n216 );
buf ( n5224 , n1642 );
buf ( n5225 , n1099 );
buf ( n5226 , n1958 );
buf ( n5227 , n1523 );
buf ( n5228 , n410 );
buf ( n5229 , n1349 );
buf ( n5230 , n1725 );
buf ( n5231 , n1372 );
buf ( n5232 , n37 );
buf ( n5233 , n1620 );
buf ( n5234 , n888 );
buf ( n5235 , n1057 );
buf ( n5236 , n352 );
buf ( n5237 , n1754 );
buf ( n5238 , n1074 );
buf ( n5239 , n931 );
buf ( n5240 , n1168 );
buf ( n5241 , n1383 );
buf ( n5242 , n2050 );
buf ( n5243 , n1376 );
buf ( n5244 , n1914 );
buf ( n5245 , n62 );
buf ( n5246 , n2006 );
buf ( n5247 , n2148 );
buf ( n5248 , n2107 );
buf ( n5249 , n782 );
buf ( n5250 , n1276 );
buf ( n5251 , n1180 );
buf ( n5252 , n2 );
buf ( n5253 , n148 );
buf ( n5254 , n1686 );
buf ( n5255 , n952 );
buf ( n5256 , n93 );
buf ( n5257 , n1887 );
buf ( n5258 , n1420 );
buf ( n5259 , n1913 );
buf ( n5260 , n512 );
buf ( n5261 , n2027 );
buf ( n5262 , n1955 );
buf ( n5263 , n402 );
buf ( n5264 , n596 );
buf ( n5265 , n440 );
buf ( n5266 , n1641 );
buf ( n5267 , n1405 );
buf ( n5268 , n2038 );
buf ( n5269 , n65 );
buf ( n5270 , n1713 );
buf ( n5271 , n829 );
buf ( n5272 , n153 );
buf ( n5273 , n1624 );
buf ( n5274 , n1617 );
buf ( n5275 , n898 );
buf ( n5276 , n934 );
buf ( n5277 , n355 );
buf ( n5278 , n1316 );
buf ( n5279 , n1185 );
buf ( n5280 , n1431 );
buf ( n5281 , n1745 );
buf ( n5282 , n1680 );
buf ( n5283 , n1085 );
buf ( n5284 , n844 );
buf ( n5285 , n35 );
buf ( n5286 , n562 );
buf ( n5287 , n161 );
buf ( n5288 , n947 );
buf ( n5289 , n409 );
buf ( n5290 , n1585 );
buf ( n5291 , n1868 );
buf ( n5292 , n1007 );
buf ( n5293 , n2000 );
buf ( n5294 , n1891 );
buf ( n5295 , n1444 );
buf ( n5296 , n1779 );
buf ( n5297 , n949 );
buf ( n5298 , n1247 );
buf ( n5299 , n1636 );
buf ( n5300 , n130 );
buf ( n5301 , n1941 );
buf ( n5302 , n2087 );
buf ( n5303 , n139 );
buf ( n5304 , n1049 );
buf ( n5305 , n1866 );
buf ( n5306 , n2052 );
buf ( n5307 , n2034 );
buf ( n5308 , n912 );
buf ( n5309 , n1401 );
buf ( n5310 , n1974 );
buf ( n5311 , n1344 );
buf ( n5312 , n744 );
buf ( n5313 , n91 );
buf ( n5314 , n987 );
buf ( n5315 , n819 );
buf ( n5316 , n644 );
buf ( n5317 , n1086 );
buf ( n5318 , n58 );
buf ( n5319 , n1501 );
buf ( n5320 , n1579 );
buf ( n5321 , n1005 );
buf ( n5322 , n839 );
buf ( n5323 , n678 );
buf ( n5324 , n1131 );
buf ( n5325 , n1503 );
buf ( n5326 , n1511 );
buf ( n5327 , n745 );
buf ( n5328 , n1305 );
buf ( n5329 , n214 );
buf ( n5330 , n73 );
buf ( n5331 , n951 );
buf ( n5332 , n1802 );
buf ( n5333 , n1791 );
buf ( n5334 , n1231 );
buf ( n5335 , n1482 );
buf ( n5336 , n606 );
buf ( n5337 , n752 );
buf ( n5338 , n75 );
buf ( n5339 , n1896 );
buf ( n5340 , n932 );
buf ( n5341 , n1457 );
buf ( n5342 , n1883 );
buf ( n5343 , n1631 );
buf ( n5344 , n1952 );
buf ( n5345 , n558 );
buf ( n5346 , n542 );
buf ( n5347 , n1733 );
buf ( n5348 , n1928 );
buf ( n5349 , n2048 );
buf ( n5350 , n295 );
buf ( n5351 , n601 );
buf ( n5352 , n524 );
buf ( n5353 , n1674 );
buf ( n5354 , n1377 );
buf ( n5355 , n657 );
buf ( n5356 , n398 );
buf ( n5357 , n2029 );
buf ( n5358 , n1878 );
buf ( n5359 , n1783 );
buf ( n5360 , n1142 );
buf ( n5361 , n1629 );
buf ( n5362 , n101 );
buf ( n5363 , n1189 );
buf ( n5364 , n508 );
buf ( n5365 , n1705 );
buf ( n5366 , n603 );
buf ( n5367 , n511 );
buf ( n5368 , n1158 );
buf ( n5369 , n364 );
buf ( n5370 , n10 );
buf ( n5371 , n1353 );
buf ( n5372 , n183 );
buf ( n5373 , n1833 );
buf ( n5374 , n716 );
buf ( n5375 , n1598 );
buf ( n5376 , n1902 );
buf ( n5377 , n1229 );
buf ( n5378 , n2090 );
buf ( n5379 , n2104 );
buf ( n5380 , n56 );
buf ( n5381 , n1707 );
buf ( n5382 , n182 );
buf ( n5383 , n2072 );
buf ( n5384 , n1360 );
buf ( n5385 , n163 );
buf ( n5386 , n1938 );
buf ( n5387 , n1370 );
buf ( n5388 , n1411 );
buf ( n5389 , n684 );
buf ( n5390 , n426 );
buf ( n5391 , n688 );
buf ( n5392 , n1043 );
buf ( n5393 , n1543 );
buf ( n5394 , n879 );
buf ( n5395 , n1849 );
buf ( n5396 , n164 );
buf ( n5397 , n1732 );
buf ( n5398 , n707 );
buf ( n5399 , n368 );
buf ( n5400 , n485 );
buf ( n5401 , n615 );
buf ( n5402 , n826 );
buf ( n5403 , n1984 );
buf ( n5404 , n695 );
buf ( n5405 , n1805 );
buf ( n5406 , n472 );
buf ( n5407 , n1026 );
buf ( n5408 , n369 );
buf ( n5409 , n2055 );
buf ( n5410 , n804 );
buf ( n5411 , n447 );
buf ( n5412 , n171 );
buf ( n5413 , n1850 );
buf ( n5414 , n1152 );
buf ( n5415 , n509 );
buf ( n5416 , n235 );
buf ( n5417 , n1135 );
buf ( n5418 , n733 );
buf ( n5419 , n972 );
buf ( n5420 , n1054 );
buf ( n5421 , n1532 );
buf ( n5422 , n1549 );
buf ( n5423 , n357 );
buf ( n5424 , n223 );
buf ( n5425 , n982 );
buf ( n5426 , n141 );
buf ( n5427 , n780 );
buf ( n5428 , n134 );
buf ( n5429 , n866 );
buf ( n5430 , n7 );
buf ( n5431 , n1003 );
buf ( n5432 , n1287 );
buf ( n5433 , n1466 );
buf ( n5434 , n167 );
buf ( n5435 , n220 );
buf ( n5436 , n1930 );
buf ( n5437 , n187 );
buf ( n5438 , n1429 );
buf ( n5439 , n802 );
buf ( n5440 , n593 );
buf ( n5441 , n767 );
buf ( n5442 , n991 );
buf ( n5443 , n1072 );
buf ( n5444 , n670 );
buf ( n5445 , n407 );
buf ( n5446 , n1290 );
buf ( n5447 , n1191 );
buf ( n5448 , n530 );
buf ( n5449 , n984 );
buf ( n5450 , n181 );
buf ( n5451 , n1687 );
buf ( n5452 , n15 );
buf ( n5453 , n877 );
buf ( n5454 , n464 );
buf ( n5455 , n416 );
buf ( n5456 , n176 );
buf ( n5457 , n1755 );
buf ( n5458 , n1826 );
buf ( n5459 , n720 );
buf ( n5460 , n996 );
buf ( n5461 , n785 );
buf ( n5462 , n310 );
buf ( n5463 , n380 );
buf ( n5464 , n708 );
buf ( n5465 , n1539 );
buf ( n5466 , n1126 );
buf ( n5467 , n1281 );
buf ( n5468 , n1192 );
buf ( n5469 , n1623 );
buf ( n5470 , n1406 );
buf ( n5471 , n0 );
buf ( n5472 , n2085 );
buf ( n5473 , n384 );
buf ( n5474 , n1311 );
buf ( n5475 , n1165 );
buf ( n5476 , n84 );
buf ( n5477 , n691 );
buf ( n5478 , n2138 );
buf ( n5479 , n669 );
buf ( n5480 , n521 );
buf ( n5481 , n1502 );
buf ( n5482 , n1038 );
buf ( n5483 , n1653 );
buf ( n5484 , n2014 );
buf ( n5485 , n392 );
buf ( n5486 , n1325 );
buf ( n5487 , n624 );
buf ( n5488 , n1178 );
buf ( n5489 , n1670 );
buf ( n5490 , n1455 );
buf ( n5491 , n1905 );
buf ( n5492 , n257 );
buf ( n5493 , n1392 );
buf ( n5494 , n518 );
buf ( n5495 , n1336 );
buf ( n5496 , n1471 );
buf ( n5497 , n1271 );
buf ( n5498 , n638 );
buf ( n5499 , n1334 );
buf ( n5500 , n1060 );
buf ( n5501 , n2095 );
buf ( n5502 , n980 );
buf ( n5503 , n174 );
buf ( n5504 , n107 );
buf ( n5505 , n847 );
buf ( n5506 , n1652 );
buf ( n5507 , n363 );
buf ( n5508 , n1017 );
buf ( n5509 , n2109 );
buf ( n5510 , n224 );
buf ( n5511 , n1141 );
buf ( n5512 , n1937 );
buf ( n5513 , n665 );
buf ( n5514 , n773 );
buf ( n5515 , n1303 );
buf ( n5516 , n1221 );
buf ( n5517 , n1516 );
buf ( n5518 , n1460 );
buf ( n5519 , n499 );
buf ( n5520 , n577 );
buf ( n5521 , n824 );
buf ( n5522 , n749 );
buf ( n5523 , n1815 );
buf ( n5524 , n1838 );
buf ( n5525 , n527 );
buf ( n5526 , n884 );
buf ( n5527 , n629 );
buf ( n5528 , n1294 );
buf ( n5529 , n1062 );
buf ( n5530 , n840 );
buf ( n5531 , n1106 );
buf ( n5532 , n1138 );
buf ( n5533 , n1527 );
buf ( n5534 , n309 );
buf ( n5535 , n1716 );
buf ( n5536 , n573 );
buf ( n5537 , n1385 );
buf ( n5538 , n1449 );
buf ( n5539 , n2083 );
buf ( n5540 , n1407 );
buf ( n5541 , n262 );
buf ( n5542 , n294 );
buf ( n5543 , n1777 );
buf ( n5544 , n1445 );
buf ( n5545 , n438 );
buf ( n5546 , n1647 );
buf ( n5547 , n1493 );
buf ( n5548 , n723 );
buf ( n5549 , n1753 );
buf ( n5550 , n1596 );
buf ( n5551 , n1799 );
buf ( n5552 , n2001 );
buf ( n5553 , n1315 );
buf ( n5554 , n1658 );
buf ( n5555 , n1433 );
buf ( n5556 , n2074 );
buf ( n5557 , n1747 );
buf ( n5558 , n2076 );
buf ( n5559 , n1992 );
buf ( n5560 , n2091 );
buf ( n5561 , n143 );
buf ( n5562 , n874 );
buf ( n5563 , n12 );
buf ( n5564 , n47 );
buf ( n5565 , n1036 );
buf ( n5566 , n1702 );
buf ( n5567 , n1083 );
buf ( n5568 , n491 );
buf ( n5569 , n431 );
buf ( n5570 , n346 );
buf ( n5571 , n1176 );
buf ( n5572 , n1488 );
buf ( n5573 , n1327 );
buf ( n5574 , n365 );
buf ( n5575 , n50 );
buf ( n5576 , n373 );
buf ( n5577 , n893 );
buf ( n5578 , n863 );
buf ( n5579 , n1836 );
buf ( n5580 , n200 );
buf ( n5581 , n1374 );
buf ( n5582 , n1246 );
buf ( n5583 , n1508 );
buf ( n5584 , n687 );
buf ( n5585 , n944 );
buf ( n5586 , n1907 );
buf ( n5587 , n1154 );
buf ( n5588 , n113 );
buf ( n5589 , n71 );
buf ( n5590 , n1656 );
buf ( n5591 , n280 );
buf ( n5592 , n1388 );
buf ( n5593 , n186 );
buf ( n5594 , n1173 );
buf ( n5595 , n2129 );
buf ( n5596 , n2051 );
buf ( n5597 , n1032 );
buf ( n5598 , n154 );
buf ( n5599 , n655 );
buf ( n5600 , n305 );
buf ( n5601 , n330 );
buf ( n5602 , n671 );
buf ( n5603 , n1375 );
buf ( n5604 , n466 );
buf ( n5605 , n1079 );
buf ( n5606 , n1048 );
buf ( n5607 , n452 );
buf ( n5608 , n779 );
buf ( n5609 , n1556 );
buf ( n5610 , n1951 );
buf ( n5611 , n781 );
buf ( n5612 , n798 );
buf ( n5613 , n889 );
buf ( n5614 , n1615 );
buf ( n5615 , n955 );
buf ( n5616 , n22 );
buf ( n5617 , n2037 );
buf ( n5618 , n1863 );
buf ( n5619 , n1550 );
buf ( n5620 , n1046 );
buf ( n5621 , n762 );
buf ( n5622 , n1839 );
buf ( n5623 , n985 );
buf ( n5624 , n2116 );
buf ( n5625 , n883 );
buf ( n5626 , n1258 );
buf ( n5627 , n835 );
buf ( n5628 , n1107 );
buf ( n5629 , n140 );
buf ( n5630 , n3 );
buf ( n5631 , n1584 );
buf ( n5632 , n656 );
buf ( n5633 , n556 );
buf ( n5634 , n1855 );
buf ( n5635 , n459 );
buf ( n5636 , n658 );
buf ( n5637 , n1260 );
buf ( n5638 , n1954 );
buf ( n5639 , n1021 );
buf ( n5640 , n450 );
buf ( n5641 , n1535 );
buf ( n5642 , n60 );
buf ( n5643 , n1760 );
buf ( n5644 , n676 );
buf ( n5645 , n1114 );
buf ( n5646 , n448 );
buf ( n5647 , n522 );
buf ( n5648 , n1264 );
buf ( n5649 , n253 );
buf ( n5650 , n1844 );
buf ( n5651 , n1157 );
buf ( n5652 , n1425 );
buf ( n5653 , n1678 );
buf ( n5654 , n1210 );
buf ( n5655 , n1398 );
buf ( n5656 , n850 );
buf ( n5657 , n1583 );
buf ( n5658 , n2101 );
buf ( n5659 , n1935 );
buf ( n5660 , n1381 );
buf ( n5661 , n1428 );
buf ( n5662 , n911 );
buf ( n5663 , n2134 );
buf ( n5664 , n868 );
buf ( n5665 , n876 );
buf ( n5666 , n228 );
buf ( n5667 , n1911 );
buf ( n5668 , n763 );
buf ( n5669 , n1273 );
buf ( n5670 , n1028 );
buf ( n5671 , n1071 );
buf ( n5672 , n523 );
buf ( n5673 , n1655 );
buf ( n5674 , n2018 );
buf ( n5675 , n905 );
buf ( n5676 , n1025 );
buf ( n5677 , n1648 );
buf ( n5678 , n95 );
buf ( n5679 , n1852 );
buf ( n5680 , n1927 );
buf ( n5681 , n1215 );
buf ( n5682 , n473 );
buf ( n5683 , n742 );
buf ( n5684 , n846 );
buf ( n5685 , n1750 );
buf ( n5686 , n962 );
buf ( n5687 , n331 );
buf ( n5688 , n225 );
buf ( n5689 , n417 );
buf ( n5690 , n793 );
buf ( n5691 , n564 );
buf ( n5692 , n1495 );
buf ( n5693 , n515 );
buf ( n5694 , n571 );
buf ( n5695 , n1369 );
buf ( n5696 , n894 );
buf ( n5697 , n1151 );
buf ( n5698 , n867 );
buf ( n5699 , n1851 );
buf ( n5700 , n1661 );
buf ( n5701 , n2140 );
buf ( n5702 , n347 );
buf ( n5703 , n1134 );
buf ( n5704 , n1742 );
buf ( n5705 , n969 );
buf ( n5706 , n1744 );
buf ( n5707 , n1676 );
buf ( n5708 , n1854 );
buf ( n5709 , n1611 );
buf ( n5710 , n2025 );
buf ( n5711 , n663 );
buf ( n5712 , n514 );
buf ( n5713 , n1118 );
buf ( n5714 , n1156 );
buf ( n5715 , n2002 );
buf ( n5716 , n1337 );
buf ( n5717 , n28 );
buf ( n5718 , n244 );
buf ( n5719 , n273 );
buf ( n5720 , n757 );
buf ( n5721 , n69 );
buf ( n5722 , n882 );
buf ( n5723 , n1696 );
buf ( n5724 , n1858 );
buf ( n5725 , n602 );
buf ( n5726 , n1967 );
buf ( n5727 , n1983 );
buf ( n5728 , n607 );
buf ( n5729 , n1811 );
buf ( n5730 , n2127 );
buf ( n5731 , n351 );
buf ( n5732 , n1355 );
buf ( n5733 , n1175 );
buf ( n5734 , n192 );
buf ( n5735 , n699 );
buf ( n5736 , n864 );
buf ( n5737 , n1553 );
buf ( n5738 , n1451 );
buf ( n5739 , n1295 );
buf ( n5740 , n1874 );
buf ( n5741 , n545 );
buf ( n5742 , n724 );
buf ( n5743 , n973 );
buf ( n5744 , n837 );
buf ( n5745 , n342 );
buf ( n5746 , n1262 );
buf ( n5747 , n666 );
buf ( n5748 , n121 );
buf ( n5749 , n378 );
buf ( n5750 , n604 );
buf ( n5751 , n2133 );
buf ( n5752 , n1701 );
buf ( n5753 , n552 );
buf ( n5754 , n2097 );
buf ( n5755 , n1782 );
buf ( n5756 , n1253 );
buf ( n5757 , n631 );
buf ( n5758 , n1869 );
buf ( n5759 , n1597 );
buf ( n5760 , n233 );
buf ( n5761 , n205 );
buf ( n5762 , n135 );
buf ( n5763 , n761 );
buf ( n5764 , n613 );
buf ( n5765 , n2092 );
buf ( n5766 , n832 );
buf ( n5767 , n1233 );
buf ( n5768 , n1143 );
buf ( n5769 , n1972 );
buf ( n5770 , n114 );
buf ( n5771 , n304 );
buf ( n5772 , n1848 );
buf ( n5773 , n608 );
buf ( n5774 , n486 );
buf ( n5775 , n783 );
buf ( n5776 , n1649 );
buf ( n5777 , n667 );
buf ( n5778 , n492 );
buf ( n5779 , n1788 );
buf ( n5780 , n626 );
buf ( n5781 , n1006 );
buf ( n5782 , n1574 );
buf ( n5783 , n1726 );
buf ( n5784 , n24 );
buf ( n5785 , n1242 );
buf ( n5786 , n818 );
buf ( n5787 , n1240 );
buf ( n5788 , n1321 );
buf ( n5789 , n118 );
buf ( n5790 , n256 );
buf ( n5791 , n302 );
buf ( n5792 , n559 );
buf ( n5793 , n1728 );
buf ( n5794 , n72 );
buf ( n5795 , n1399 );
buf ( n5796 , n43 );
buf ( n5797 , n456 );
buf ( n5798 , n422 );
buf ( n5799 , n96 );
buf ( n5800 , n1304 );
buf ( n5801 , n1918 );
buf ( n5802 , n1722 );
buf ( n5803 , n698 );
buf ( n5804 , n2141 );
buf ( n5805 , n419 );
buf ( n5806 , n423 );
buf ( n5807 , n1310 );
buf ( n5808 , n637 );
buf ( n5809 , n1947 );
buf ( n5810 , n1807 );
buf ( n5811 , n1000 );
buf ( n5812 , n568 );
buf ( n5813 , n770 );
buf ( n5814 , n627 );
buf ( n5815 , n1738 );
buf ( n5816 , n1468 );
buf ( n5817 , n1572 );
buf ( n5818 , n437 );
buf ( n5819 , n822 );
buf ( n5820 , n632 );
buf ( n5821 , n1174 );
buf ( n5822 , n1654 );
buf ( n5823 , n1565 );
buf ( n5824 , n430 );
buf ( n5825 , n1630 );
buf ( n5826 , n1345 );
buf ( n5827 , n566 );
buf ( n5828 , n1780 );
buf ( n5829 , n2131 );
buf ( n5830 , n1439 );
buf ( n5831 , n269 );
buf ( n5832 , n937 );
buf ( n5833 , n1121 );
buf ( n5834 , n115 );
buf ( n5835 , n1605 );
buf ( n5836 , n1766 );
buf ( n5837 , n1613 );
buf ( n5838 , n1604 );
buf ( n5839 , n1645 );
buf ( n5840 , n1056 );
buf ( n5841 , n350 );
buf ( n5842 , n1734 );
buf ( n5843 , n890 );
buf ( n5844 , n2063 );
buf ( n5845 , n54 );
buf ( n5846 , n1306 );
buf ( n5847 , n1346 );
buf ( n5848 , n1886 );
buf ( n5849 , n117 );
buf ( n5850 , n875 );
buf ( n5851 , n1500 );
buf ( n5852 , n1545 );
buf ( n5853 , n1104 );
buf ( n5854 , n1775 );
buf ( n5855 , n1606 );
buf ( n5856 , n1020 );
buf ( n5857 , n1717 );
buf ( n5858 , n1916 );
buf ( n5859 , n1354 );
buf ( n5860 , n285 );
buf ( n5861 , n202 );
buf ( n5862 , n2030 );
buf ( n5863 , n897 );
buf ( n5864 , n1236 );
buf ( n5865 , n1957 );
buf ( n5866 , n359 );
buf ( n5867 , n610 );
buf ( n5868 , n429 );
buf ( n5869 , n339 );
buf ( n5870 , n623 );
buf ( n5871 , n1864 );
buf ( n5872 , n1960 );
buf ( n5873 , n565 );
buf ( n5874 , n78 );
buf ( n5875 , n1818 );
buf ( n5876 , n385 );
buf ( n5877 , n1012 );
buf ( n5878 , n668 );
buf ( n5879 , n1578 );
buf ( n5880 , n652 );
buf ( n5881 , n387 );
buf ( n5882 , n1441 );
buf ( n5883 , n550 );
buf ( n5884 , n279 );
buf ( n5885 , n531 );
buf ( n5886 , n411 );
buf ( n5887 , n1480 );
buf ( n5888 , n1758 );
buf ( n5889 , n906 );
buf ( n5890 , n1475 );
buf ( n5891 , n664 );
buf ( n5892 , n2126 );
buf ( n5893 , n105 );
buf ( n5894 , n493 );
buf ( n5895 , n589 );
buf ( n5896 , n506 );
buf ( n5897 , n1217 );
buf ( n5898 , n81 );
buf ( n5899 , n189 );
buf ( n5900 , n2073 );
buf ( n5901 , n126 );
buf ( n5902 , n31 );
buf ( n5903 , n1997 );
buf ( n5904 , n1188 );
buf ( n5905 , n239 );
buf ( n5906 , n1479 );
buf ( n5907 , n1614 );
buf ( n5908 , n2100 );
buf ( n5909 , n151 );
buf ( n5910 , n110 );
buf ( n5911 , n88 );
buf ( n5912 , n325 );
buf ( n5913 , n887 );
buf ( n5914 , n1973 );
buf ( n5915 , n1956 );
buf ( n5916 , n467 );
buf ( n5917 , n166 );
buf ( n5918 , n1627 );
buf ( n5919 , n2059 );
buf ( n5920 , n284 );
buf ( n5921 , n1013 );
buf ( n5922 , n800 );
buf ( n5923 , n1237 );
buf ( n5924 , n1296 );
buf ( n5925 , n1513 );
buf ( n5926 , n1996 );
buf ( n5927 , n1335 );
buf ( n5928 , n379 );
buf ( n5929 , n137 );
buf ( n5930 , n55 );
buf ( n5931 , n674 );
buf ( n5932 , n975 );
buf ( n5933 , n1498 );
buf ( n5934 , n1509 );
buf ( n5935 , n1009 );
buf ( n5936 , n635 );
buf ( n5937 , n642 );
buf ( n5938 , n755 );
buf ( n5939 , n736 );
buf ( n5940 , n1080 );
buf ( n5941 , n1586 );
buf ( n5942 , n1776 );
buf ( n5943 , n89 );
buf ( n5944 , n555 );
buf ( n5945 , n2139 );
buf ( n5946 , n326 );
buf ( n5947 , n297 );
buf ( n5948 , n1748 );
buf ( n5949 , n420 );
buf ( n5950 , n1166 );
buf ( n5951 , n541 );
buf ( n5952 , n2061 );
buf ( n5953 , n959 );
buf ( n5954 , n1588 );
buf ( n5955 , n1243 );
buf ( n5956 , n505 );
buf ( n5957 , n159 );
buf ( n5958 , n1423 );
buf ( n5959 , n696 );
buf ( n5960 , n336 );
buf ( n5961 , n1662 );
buf ( n5962 , n397 );
buf ( n5963 , n252 );
buf ( n5964 , n2007 );
buf ( n5965 , n1084 );
buf ( n5966 , n774 );
buf ( n5967 , n1113 );
buf ( n5968 , n1328 );
buf ( n5969 , n1058 );
buf ( n5970 , n286 );
buf ( n5971 , n120 );
buf ( n5972 , n2147 );
buf ( n5973 , n1459 );
buf ( n5974 , n1988 );
buf ( n5975 , n1132 );
buf ( n5976 , n1331 );
buf ( n5977 , n241 );
buf ( n5978 , n1470 );
buf ( n5979 , n1759 );
buf ( n5980 , n1446 );
buf ( n5981 , n488 );
buf ( n5982 , n1924 );
buf ( n5983 , n1719 );
buf ( n5984 , n858 );
buf ( n5985 , n138 );
buf ( n5986 , n963 );
buf ( n5987 , n1904 );
buf ( n5988 , n650 );
buf ( n5989 , n2125 );
buf ( n5990 , n1740 );
buf ( n5991 , n1101 );
buf ( n5992 , n704 );
buf ( n5993 , n581 );
buf ( n5994 , n1666 );
buf ( n5995 , n1879 );
buf ( n5996 , n300 );
buf ( n5997 , n80 );
buf ( n5998 , n1612 );
buf ( n5999 , n255 );
buf ( n6000 , n954 );
buf ( n6001 , n1727 );
buf ( n6002 , n215 );
buf ( n6003 , n945 );
buf ( n6004 , n870 );
buf ( n6005 , n2136 );
buf ( n6006 , n1581 );
buf ( n6007 , n1391 );
buf ( n6008 , n1915 );
buf ( n6009 , n1789 );
buf ( n6010 , n1129 );
buf ( n6011 , n29 );
buf ( n6012 , n377 );
buf ( n6013 , n6 );
buf ( n6014 , n1544 );
buf ( n6015 , n1936 );
buf ( n6016 , n17 );
buf ( n6017 , n1285 );
buf ( n6018 , n1846 );
buf ( n6019 , n712 );
buf ( n6020 , n1853 );
buf ( n6021 , n1693 );
buf ( n6022 , n1179 );
buf ( n6023 , n968 );
buf ( n6024 , n2057 );
buf ( n6025 , n585 );
buf ( n6026 , n1418 );
buf ( n6027 , n484 );
buf ( n6028 , n2005 );
buf ( n6029 , n989 );
buf ( n6030 , n1741 );
buf ( n6031 , n1228 );
buf ( n6032 , n1184 );
buf ( n6033 , n1520 );
buf ( n6034 , n1940 );
buf ( n6035 , n702 );
buf ( n6036 , n1533 );
buf ( n6037 , n2124 );
buf ( n6038 , n1078 );
buf ( n6039 , n640 );
buf ( n6040 , n852 );
buf ( n6041 , n902 );
buf ( n6042 , n690 );
buf ( n6043 , n2062 );
buf ( n6044 , n1528 );
buf ( n6045 , n1638 );
buf ( n6046 , n1257 );
buf ( n6047 , n1382 );
buf ( n6048 , n1576 );
buf ( n6049 , n1245 );
buf ( n6050 , n1892 );
buf ( n6051 , n1066 );
buf ( n6052 , n1235 );
buf ( n6053 , n1302 );
buf ( n6054 , n345 );
buf ( n6055 , n1923 );
buf ( n6056 , n1986 );
buf ( n6057 , n563 );
buf ( n6058 , n549 );
buf ( n6059 , n1205 );
buf ( n6060 , n741 );
buf ( n6061 , n1077 );
buf ( n6062 , n61 );
buf ( n6063 , n796 );
buf ( n6064 , n776 );
buf ( n6065 , n1212 );
buf ( n6066 , n871 );
buf ( n6067 , n1692 );
buf ( n6068 , n578 );
buf ( n6069 , n372 );
buf ( n6070 , n1059 );
buf ( n6071 , n1064 );
buf ( n6072 , n1765 );
buf ( n6073 , n917 );
buf ( n6074 , n1312 );
buf ( n6075 , n738 );
buf ( n6076 , n865 );
buf ( n6077 , n1969 );
buf ( n6078 , n1595 );
buf ( n6079 , n1798 );
buf ( n6080 , n1507 );
buf ( n6081 , n1105 );
buf ( n6082 , n1093 );
buf ( n6083 , n675 );
buf ( n6084 , n1333 );
buf ( n6085 , n1069 );
buf ( n6086 , n333 );
buf ( n6087 , n797 );
buf ( n6088 , n208 );
buf ( n6089 , n1573 );
buf ( n6090 , n936 );
buf ( n6091 , n13 );
buf ( n6092 , n729 );
buf ( n6093 , n1366 );
buf ( n6094 , n2143 );
buf ( n6095 , n1813 );
buf ( n6096 , n399 );
buf ( n6097 , n591 );
buf ( n6098 , n582 );
buf ( n6099 , n322 );
buf ( n6100 , n2106 );
buf ( n6101 , n1010 );
buf ( n6102 , n277 );
buf ( n6103 , n1146 );
buf ( n6104 , n648 );
buf ( n6105 , n1823 );
buf ( n6106 , n259 );
buf ( n6107 , n1476 );
buf ( n6108 , n1265 );
buf ( n6109 , n290 );
buf ( n6110 , n90 );
buf ( n6111 , n41 );
buf ( n6112 , n1746 );
buf ( n6113 , n1417 );
buf ( n6114 , n861 );
buf ( n6115 , n2075 );
buf ( n6116 , n125 );
buf ( n6117 , n1203 );
buf ( n6118 , n1835 );
buf ( n6119 , n828 );
buf ( n6120 , n953 );
buf ( n6121 , n1769 );
buf ( n6122 , n908 );
buf ( n6123 , n477 );
buf ( n6124 , n622 );
buf ( n6125 , n1723 );
buf ( n6126 , n329 );
buf ( n6127 , n1634 );
buf ( n6128 , n1416 );
buf ( n6129 , n2099 );
buf ( n6130 , n786 );
buf ( n6131 , n1396 );
buf ( n6132 , n2039 );
buf ( n6133 , n1256 );
buf ( n6134 , n525 );
buf ( n6135 , n401 );
buf ( n6136 , n1621 );
buf ( n6137 , n1368 );
buf ( n6138 , n2071 );
buf ( n6139 , n483 );
buf ( n6140 , n1268 );
buf ( n6141 , n1518 );
buf ( n6142 , n597 );
buf ( n6143 , n660 );
buf ( n6144 , n2011 );
buf ( n6145 , n2094 );
buf ( n6146 , n685 );
buf ( n6147 , n1200 );
buf ( n6148 , n1590 );
buf ( n6149 , n1778 );
buf ( n6150 , n1774 );
buf ( n6151 , n1593 );
buf ( n6152 , n272 );
buf ( n6153 , n1219 );
buf ( n6154 , n1667 );
buf ( n6155 , n1408 );
buf ( n6156 , n595 );
buf ( n6157 , n994 );
buf ( n6158 , n1147 );
buf ( n6159 , n1821 );
buf ( n6160 , n1761 );
buf ( n6161 , n1577 );
buf ( n6162 , n1330 );
buf ( n6163 , n1095 );
buf ( n6164 , n175 );
buf ( n6165 , n1796 );
buf ( n6166 , n204 );
buf ( n6167 , n1269 );
buf ( n6168 , n1162 );
buf ( n6169 , n1694 );
buf ( n6170 , n1663 );
buf ( n6171 , n519 );
buf ( n6172 , n1254 );
buf ( n6173 , n981 );
buf ( n6174 , n1626 );
buf ( n6175 , n52 );
buf ( n6176 , n237 );
buf ( n6177 , n721 );
buf ( n6178 , n859 );
buf ( n6179 , n1351 );
buf ( n6180 , n1555 );
buf ( n6181 , n1607 );
buf ( n6182 , n1684 );
buf ( n6183 , n2117 );
buf ( n6184 , n2118 );
buf ( n6185 , n1186 );
buf ( n6186 , n1735 );
buf ( n6187 , n1781 );
buf ( n6188 , n1877 );
buf ( n6189 , n1022 );
buf ( n6190 , n584 );
buf ( n6191 , n1227 );
buf ( n6192 , n358 );
buf ( n6193 , n463 );
buf ( n6194 , n1989 );
buf ( n6195 , n1633 );
buf ( n6196 , n1122 );
buf ( n6197 , n1453 );
buf ( n6198 , n634 );
buf ( n6199 , n1698 );
buf ( n6200 , n1982 );
buf ( n6201 , n1403 );
buf ( n6202 , n99 );
buf ( n6203 , n735 );
buf ( n6204 , n756 );
buf ( n6205 , n926 );
buf ( n6206 , n268 );
buf ( n6207 , n1566 );
buf ( n6208 , n289 );
buf ( n6209 , n1073 );
buf ( n6210 , n526 );
buf ( n6211 , n316 );
buf ( n6212 , n1299 );
buf ( n6213 , n1587 );
buf ( n6214 , n76 );
buf ( n6215 , n957 );
buf ( n6216 , n2008 );
buf ( n6217 , n1011 );
buf ( n6218 , n1053 );
buf ( n6219 , n455 );
buf ( n6220 , n36 );
buf ( n6221 , n1843 );
buf ( n6222 , n439 );
buf ( n6223 , n1035 );
buf ( n6224 , n474 );
buf ( n6225 , n677 );
buf ( n6226 , n178 );
buf ( n6227 , n2003 );
buf ( n6228 , n1137 );
buf ( n6229 , n548 );
buf ( n6230 , n221 );
buf ( n6231 , n1272 );
buf ( n6232 , n142 );
buf ( n6233 , n924 );
buf ( n6234 , n264 );
buf ( n6235 , n1352 );
buf ( n6236 , n1201 );
buf ( n6237 , n1499 );
buf ( n6238 , n496 );
buf ( n6239 , n567 );
buf ( n6240 , n1427 );
buf ( n6241 , n941 );
buf ( n6242 , n750 );
buf ( n6243 , n1097 );
buf ( n6244 , n693 );
buf ( n6245 , n1076 );
buf ( n6246 , n230 );
buf ( n6247 , n1278 );
buf ( n6248 , n845 );
buf ( n6249 , n63 );
buf ( n6250 , n213 );
buf ( n6251 , n2128 );
buf ( n6252 , n2040 );
buf ( n6253 , n705 );
buf ( n6254 , n958 );
buf ( n6255 , n1400 );
buf ( n6256 , n854 );
buf ( n6257 , n313 );
buf ( n6258 , n856 );
buf ( n6259 , n689 );
buf ( n6260 , n923 );
buf ( n6261 , n1679 );
buf ( n6262 , n1842 );
buf ( n6263 , n2142 );
buf ( n6264 , n1112 );
buf ( n6265 , n412 );
buf ( n6266 , n1289 );
buf ( n6267 , n162 );
buf ( n6268 , n282 );
buf ( n6269 , n1409 );
buf ( n6270 , n229 );
buf ( n6271 , n1029 );
buf ( n6272 , n195 );
buf ( n6273 , n155 );
buf ( n6274 , n1514 );
buf ( n6275 , n1402 );
buf ( n6276 , n1724 );
buf ( n6277 , n659 );
buf ( n6278 , n406 );
buf ( n6279 , n633 );
buf ( n6280 , n2035 );
buf ( n6281 , n1206 );
buf ( n6282 , n909 );
buf ( n6283 , n561 );
buf ( n6284 , n1880 );
buf ( n6285 , n337 );
buf ( n6286 , n389 );
buf ( n6287 , n1504 );
buf ( n6288 , n1945 );
buf ( n6289 , n1786 );
buf ( n6290 , n122 );
buf ( n6291 , n479 );
buf ( n6292 , n1259 );
buf ( n6293 , n547 );
buf ( n6294 , n537 );
buf ( n6295 , n160 );
buf ( n6296 , n806 );
buf ( n6297 , n1051 );
buf ( n6298 , n1921 );
buf ( n6299 , n851 );
buf ( n6300 , n1552 );
buf ( n6301 , n986 );
buf ( n6302 , n232 );
buf ( n6303 , n203 );
buf ( n6304 , n1384 );
buf ( n6305 , n586 );
buf ( n6306 , n1512 );
buf ( n6307 , n939 );
buf ( n6308 , n672 );
buf ( n6309 , n1002 );
buf ( n6310 , n2077 );
buf ( n6311 , n1816 );
buf ( n6312 , n451 );
buf ( n6313 , n971 );
buf ( n6314 , n706 );
buf ( n6315 , n1300 );
buf ( n6316 , n207 );
buf ( n6317 , n1167 );
buf ( n6318 , n424 );
buf ( n6319 , n1932 );
buf ( n6320 , n251 );
buf ( n6321 , n673 );
buf ( n6322 , n860 );
buf ( n6323 , n1953 );
buf ( n6324 , n2121 );
buf ( n6325 , n1211 );
buf ( n6326 , n1421 );
buf ( n6327 , n701 );
buf ( n6328 , n1148 );
buf ( n6329 , n258 );
buf ( n6330 , n1857 );
buf ( n6331 , n1637 );
buf ( n6332 , n1055 );
buf ( n6333 , n1847 );
buf ( n6334 , n128 );
buf ( n6335 , n1463 );
buf ( n6336 , n928 );
buf ( n6337 , n25 );
buf ( n6338 , n1288 );
buf ( n6339 , n1793 );
buf ( n6340 , n468 );
buf ( n6341 , n132 );
buf ( n6342 , n817 );
buf ( n6343 , n726 );
buf ( n6344 , n921 );
buf ( n6345 , n49 );
buf ( n6346 , n1120 );
buf ( n6347 , n611 );
buf ( n6348 , n308 );
buf ( n6349 , n1313 );
buf ( n6350 , n210 );
buf ( n6351 , n1373 );
buf ( n6352 , n1714 );
buf ( n6353 , n1763 );
buf ( n6354 , n1795 );
buf ( n6355 , n919 );
buf ( n6356 , n830 );
buf ( n6357 , n70 );
buf ( n6358 , n831 );
buf ( n6359 , n915 );
buf ( n6360 , n1270 );
buf ( n6361 , n127 );
buf ( n6362 , n319 );
buf ( n6363 , n1082 );
buf ( n6364 , n1343 );
buf ( n6365 , n482 );
buf ( n6366 , n820 );
buf ( n6367 , n1551 );
buf ( n6368 , n197 );
buf ( n6369 , n769 );
buf ( n6370 , n1371 );
buf ( n6371 , n1668 );
buf ( n6372 , n1422 );
buf ( n6373 , n321 );
buf ( n6374 , n1592 );
buf ( n6375 , n1689 );
buf ( n6376 , n2081 );
buf ( n6377 , n1534 );
buf ( n6378 , n1756 );
buf ( n6379 , n51 );
buf ( n6380 , n948 );
buf ( n6381 , n1348 );
buf ( n6382 , n713 );
buf ( n6383 , n265 );
buf ( n6384 , n116 );
buf ( n6385 , n348 );
buf ( n6386 , n1363 );
buf ( n6387 , n1968 );
buf ( n6388 , n1286 );
buf ( n6389 , n427 );
buf ( n6390 , n442 );
buf ( n6391 , n815 );
buf ( n6392 , n1386 );
buf ( n6393 , n152 );
buf ( n6394 , n307 );
buf ( n6395 , n2111 );
buf ( n6396 , n374 );
buf ( n6397 , n390 );
buf ( n6398 , n2110 );
buf ( n6399 , n885 );
buf ( n6400 , n653 );
buf ( n6401 , n575 );
buf ( n6402 , n641 );
buf ( n6403 , n903 );
buf ( n6404 , n718 );
buf ( n6405 , n1768 );
buf ( n6406 , n1524 );
buf ( n6407 , n435 );
buf ( n6408 , n2032 );
buf ( n6409 , n935 );
buf ( n6410 , n1899 );
buf ( n6411 , n1379 );
buf ( n6412 , n1292 );
buf ( n6413 , n124 );
buf ( n6414 , n1350 );
buf ( n6415 , n149 );
buf ( n6416 , n1164 );
buf ( n6417 , n46 );
buf ( n6418 , n2056 );
buf ( n6419 , n1477 );
buf ( n6420 , n469 );
buf ( n6421 , n1834 );
buf ( n6422 , n109 );
buf ( n6423 , n1317 );
buf ( n6424 , n1810 );
buf ( n6425 , n1582 );
buf ( n6426 , n590 );
buf ( n6427 , n238 );
buf ( n6428 , n14 );
buf ( n6429 , n553 );
buf ( n6430 , n799 );
buf ( n6431 , n217 );
buf ( n6432 , n1767 );
buf ( n6433 , n1489 );
buf ( n6434 , n97 );
buf ( n6435 , n616 );
buf ( n6436 , n1715 );
buf ( n6437 , n271 );
buf ( n6438 , n1090 );
buf ( n6439 , n341 );
buf ( n6440 , n950 );
buf ( n6441 , n734 );
buf ( n6442 , n1929 );
buf ( n6443 , n457 );
buf ( n6444 , n168 );
buf ( n6445 , n967 );
buf ( n6446 , n1712 );
buf ( n6447 , n2113 );
buf ( n6448 , n283 );
buf ( n6449 , n1817 );
buf ( n6450 , n1098 );
buf ( n6451 , n1820 );
buf ( n6452 , n1150 );
buf ( n6453 , n896 );
buf ( n6454 , n576 );
buf ( n6455 , n102 );
buf ( n6456 , n1990 );
buf ( n6457 , n2010 );
buf ( n6458 , n772 );
buf ( n6459 , n311 );
buf ( n6460 , n1704 );
buf ( n6461 , n2102 );
buf ( n6462 , n314 );
buf ( n6463 , n2132 );
buf ( n6464 , n434 );
buf ( n6465 , n630 );
buf ( n6466 , n759 );
buf ( n6467 , n44 );
buf ( n6468 , n196 );
buf ( n6469 , n4324 );
not ( n6470 , n6469 );
buf ( n6471 , n4325 );
buf ( n6472 , n4326 );
not ( n6473 , n6471 );
and ( n6474 , n6472 , n6473 );
or ( n6475 , n6471 , n6474 );
not ( n6476 , n6475 );
buf ( n6477 , n4327 );
and ( n6478 , n6476 , n6477 );
buf ( n6479 , n4328 );
not ( n6480 , n6474 );
buf ( n6481 , n4329 );
and ( n6482 , n6480 , n6481 );
buf ( n6483 , n4330 );
xor ( n6484 , n6483 , n6481 );
and ( n6485 , n6484 , n6474 );
or ( n6486 , n6482 , n6485 );
not ( n6487 , n6474 );
buf ( n6488 , n4331 );
and ( n6489 , n6487 , n6488 );
buf ( n6490 , n4332 );
xor ( n6491 , n6490 , n6488 );
and ( n6492 , n6491 , n6474 );
or ( n6493 , n6489 , n6492 );
xor ( n6494 , n6486 , n6493 );
buf ( n6495 , n4333 );
xor ( n6496 , n6494 , n6495 );
buf ( n6497 , n4334 );
xor ( n6498 , n6496 , n6497 );
buf ( n6499 , n4335 );
xor ( n6500 , n6498 , n6499 );
xor ( n6501 , n6479 , n6500 );
not ( n6502 , n6474 );
buf ( n6503 , n4336 );
and ( n6504 , n6502 , n6503 );
buf ( n6505 , n4337 );
xor ( n6506 , n6505 , n6503 );
and ( n6507 , n6506 , n6474 );
or ( n6508 , n6504 , n6507 );
buf ( n6509 , n4338 );
xor ( n6510 , n6508 , n6509 );
buf ( n6511 , n4339 );
xor ( n6512 , n6510 , n6511 );
buf ( n6513 , n4340 );
xor ( n6514 , n6512 , n6513 );
buf ( n6515 , n4341 );
xor ( n6516 , n6514 , n6515 );
xor ( n6517 , n6501 , n6516 );
buf ( n6518 , n4342 );
not ( n6519 , n6474 );
not ( n6520 , n4343 );
buf ( n6521 , n6520 );
and ( n6522 , n6519 , n6521 );
buf ( n6523 , n6474 );
or ( n6524 , n6522 , n6523 );
not ( n6525 , n6474 );
buf ( n6526 , n4344 );
and ( n6527 , n6525 , n6526 );
buf ( n6528 , n4345 );
xor ( n6529 , n6528 , n6526 );
and ( n6530 , n6529 , n6474 );
or ( n6531 , n6527 , n6530 );
xor ( n6532 , n6524 , n6531 );
buf ( n6533 , n4346 );
xor ( n6534 , n6532 , n6533 );
buf ( n6535 , n4347 );
xor ( n6536 , n6534 , n6535 );
buf ( n6537 , n4348 );
xor ( n6538 , n6536 , n6537 );
xor ( n6539 , n6518 , n6538 );
not ( n6540 , n6474 );
buf ( n6541 , n4349 );
and ( n6542 , n6540 , n6541 );
buf ( n6543 , n4350 );
xor ( n6544 , n6543 , n6541 );
and ( n6545 , n6544 , n6474 );
or ( n6546 , n6542 , n6545 );
not ( n6547 , n6474 );
buf ( n6548 , n4351 );
and ( n6549 , n6547 , n6548 );
buf ( n6550 , n4352 );
xor ( n6551 , n6550 , n6548 );
and ( n6552 , n6551 , n6474 );
or ( n6553 , n6549 , n6552 );
xor ( n6554 , n6546 , n6553 );
buf ( n6555 , n4353 );
xor ( n6556 , n6554 , n6555 );
buf ( n6557 , n4354 );
xor ( n6558 , n6556 , n6557 );
buf ( n6559 , n4355 );
xor ( n6560 , n6558 , n6559 );
xor ( n6561 , n6539 , n6560 );
not ( n6562 , n6561 );
not ( n6563 , n6474 );
buf ( n6564 , n4356 );
and ( n6565 , n6563 , n6564 );
buf ( n6566 , n4357 );
xor ( n6567 , n6566 , n6564 );
and ( n6568 , n6567 , n6474 );
or ( n6569 , n6565 , n6568 );
not ( n6570 , n6474 );
buf ( n6571 , n4358 );
and ( n6572 , n6570 , n6571 );
buf ( n6573 , n4359 );
xor ( n6574 , n6573 , n6571 );
and ( n6575 , n6574 , n6474 );
or ( n6576 , n6572 , n6575 );
buf ( n6577 , n4360 );
xor ( n6578 , n6576 , n6577 );
buf ( n6579 , n4361 );
xor ( n6580 , n6578 , n6579 );
buf ( n6581 , n4362 );
xor ( n6582 , n6580 , n6581 );
buf ( n6583 , n4363 );
xor ( n6584 , n6582 , n6583 );
xor ( n6585 , n6569 , n6584 );
not ( n6586 , n6474 );
buf ( n6587 , n4364 );
and ( n6588 , n6586 , n6587 );
buf ( n6589 , n4365 );
xor ( n6590 , n6589 , n6587 );
and ( n6591 , n6590 , n6474 );
or ( n6592 , n6588 , n6591 );
not ( n6593 , n6474 );
buf ( n6594 , n4366 );
and ( n6595 , n6593 , n6594 );
buf ( n6596 , n4367 );
xor ( n6597 , n6596 , n6594 );
and ( n6598 , n6597 , n6474 );
or ( n6599 , n6595 , n6598 );
xor ( n6600 , n6592 , n6599 );
buf ( n6601 , n4368 );
xor ( n6602 , n6600 , n6601 );
buf ( n6603 , n4369 );
xor ( n6604 , n6602 , n6603 );
buf ( n6605 , n4370 );
xor ( n6606 , n6604 , n6605 );
xor ( n6607 , n6585 , n6606 );
and ( n6608 , n6562 , n6607 );
xor ( n6609 , n6517 , n6608 );
buf ( n6610 , n4371 );
not ( n6611 , n6474 );
buf ( n6612 , n4372 );
and ( n6613 , n6611 , n6612 );
buf ( n6614 , n4373 );
xor ( n6615 , n6614 , n6612 );
and ( n6616 , n6615 , n6474 );
or ( n6617 , n6613 , n6616 );
not ( n6618 , n6474 );
buf ( n6619 , n4374 );
and ( n6620 , n6618 , n6619 );
buf ( n6621 , n4375 );
xor ( n6622 , n6621 , n6619 );
and ( n6623 , n6622 , n6474 );
or ( n6624 , n6620 , n6623 );
xor ( n6625 , n6617 , n6624 );
buf ( n6626 , n4376 );
xor ( n6627 , n6625 , n6626 );
buf ( n6628 , n4377 );
xor ( n6629 , n6627 , n6628 );
buf ( n6630 , n4378 );
xor ( n6631 , n6629 , n6630 );
xor ( n6632 , n6610 , n6631 );
not ( n6633 , n6474 );
buf ( n6634 , n4379 );
and ( n6635 , n6633 , n6634 );
buf ( n6636 , n4380 );
xor ( n6637 , n6636 , n6634 );
and ( n6638 , n6637 , n6474 );
or ( n6639 , n6635 , n6638 );
not ( n6640 , n6474 );
buf ( n6641 , n4381 );
and ( n6642 , n6640 , n6641 );
buf ( n6643 , n4382 );
xor ( n6644 , n6643 , n6641 );
and ( n6645 , n6644 , n6474 );
or ( n6646 , n6642 , n6645 );
xor ( n6647 , n6639 , n6646 );
buf ( n6648 , n4383 );
xor ( n6649 , n6647 , n6648 );
buf ( n6650 , n4384 );
xor ( n6651 , n6649 , n6650 );
buf ( n6652 , n4385 );
xor ( n6653 , n6651 , n6652 );
xor ( n6654 , n6632 , n6653 );
not ( n6655 , n6517 );
and ( n6656 , n6655 , n6561 );
xor ( n6657 , n6654 , n6656 );
buf ( n6658 , n4386 );
not ( n6659 , n6474 );
buf ( n6660 , n4387 );
and ( n6661 , n6659 , n6660 );
buf ( n6662 , n4388 );
xor ( n6663 , n6662 , n6660 );
and ( n6664 , n6663 , n6474 );
or ( n6665 , n6661 , n6664 );
buf ( n6666 , n4389 );
xor ( n6667 , n6665 , n6666 );
buf ( n6668 , n4390 );
xor ( n6669 , n6667 , n6668 );
buf ( n6670 , n4391 );
xor ( n6671 , n6669 , n6670 );
buf ( n6672 , n4392 );
xor ( n6673 , n6671 , n6672 );
xor ( n6674 , n6658 , n6673 );
not ( n6675 , n6474 );
buf ( n6676 , n4393 );
and ( n6677 , n6675 , n6676 );
buf ( n6678 , n4394 );
xor ( n6679 , n6678 , n6676 );
and ( n6680 , n6679 , n6474 );
or ( n6681 , n6677 , n6680 );
not ( n6682 , n6474 );
buf ( n6683 , n4395 );
and ( n6684 , n6682 , n6683 );
buf ( n6685 , n4396 );
xor ( n6686 , n6685 , n6683 );
and ( n6687 , n6686 , n6474 );
or ( n6688 , n6684 , n6687 );
xor ( n6689 , n6681 , n6688 );
buf ( n6690 , n4397 );
xor ( n6691 , n6689 , n6690 );
buf ( n6692 , n4398 );
xor ( n6693 , n6691 , n6692 );
buf ( n6694 , n4399 );
xor ( n6695 , n6693 , n6694 );
xor ( n6696 , n6674 , n6695 );
buf ( n6697 , n4400 );
not ( n6698 , n6474 );
buf ( n6699 , n4401 );
and ( n6700 , n6698 , n6699 );
buf ( n6701 , n6699 );
and ( n6702 , n6701 , n6474 );
or ( n6703 , n6700 , n6702 );
not ( n6704 , n6474 );
buf ( n6705 , n4402 );
and ( n6706 , n6704 , n6705 );
buf ( n6707 , n4403 );
xor ( n6708 , n6707 , n6705 );
and ( n6709 , n6708 , n6474 );
or ( n6710 , n6706 , n6709 );
xor ( n6711 , n6703 , n6710 );
buf ( n6712 , n4404 );
xor ( n6713 , n6711 , n6712 );
buf ( n6714 , n4405 );
xor ( n6715 , n6713 , n6714 );
buf ( n6716 , n4406 );
xor ( n6717 , n6715 , n6716 );
xor ( n6718 , n6697 , n6717 );
not ( n6719 , n6474 );
buf ( n6720 , n4407 );
and ( n6721 , n6719 , n6720 );
buf ( n6722 , n4408 );
xor ( n6723 , n6722 , n6720 );
and ( n6724 , n6723 , n6474 );
or ( n6725 , n6721 , n6724 );
not ( n6726 , n6474 );
buf ( n6727 , n4409 );
and ( n6728 , n6726 , n6727 );
buf ( n6729 , n4410 );
xor ( n6730 , n6729 , n6727 );
and ( n6731 , n6730 , n6474 );
or ( n6732 , n6728 , n6731 );
xor ( n6733 , n6725 , n6732 );
buf ( n6734 , n4411 );
xor ( n6735 , n6733 , n6734 );
buf ( n6736 , n4412 );
xor ( n6737 , n6735 , n6736 );
buf ( n6738 , n4413 );
xor ( n6739 , n6737 , n6738 );
xor ( n6740 , n6718 , n6739 );
not ( n6741 , n6740 );
buf ( n6742 , n4414 );
not ( n6743 , n6474 );
buf ( n6744 , n4415 );
and ( n6745 , n6743 , n6744 );
buf ( n6746 , n4416 );
xor ( n6747 , n6746 , n6744 );
and ( n6748 , n6747 , n6474 );
or ( n6749 , n6745 , n6748 );
not ( n6750 , n6474 );
buf ( n6751 , n4417 );
and ( n6752 , n6750 , n6751 );
buf ( n6753 , n4418 );
xor ( n6754 , n6753 , n6751 );
and ( n6755 , n6754 , n6474 );
or ( n6756 , n6752 , n6755 );
xor ( n6757 , n6749 , n6756 );
buf ( n6758 , n4419 );
xor ( n6759 , n6757 , n6758 );
buf ( n6760 , n4420 );
xor ( n6761 , n6759 , n6760 );
buf ( n6762 , n4421 );
xor ( n6763 , n6761 , n6762 );
xor ( n6764 , n6742 , n6763 );
not ( n6765 , n6474 );
buf ( n6766 , n4422 );
and ( n6767 , n6765 , n6766 );
buf ( n6768 , n4423 );
xor ( n6769 , n6768 , n6766 );
and ( n6770 , n6769 , n6474 );
or ( n6771 , n6767 , n6770 );
not ( n6772 , n6474 );
buf ( n6773 , n4424 );
and ( n6774 , n6772 , n6773 );
buf ( n6775 , n4425 );
xor ( n6776 , n6775 , n6773 );
and ( n6777 , n6776 , n6474 );
or ( n6778 , n6774 , n6777 );
xor ( n6779 , n6771 , n6778 );
buf ( n6780 , n4426 );
xor ( n6781 , n6779 , n6780 );
buf ( n6782 , n4427 );
xor ( n6783 , n6781 , n6782 );
buf ( n6784 , n4428 );
xor ( n6785 , n6783 , n6784 );
xor ( n6786 , n6764 , n6785 );
and ( n6787 , n6741 , n6786 );
xor ( n6788 , n6696 , n6787 );
xor ( n6789 , n6657 , n6788 );
buf ( n6790 , n4429 );
not ( n6791 , n6474 );
buf ( n6792 , n4430 );
and ( n6793 , n6791 , n6792 );
buf ( n6794 , n4431 );
xor ( n6795 , n6794 , n6792 );
and ( n6796 , n6795 , n6474 );
or ( n6797 , n6793 , n6796 );
not ( n6798 , n6474 );
buf ( n6799 , n4432 );
and ( n6800 , n6798 , n6799 );
buf ( n6801 , n4433 );
xor ( n6802 , n6801 , n6799 );
and ( n6803 , n6802 , n6474 );
or ( n6804 , n6800 , n6803 );
xor ( n6805 , n6797 , n6804 );
buf ( n6806 , n4434 );
xor ( n6807 , n6805 , n6806 );
buf ( n6808 , n4435 );
xor ( n6809 , n6807 , n6808 );
buf ( n6810 , n4436 );
xor ( n6811 , n6809 , n6810 );
xor ( n6812 , n6790 , n6811 );
not ( n6813 , n6474 );
buf ( n6814 , n4437 );
and ( n6815 , n6813 , n6814 );
buf ( n6816 , n4438 );
xor ( n6817 , n6816 , n6814 );
and ( n6818 , n6817 , n6474 );
or ( n6819 , n6815 , n6818 );
buf ( n6820 , n4439 );
xor ( n6821 , n6819 , n6820 );
buf ( n6822 , n4440 );
xor ( n6823 , n6821 , n6822 );
buf ( n6824 , n4441 );
xor ( n6825 , n6823 , n6824 );
buf ( n6826 , n4442 );
xor ( n6827 , n6825 , n6826 );
xor ( n6828 , n6812 , n6827 );
buf ( n6829 , n4443 );
not ( n6830 , n6474 );
buf ( n6831 , n4444 );
and ( n6832 , n6830 , n6831 );
buf ( n6833 , n4445 );
xor ( n6834 , n6833 , n6831 );
and ( n6835 , n6834 , n6474 );
or ( n6836 , n6832 , n6835 );
not ( n6837 , n6474 );
buf ( n6838 , n4446 );
and ( n6839 , n6837 , n6838 );
buf ( n6840 , n4447 );
xor ( n6841 , n6840 , n6838 );
and ( n6842 , n6841 , n6474 );
or ( n6843 , n6839 , n6842 );
xor ( n6844 , n6836 , n6843 );
buf ( n6845 , n4448 );
xor ( n6846 , n6844 , n6845 );
buf ( n6847 , n4449 );
xor ( n6848 , n6846 , n6847 );
buf ( n6849 , n4450 );
xor ( n6850 , n6848 , n6849 );
xor ( n6851 , n6829 , n6850 );
not ( n6852 , n6474 );
buf ( n6853 , n4451 );
and ( n6854 , n6852 , n6853 );
buf ( n6855 , n4452 );
xor ( n6856 , n6855 , n6853 );
and ( n6857 , n6856 , n6474 );
or ( n6858 , n6854 , n6857 );
not ( n6859 , n6474 );
buf ( n6860 , n4453 );
and ( n6861 , n6859 , n6860 );
buf ( n6862 , n4454 );
xor ( n6863 , n6862 , n6860 );
and ( n6864 , n6863 , n6474 );
or ( n6865 , n6861 , n6864 );
xor ( n6866 , n6858 , n6865 );
buf ( n6867 , n4455 );
xor ( n6868 , n6866 , n6867 );
buf ( n6869 , n4456 );
xor ( n6870 , n6868 , n6869 );
buf ( n6871 , n4457 );
xor ( n6872 , n6870 , n6871 );
xor ( n6873 , n6851 , n6872 );
not ( n6874 , n6873 );
buf ( n6875 , n4458 );
not ( n6876 , n6474 );
buf ( n6877 , n4459 );
and ( n6878 , n6876 , n6877 );
buf ( n6879 , n4460 );
xor ( n6880 , n6879 , n6877 );
and ( n6881 , n6880 , n6474 );
or ( n6882 , n6878 , n6881 );
buf ( n6883 , n4461 );
xor ( n6884 , n6882 , n6883 );
buf ( n6885 , n4462 );
xor ( n6886 , n6884 , n6885 );
buf ( n6887 , n4463 );
buf ( n6888 , n6887 );
xor ( n6889 , n6886 , n6888 );
buf ( n6890 , n4464 );
xor ( n6891 , n6889 , n6890 );
xor ( n6892 , n6875 , n6891 );
not ( n6893 , n6474 );
buf ( n6894 , n4465 );
and ( n6895 , n6893 , n6894 );
buf ( n6896 , n4466 );
xor ( n6897 , n6896 , n6894 );
and ( n6898 , n6897 , n6474 );
or ( n6899 , n6895 , n6898 );
not ( n6900 , n6474 );
buf ( n6901 , n4467 );
and ( n6902 , n6900 , n6901 );
buf ( n6903 , n4468 );
xor ( n6904 , n6903 , n6901 );
and ( n6905 , n6904 , n6474 );
or ( n6906 , n6902 , n6905 );
xor ( n6907 , n6899 , n6906 );
buf ( n6908 , n4469 );
xor ( n6909 , n6907 , n6908 );
buf ( n6910 , n4470 );
xor ( n6911 , n6909 , n6910 );
buf ( n6912 , n4471 );
xor ( n6913 , n6911 , n6912 );
xor ( n6914 , n6892 , n6913 );
and ( n6915 , n6874 , n6914 );
xor ( n6916 , n6828 , n6915 );
xor ( n6917 , n6789 , n6916 );
buf ( n6918 , n4472 );
not ( n6919 , n6474 );
buf ( n6920 , n4473 );
and ( n6921 , n6919 , n6920 );
buf ( n6922 , n4474 );
xor ( n6923 , n6922 , n6920 );
and ( n6924 , n6923 , n6474 );
or ( n6925 , n6921 , n6924 );
not ( n6926 , n6474 );
buf ( n6927 , n4475 );
and ( n6928 , n6926 , n6927 );
buf ( n6929 , n4476 );
xor ( n6930 , n6929 , n6927 );
and ( n6931 , n6930 , n6474 );
or ( n6932 , n6928 , n6931 );
xor ( n6933 , n6925 , n6932 );
buf ( n6934 , n4477 );
xor ( n6935 , n6933 , n6934 );
buf ( n6936 , n4478 );
xor ( n6937 , n6935 , n6936 );
buf ( n6938 , n4479 );
xor ( n6939 , n6937 , n6938 );
xor ( n6940 , n6918 , n6939 );
not ( n6941 , n6474 );
buf ( n6942 , n4480 );
and ( n6943 , n6941 , n6942 );
buf ( n6944 , n4481 );
xor ( n6945 , n6944 , n6942 );
and ( n6946 , n6945 , n6474 );
or ( n6947 , n6943 , n6946 );
not ( n6948 , n6474 );
buf ( n6949 , n4482 );
and ( n6950 , n6948 , n6949 );
buf ( n6951 , n4483 );
xor ( n6952 , n6951 , n6949 );
and ( n6953 , n6952 , n6474 );
or ( n6954 , n6950 , n6953 );
xor ( n6955 , n6947 , n6954 );
buf ( n6956 , n4484 );
xor ( n6957 , n6955 , n6956 );
buf ( n6958 , n4485 );
xor ( n6959 , n6957 , n6958 );
buf ( n6960 , n4486 );
xor ( n6961 , n6959 , n6960 );
xor ( n6962 , n6940 , n6961 );
buf ( n6963 , n4487 );
not ( n6964 , n6474 );
buf ( n6965 , n4488 );
and ( n6966 , n6964 , n6965 );
buf ( n6967 , n4489 );
xor ( n6968 , n6967 , n6965 );
and ( n6969 , n6968 , n6474 );
or ( n6970 , n6966 , n6969 );
not ( n6971 , n6474 );
buf ( n6972 , n4490 );
and ( n6973 , n6971 , n6972 );
buf ( n6974 , n4491 );
xor ( n6975 , n6974 , n6972 );
and ( n6976 , n6975 , n6474 );
or ( n6977 , n6973 , n6976 );
xor ( n6978 , n6970 , n6977 );
buf ( n6979 , n4492 );
xor ( n6980 , n6978 , n6979 );
buf ( n6981 , n4493 );
xor ( n6982 , n6980 , n6981 );
buf ( n6983 , n4494 );
xor ( n6984 , n6982 , n6983 );
xor ( n6985 , n6963 , n6984 );
not ( n6986 , n6474 );
buf ( n6987 , n4495 );
and ( n6988 , n6986 , n6987 );
buf ( n6989 , n4496 );
xor ( n6990 , n6989 , n6987 );
and ( n6991 , n6990 , n6474 );
or ( n6992 , n6988 , n6991 );
not ( n6993 , n6474 );
buf ( n6994 , n4497 );
and ( n6995 , n6993 , n6994 );
buf ( n6996 , n4498 );
xor ( n6997 , n6996 , n6994 );
and ( n6998 , n6997 , n6474 );
or ( n6999 , n6995 , n6998 );
xor ( n7000 , n6992 , n6999 );
buf ( n7001 , n4499 );
xor ( n7002 , n7000 , n7001 );
buf ( n7003 , n4500 );
xor ( n7004 , n7002 , n7003 );
buf ( n7005 , n4501 );
xor ( n7006 , n7004 , n7005 );
xor ( n7007 , n6985 , n7006 );
not ( n7008 , n7007 );
buf ( n7009 , n4502 );
not ( n7010 , n6474 );
buf ( n7011 , n4503 );
and ( n7012 , n7010 , n7011 );
buf ( n7013 , n4504 );
xor ( n7014 , n7013 , n7011 );
and ( n7015 , n7014 , n6474 );
or ( n7016 , n7012 , n7015 );
not ( n7017 , n6474 );
buf ( n7018 , n4505 );
and ( n7019 , n7017 , n7018 );
buf ( n7020 , n4506 );
xor ( n7021 , n7020 , n7018 );
and ( n7022 , n7021 , n6474 );
or ( n7023 , n7019 , n7022 );
xor ( n7024 , n7016 , n7023 );
buf ( n7025 , n4507 );
xor ( n7026 , n7024 , n7025 );
buf ( n7027 , n4508 );
xor ( n7028 , n7026 , n7027 );
buf ( n7029 , n4509 );
xor ( n7030 , n7028 , n7029 );
xor ( n7031 , n7009 , n7030 );
not ( n7032 , n6474 );
buf ( n7033 , n4510 );
and ( n7034 , n7032 , n7033 );
buf ( n7035 , n4511 );
xor ( n7036 , n7035 , n7033 );
and ( n7037 , n7036 , n6474 );
or ( n7038 , n7034 , n7037 );
buf ( n7039 , n4512 );
xor ( n7040 , n7038 , n7039 );
buf ( n7041 , n4513 );
xor ( n7042 , n7040 , n7041 );
buf ( n7043 , n4514 );
xor ( n7044 , n7042 , n7043 );
buf ( n7045 , n4515 );
xor ( n7046 , n7044 , n7045 );
xor ( n7047 , n7031 , n7046 );
and ( n7048 , n7008 , n7047 );
xor ( n7049 , n6962 , n7048 );
xor ( n7050 , n6917 , n7049 );
buf ( n7051 , n4516 );
not ( n7052 , n6474 );
buf ( n7053 , n4517 );
and ( n7054 , n7052 , n7053 );
buf ( n7055 , n4518 );
xor ( n7056 , n7055 , n7053 );
and ( n7057 , n7056 , n6474 );
or ( n7058 , n7054 , n7057 );
not ( n7059 , n6474 );
buf ( n7060 , n4519 );
and ( n7061 , n7059 , n7060 );
buf ( n7062 , n4520 );
xor ( n7063 , n7062 , n7060 );
and ( n7064 , n7063 , n6474 );
or ( n7065 , n7061 , n7064 );
xor ( n7066 , n7058 , n7065 );
buf ( n7067 , n4521 );
xor ( n7068 , n7066 , n7067 );
buf ( n7069 , n4522 );
xor ( n7070 , n7068 , n7069 );
buf ( n7071 , n4523 );
xor ( n7072 , n7070 , n7071 );
xor ( n7073 , n7051 , n7072 );
not ( n7074 , n6474 );
buf ( n7075 , n4524 );
and ( n7076 , n7074 , n7075 );
buf ( n7077 , n4525 );
xor ( n7078 , n7077 , n7075 );
and ( n7079 , n7078 , n6474 );
or ( n7080 , n7076 , n7079 );
not ( n7081 , n6474 );
buf ( n7082 , n4526 );
and ( n7083 , n7081 , n7082 );
buf ( n7084 , n4527 );
xor ( n7085 , n7084 , n7082 );
and ( n7086 , n7085 , n6474 );
or ( n7087 , n7083 , n7086 );
xor ( n7088 , n7080 , n7087 );
buf ( n7089 , n4528 );
xor ( n7090 , n7088 , n7089 );
buf ( n7091 , n4529 );
buf ( n7092 , n7091 );
xor ( n7093 , n7090 , n7092 );
buf ( n7094 , n4530 );
xor ( n7095 , n7093 , n7094 );
xor ( n7096 , n7073 , n7095 );
buf ( n7097 , n4531 );
not ( n7098 , n6474 );
buf ( n7099 , n4532 );
and ( n7100 , n7098 , n7099 );
buf ( n7101 , n4533 );
xor ( n7102 , n7101 , n7099 );
and ( n7103 , n7102 , n6474 );
or ( n7104 , n7100 , n7103 );
buf ( n7105 , n4534 );
xor ( n7106 , n7104 , n7105 );
buf ( n7107 , n4535 );
xor ( n7108 , n7106 , n7107 );
buf ( n7109 , n4536 );
xor ( n7110 , n7108 , n7109 );
buf ( n7111 , n4537 );
xor ( n7112 , n7110 , n7111 );
xor ( n7113 , n7097 , n7112 );
not ( n7114 , n6474 );
buf ( n7115 , n4538 );
and ( n7116 , n7114 , n7115 );
buf ( n7117 , n4539 );
xor ( n7118 , n7117 , n7115 );
and ( n7119 , n7118 , n6474 );
or ( n7120 , n7116 , n7119 );
not ( n7121 , n6474 );
buf ( n7122 , n4540 );
and ( n7123 , n7121 , n7122 );
buf ( n7124 , n4541 );
xor ( n7125 , n7124 , n7122 );
and ( n7126 , n7125 , n6474 );
or ( n7127 , n7123 , n7126 );
xor ( n7128 , n7120 , n7127 );
buf ( n7129 , n4542 );
xor ( n7130 , n7128 , n7129 );
buf ( n7131 , n4543 );
xor ( n7132 , n7130 , n7131 );
buf ( n7133 , n4544 );
xor ( n7134 , n7132 , n7133 );
xor ( n7135 , n7113 , n7134 );
not ( n7136 , n7135 );
buf ( n7137 , n4545 );
not ( n7138 , n6474 );
buf ( n7139 , n4546 );
and ( n7140 , n7138 , n7139 );
buf ( n7141 , n4547 );
xor ( n7142 , n7141 , n7139 );
and ( n7143 , n7142 , n6474 );
or ( n7144 , n7140 , n7143 );
not ( n7145 , n6474 );
buf ( n7146 , n4548 );
and ( n7147 , n7145 , n7146 );
buf ( n7148 , n4549 );
xor ( n7149 , n7148 , n7146 );
and ( n7150 , n7149 , n6474 );
or ( n7151 , n7147 , n7150 );
xor ( n7152 , n7144 , n7151 );
buf ( n7153 , n4550 );
xor ( n7154 , n7152 , n7153 );
buf ( n7155 , n4551 );
xor ( n7156 , n7154 , n7155 );
buf ( n7157 , n4552 );
buf ( n7158 , n7157 );
xor ( n7159 , n7156 , n7158 );
xor ( n7160 , n7137 , n7159 );
not ( n7161 , n6474 );
buf ( n7162 , n4553 );
and ( n7163 , n7161 , n7162 );
buf ( n7164 , n4554 );
xor ( n7165 , n7164 , n7162 );
and ( n7166 , n7165 , n6474 );
or ( n7167 , n7163 , n7166 );
not ( n7168 , n6474 );
buf ( n7169 , n4555 );
and ( n7170 , n7168 , n7169 );
buf ( n7171 , n4556 );
xor ( n7172 , n7171 , n7169 );
and ( n7173 , n7172 , n6474 );
or ( n7174 , n7170 , n7173 );
xor ( n7175 , n7167 , n7174 );
buf ( n7176 , n4557 );
xor ( n7177 , n7175 , n7176 );
buf ( n7178 , n4558 );
xor ( n7179 , n7177 , n7178 );
buf ( n7180 , n4559 );
xor ( n7181 , n7179 , n7180 );
xor ( n7182 , n7160 , n7181 );
and ( n7183 , n7136 , n7182 );
xor ( n7184 , n7096 , n7183 );
xor ( n7185 , n7050 , n7184 );
xor ( n7186 , n6609 , n7185 );
buf ( n7187 , n4560 );
not ( n7188 , n6474 );
buf ( n7189 , n4561 );
and ( n7190 , n7188 , n7189 );
buf ( n7191 , n4562 );
xor ( n7192 , n7191 , n7189 );
and ( n7193 , n7192 , n6474 );
or ( n7194 , n7190 , n7193 );
not ( n7195 , n6474 );
buf ( n7196 , n4563 );
and ( n7197 , n7195 , n7196 );
buf ( n7198 , n4564 );
xor ( n7199 , n7198 , n7196 );
and ( n7200 , n7199 , n6474 );
or ( n7201 , n7197 , n7200 );
xor ( n7202 , n7194 , n7201 );
buf ( n7203 , n4565 );
xor ( n7204 , n7202 , n7203 );
buf ( n7205 , n4566 );
xor ( n7206 , n7204 , n7205 );
buf ( n7207 , n4567 );
xor ( n7208 , n7206 , n7207 );
xor ( n7209 , n7187 , n7208 );
not ( n7210 , n6474 );
buf ( n7211 , n4568 );
and ( n7212 , n7210 , n7211 );
buf ( n7213 , n4569 );
xor ( n7214 , n7213 , n7211 );
and ( n7215 , n7214 , n6474 );
or ( n7216 , n7212 , n7215 );
not ( n7217 , n6474 );
buf ( n7218 , n4570 );
and ( n7219 , n7217 , n7218 );
buf ( n7220 , n4571 );
xor ( n7221 , n7220 , n7218 );
and ( n7222 , n7221 , n6474 );
or ( n7223 , n7219 , n7222 );
xor ( n7224 , n7216 , n7223 );
buf ( n7225 , n4572 );
xor ( n7226 , n7224 , n7225 );
buf ( n7227 , n4573 );
xor ( n7228 , n7226 , n7227 );
buf ( n7229 , n4574 );
xor ( n7230 , n7228 , n7229 );
xor ( n7231 , n7209 , n7230 );
not ( n7232 , n6474 );
buf ( n7233 , n4575 );
and ( n7234 , n7232 , n7233 );
buf ( n7235 , n4576 );
xor ( n7236 , n7235 , n7233 );
and ( n7237 , n7236 , n6474 );
or ( n7238 , n7234 , n7237 );
not ( n7239 , n6474 );
buf ( n7240 , n4577 );
and ( n7241 , n7239 , n7240 );
buf ( n7242 , n4578 );
xor ( n7243 , n7242 , n7240 );
and ( n7244 , n7243 , n6474 );
or ( n7245 , n7241 , n7244 );
buf ( n7246 , n4579 );
xor ( n7247 , n7245 , n7246 );
buf ( n7248 , n4580 );
xor ( n7249 , n7247 , n7248 );
buf ( n7250 , n4581 );
xor ( n7251 , n7249 , n7250 );
buf ( n7252 , n4582 );
xor ( n7253 , n7251 , n7252 );
xor ( n7254 , n7238 , n7253 );
not ( n7255 , n6474 );
buf ( n7256 , n4583 );
and ( n7257 , n7255 , n7256 );
buf ( n7258 , n4584 );
xor ( n7259 , n7258 , n7256 );
and ( n7260 , n7259 , n6474 );
or ( n7261 , n7257 , n7260 );
not ( n7262 , n6474 );
buf ( n7263 , n4585 );
and ( n7264 , n7262 , n7263 );
buf ( n7265 , n4586 );
xor ( n7266 , n7265 , n7263 );
and ( n7267 , n7266 , n6474 );
or ( n7268 , n7264 , n7267 );
xor ( n7269 , n7261 , n7268 );
buf ( n7270 , n4587 );
xor ( n7271 , n7269 , n7270 );
buf ( n7272 , n4588 );
xor ( n7273 , n7271 , n7272 );
xor ( n7274 , n7273 , n7137 );
xor ( n7275 , n7254 , n7274 );
not ( n7276 , n7275 );
not ( n7277 , n6474 );
buf ( n7278 , n4589 );
and ( n7279 , n7277 , n7278 );
buf ( n7280 , n4590 );
xor ( n7281 , n7280 , n7278 );
and ( n7282 , n7281 , n6474 );
or ( n7283 , n7279 , n7282 );
xor ( n7284 , n7283 , n6717 );
xor ( n7285 , n7284 , n6739 );
and ( n7286 , n7276 , n7285 );
xor ( n7287 , n7231 , n7286 );
buf ( n7288 , n4591 );
not ( n7289 , n6474 );
buf ( n7290 , n4592 );
and ( n7291 , n7289 , n7290 );
buf ( n7292 , n4593 );
xor ( n7293 , n7292 , n7290 );
and ( n7294 , n7293 , n6474 );
or ( n7295 , n7291 , n7294 );
not ( n7296 , n6474 );
buf ( n7297 , n4594 );
and ( n7298 , n7296 , n7297 );
buf ( n7299 , n4595 );
xor ( n7300 , n7299 , n7297 );
and ( n7301 , n7300 , n6474 );
or ( n7302 , n7298 , n7301 );
xor ( n7303 , n7295 , n7302 );
buf ( n7304 , n4596 );
xor ( n7305 , n7303 , n7304 );
buf ( n7306 , n4597 );
xor ( n7307 , n7305 , n7306 );
buf ( n7308 , n4598 );
xor ( n7309 , n7307 , n7308 );
xor ( n7310 , n7288 , n7309 );
not ( n7311 , n6474 );
buf ( n7312 , n4599 );
and ( n7313 , n7311 , n7312 );
buf ( n7314 , n4600 );
xor ( n7315 , n7314 , n7312 );
and ( n7316 , n7315 , n6474 );
or ( n7317 , n7313 , n7316 );
not ( n7318 , n6474 );
buf ( n7319 , n4601 );
and ( n7320 , n7318 , n7319 );
buf ( n7321 , n4602 );
xor ( n7322 , n7321 , n7319 );
and ( n7323 , n7322 , n6474 );
or ( n7324 , n7320 , n7323 );
xor ( n7325 , n7317 , n7324 );
buf ( n7326 , n4603 );
xor ( n7327 , n7325 , n7326 );
buf ( n7328 , n4604 );
xor ( n7329 , n7327 , n7328 );
buf ( n7330 , n4605 );
xor ( n7331 , n7329 , n7330 );
xor ( n7332 , n7310 , n7331 );
not ( n7333 , n6474 );
buf ( n7334 , n4606 );
and ( n7335 , n7333 , n7334 );
buf ( n7336 , n4607 );
xor ( n7337 , n7336 , n7334 );
and ( n7338 , n7337 , n6474 );
or ( n7339 , n7335 , n7338 );
not ( n7340 , n6474 );
buf ( n7341 , n4608 );
and ( n7342 , n7340 , n7341 );
buf ( n7343 , n4609 );
xor ( n7344 , n7343 , n7341 );
and ( n7345 , n7344 , n6474 );
or ( n7346 , n7342 , n7345 );
not ( n7347 , n6474 );
buf ( n7348 , n4610 );
and ( n7349 , n7347 , n7348 );
buf ( n7350 , n4611 );
xor ( n7351 , n7350 , n7348 );
and ( n7352 , n7351 , n6474 );
or ( n7353 , n7349 , n7352 );
xor ( n7354 , n7346 , n7353 );
buf ( n7355 , n4612 );
xor ( n7356 , n7354 , n7355 );
buf ( n7357 , n4613 );
xor ( n7358 , n7356 , n7357 );
buf ( n7359 , n4614 );
xor ( n7360 , n7358 , n7359 );
xor ( n7361 , n7339 , n7360 );
not ( n7362 , n6474 );
buf ( n7363 , n4615 );
and ( n7364 , n7362 , n7363 );
buf ( n7365 , n4616 );
xor ( n7366 , n7365 , n7363 );
and ( n7367 , n7366 , n6474 );
or ( n7368 , n7364 , n7367 );
buf ( n7369 , n4617 );
xor ( n7370 , n7368 , n7369 );
buf ( n7371 , n4618 );
xor ( n7372 , n7370 , n7371 );
buf ( n7373 , n4619 );
xor ( n7374 , n7372 , n7373 );
buf ( n7375 , n4620 );
xor ( n7376 , n7374 , n7375 );
xor ( n7377 , n7361 , n7376 );
not ( n7378 , n7377 );
buf ( n7379 , n4621 );
not ( n7380 , n6474 );
buf ( n7381 , n4622 );
and ( n7382 , n7380 , n7381 );
buf ( n7383 , n4623 );
xor ( n7384 , n7383 , n7381 );
and ( n7385 , n7384 , n6474 );
or ( n7386 , n7382 , n7385 );
not ( n7387 , n6474 );
buf ( n7388 , n4624 );
and ( n7389 , n7387 , n7388 );
buf ( n7390 , n4625 );
xor ( n7391 , n7390 , n7388 );
and ( n7392 , n7391 , n6474 );
or ( n7393 , n7389 , n7392 );
xor ( n7394 , n7386 , n7393 );
buf ( n7395 , n4626 );
xor ( n7396 , n7394 , n7395 );
xor ( n7397 , n7396 , n6479 );
buf ( n7398 , n4627 );
xor ( n7399 , n7397 , n7398 );
xor ( n7400 , n7379 , n7399 );
not ( n7401 , n6474 );
buf ( n7402 , n4628 );
and ( n7403 , n7401 , n7402 );
buf ( n7404 , n4629 );
xor ( n7405 , n7404 , n7402 );
and ( n7406 , n7405 , n6474 );
or ( n7407 , n7403 , n7406 );
not ( n7408 , n6474 );
buf ( n7409 , n4630 );
and ( n7410 , n7408 , n7409 );
buf ( n7411 , n4631 );
xor ( n7412 , n7411 , n7409 );
and ( n7413 , n7412 , n6474 );
or ( n7414 , n7410 , n7413 );
xor ( n7415 , n7407 , n7414 );
buf ( n7416 , n4632 );
xor ( n7417 , n7415 , n7416 );
buf ( n7418 , n4633 );
xor ( n7419 , n7417 , n7418 );
buf ( n7420 , n4634 );
xor ( n7421 , n7419 , n7420 );
xor ( n7422 , n7400 , n7421 );
and ( n7423 , n7378 , n7422 );
xor ( n7424 , n7332 , n7423 );
xor ( n7425 , n7287 , n7424 );
buf ( n7426 , n4635 );
not ( n7427 , n6474 );
buf ( n7428 , n4636 );
and ( n7429 , n7427 , n7428 );
buf ( n7430 , n4637 );
xor ( n7431 , n7430 , n7428 );
and ( n7432 , n7431 , n6474 );
or ( n7433 , n7429 , n7432 );
buf ( n7434 , n4638 );
xor ( n7435 , n7433 , n7434 );
buf ( n7436 , n4639 );
xor ( n7437 , n7435 , n7436 );
buf ( n7438 , n4640 );
xor ( n7439 , n7437 , n7438 );
buf ( n7440 , n4641 );
xor ( n7441 , n7439 , n7440 );
xor ( n7442 , n7426 , n7441 );
not ( n7443 , n6474 );
buf ( n7444 , n4642 );
and ( n7445 , n7443 , n7444 );
buf ( n7446 , n4643 );
xor ( n7447 , n7446 , n7444 );
and ( n7448 , n7447 , n6474 );
or ( n7449 , n7445 , n7448 );
not ( n7450 , n6474 );
buf ( n7451 , n4644 );
and ( n7452 , n7450 , n7451 );
buf ( n7453 , n4645 );
xor ( n7454 , n7453 , n7451 );
and ( n7455 , n7454 , n6474 );
or ( n7456 , n7452 , n7455 );
xor ( n7457 , n7449 , n7456 );
buf ( n7458 , n4646 );
xor ( n7459 , n7457 , n7458 );
buf ( n7460 , n4647 );
xor ( n7461 , n7459 , n7460 );
buf ( n7462 , n4648 );
xor ( n7463 , n7461 , n7462 );
xor ( n7464 , n7442 , n7463 );
xor ( n7465 , n7261 , n7159 );
xor ( n7466 , n7465 , n7181 );
not ( n7467 , n7466 );
not ( n7468 , n6474 );
buf ( n7469 , n4649 );
and ( n7470 , n7468 , n7469 );
buf ( n7471 , n4650 );
xor ( n7472 , n7471 , n7469 );
and ( n7473 , n7472 , n6474 );
or ( n7474 , n7470 , n7473 );
not ( n7475 , n6474 );
buf ( n7476 , n7475 );
buf ( n7477 , n4651 );
not ( n7478 , n7477 );
and ( n7479 , n7478 , n6474 );
or ( n7480 , n7476 , n7479 );
not ( n7481 , n6474 );
buf ( n7482 , n4652 );
and ( n7483 , n7481 , n7482 );
buf ( n7484 , n4653 );
xor ( n7485 , n7484 , n7482 );
and ( n7486 , n7485 , n6474 );
or ( n7487 , n7483 , n7486 );
xor ( n7488 , n7480 , n7487 );
buf ( n7489 , n4654 );
xor ( n7490 , n7488 , n7489 );
buf ( n7491 , n4655 );
xor ( n7492 , n7490 , n7491 );
buf ( n7493 , n4656 );
xor ( n7494 , n7492 , n7493 );
xor ( n7495 , n7474 , n7494 );
xor ( n7496 , n7495 , n6850 );
and ( n7497 , n7467 , n7496 );
xor ( n7498 , n7464 , n7497 );
xor ( n7499 , n7425 , n7498 );
buf ( n7500 , n4657 );
not ( n7501 , n6474 );
buf ( n7502 , n4658 );
and ( n7503 , n7501 , n7502 );
buf ( n7504 , n4659 );
xor ( n7505 , n7504 , n7502 );
and ( n7506 , n7505 , n6474 );
or ( n7507 , n7503 , n7506 );
not ( n7508 , n6474 );
buf ( n7509 , n4660 );
and ( n7510 , n7508 , n7509 );
buf ( n7511 , n4661 );
xor ( n7512 , n7511 , n7509 );
and ( n7513 , n7512 , n6474 );
or ( n7514 , n7510 , n7513 );
xor ( n7515 , n7507 , n7514 );
buf ( n7516 , n4662 );
xor ( n7517 , n7515 , n7516 );
buf ( n7518 , n4663 );
xor ( n7519 , n7517 , n7518 );
buf ( n7520 , n4664 );
xor ( n7521 , n7519 , n7520 );
xor ( n7522 , n7500 , n7521 );
not ( n7523 , n6474 );
buf ( n7524 , n4665 );
and ( n7525 , n7523 , n7524 );
buf ( n7526 , n4666 );
xor ( n7527 , n7526 , n7524 );
and ( n7528 , n7527 , n6474 );
or ( n7529 , n7525 , n7528 );
buf ( n7530 , n4667 );
xor ( n7531 , n7529 , n7530 );
buf ( n7532 , n4668 );
xor ( n7533 , n7531 , n7532 );
buf ( n7534 , n4669 );
xor ( n7535 , n7533 , n7534 );
buf ( n7536 , n4670 );
xor ( n7537 , n7535 , n7536 );
xor ( n7538 , n7522 , n7537 );
not ( n7539 , n6474 );
buf ( n7540 , n4671 );
and ( n7541 , n7539 , n7540 );
buf ( n7542 , n4672 );
xor ( n7543 , n7542 , n7540 );
and ( n7544 , n7543 , n6474 );
or ( n7545 , n7541 , n7544 );
not ( n7546 , n6474 );
buf ( n7547 , n4673 );
and ( n7548 , n7546 , n7547 );
buf ( n7549 , n4674 );
xor ( n7550 , n7549 , n7547 );
and ( n7551 , n7550 , n6474 );
or ( n7552 , n7548 , n7551 );
not ( n7553 , n6474 );
buf ( n7554 , n4675 );
and ( n7555 , n7553 , n7554 );
buf ( n7556 , n4676 );
xor ( n7557 , n7556 , n7554 );
and ( n7558 , n7557 , n6474 );
or ( n7559 , n7555 , n7558 );
xor ( n7560 , n7552 , n7559 );
buf ( n7561 , n4677 );
xor ( n7562 , n7560 , n7561 );
buf ( n7563 , n4678 );
xor ( n7564 , n7562 , n7563 );
buf ( n7565 , n4679 );
xor ( n7566 , n7564 , n7565 );
xor ( n7567 , n7545 , n7566 );
not ( n7568 , n6474 );
buf ( n7569 , n4680 );
and ( n7570 , n7568 , n7569 );
buf ( n7571 , n4681 );
xor ( n7572 , n7571 , n7569 );
and ( n7573 , n7572 , n6474 );
or ( n7574 , n7570 , n7573 );
not ( n7575 , n6474 );
buf ( n7576 , n4682 );
and ( n7577 , n7575 , n7576 );
buf ( n7578 , n4683 );
xor ( n7579 , n7578 , n7576 );
and ( n7580 , n7579 , n6474 );
or ( n7581 , n7577 , n7580 );
xor ( n7582 , n7574 , n7581 );
buf ( n7583 , n4684 );
xor ( n7584 , n7582 , n7583 );
buf ( n7585 , n4685 );
xor ( n7586 , n7584 , n7585 );
buf ( n7587 , n4686 );
xor ( n7588 , n7586 , n7587 );
xor ( n7589 , n7567 , n7588 );
not ( n7590 , n7589 );
not ( n7591 , n6474 );
buf ( n7592 , n4687 );
and ( n7593 , n7591 , n7592 );
buf ( n7594 , n4688 );
xor ( n7595 , n7594 , n7592 );
and ( n7596 , n7595 , n6474 );
or ( n7597 , n7593 , n7596 );
not ( n7598 , n6474 );
buf ( n7599 , n4689 );
and ( n7600 , n7598 , n7599 );
buf ( n7601 , n4690 );
xor ( n7602 , n7601 , n7599 );
and ( n7603 , n7602 , n6474 );
or ( n7604 , n7600 , n7603 );
buf ( n7605 , n4691 );
xor ( n7606 , n7604 , n7605 );
buf ( n7607 , n4692 );
xor ( n7608 , n7606 , n7607 );
buf ( n7609 , n4693 );
xor ( n7610 , n7608 , n7609 );
buf ( n7611 , n4694 );
xor ( n7612 , n7610 , n7611 );
xor ( n7613 , n7597 , n7612 );
not ( n7614 , n6474 );
buf ( n7615 , n4695 );
and ( n7616 , n7614 , n7615 );
buf ( n7617 , n4696 );
xor ( n7618 , n7617 , n7615 );
and ( n7619 , n7618 , n6474 );
or ( n7620 , n7616 , n7619 );
not ( n7621 , n6474 );
buf ( n7622 , n4697 );
and ( n7623 , n7621 , n7622 );
buf ( n7624 , n4698 );
xor ( n7625 , n7624 , n7622 );
and ( n7626 , n7625 , n6474 );
or ( n7627 , n7623 , n7626 );
xor ( n7628 , n7620 , n7627 );
buf ( n7629 , n4699 );
xor ( n7630 , n7628 , n7629 );
buf ( n7631 , n4700 );
xor ( n7632 , n7630 , n7631 );
buf ( n7633 , n4701 );
xor ( n7634 , n7632 , n7633 );
xor ( n7635 , n7613 , n7634 );
and ( n7636 , n7590 , n7635 );
xor ( n7637 , n7538 , n7636 );
xor ( n7638 , n7499 , n7637 );
buf ( n7639 , n4702 );
not ( n7640 , n6474 );
buf ( n7641 , n4703 );
and ( n7642 , n7640 , n7641 );
buf ( n7643 , n4704 );
xor ( n7644 , n7643 , n7641 );
and ( n7645 , n7644 , n6474 );
or ( n7646 , n7642 , n7645 );
not ( n7647 , n6474 );
buf ( n7648 , n4705 );
and ( n7649 , n7647 , n7648 );
buf ( n7650 , n4706 );
xor ( n7651 , n7650 , n7648 );
and ( n7652 , n7651 , n6474 );
or ( n7653 , n7649 , n7652 );
xor ( n7654 , n7646 , n7653 );
xor ( n7655 , n7654 , n6658 );
buf ( n7656 , n4707 );
xor ( n7657 , n7655 , n7656 );
buf ( n7658 , n4708 );
xor ( n7659 , n7657 , n7658 );
xor ( n7660 , n7639 , n7659 );
not ( n7661 , n6474 );
buf ( n7662 , n4709 );
and ( n7663 , n7661 , n7662 );
buf ( n7664 , n4710 );
xor ( n7665 , n7664 , n7662 );
and ( n7666 , n7665 , n6474 );
or ( n7667 , n7663 , n7666 );
not ( n7668 , n6474 );
buf ( n7669 , n4711 );
and ( n7670 , n7668 , n7669 );
buf ( n7671 , n4712 );
xor ( n7672 , n7671 , n7669 );
and ( n7673 , n7672 , n6474 );
or ( n7674 , n7670 , n7673 );
xor ( n7675 , n7667 , n7674 );
buf ( n7676 , n4713 );
xor ( n7677 , n7675 , n7676 );
buf ( n7678 , n4714 );
xor ( n7679 , n7677 , n7678 );
buf ( n7680 , n4715 );
xor ( n7681 , n7679 , n7680 );
xor ( n7682 , n7660 , n7681 );
not ( n7683 , n6474 );
buf ( n7684 , n4716 );
and ( n7685 , n7683 , n7684 );
buf ( n7686 , n4717 );
xor ( n7687 , n7686 , n7684 );
and ( n7688 , n7687 , n6474 );
or ( n7689 , n7685 , n7688 );
not ( n7690 , n6474 );
buf ( n7691 , n4718 );
and ( n7692 , n7690 , n7691 );
buf ( n7693 , n4719 );
xor ( n7694 , n7693 , n7691 );
and ( n7695 , n7694 , n6474 );
or ( n7696 , n7692 , n7695 );
not ( n7697 , n6474 );
buf ( n7698 , n4720 );
and ( n7699 , n7697 , n7698 );
buf ( n7700 , n4721 );
xor ( n7701 , n7700 , n7698 );
and ( n7702 , n7701 , n6474 );
or ( n7703 , n7699 , n7702 );
xor ( n7704 , n7696 , n7703 );
buf ( n7705 , n4722 );
xor ( n7706 , n7704 , n7705 );
buf ( n7707 , n4723 );
xor ( n7708 , n7706 , n7707 );
buf ( n7709 , n4724 );
xor ( n7710 , n7708 , n7709 );
xor ( n7711 , n7689 , n7710 );
not ( n7712 , n6474 );
buf ( n7713 , n4725 );
and ( n7714 , n7712 , n7713 );
buf ( n7715 , n4726 );
xor ( n7716 , n7715 , n7713 );
and ( n7717 , n7716 , n6474 );
or ( n7718 , n7714 , n7717 );
not ( n7719 , n6474 );
buf ( n7720 , n4727 );
and ( n7721 , n7719 , n7720 );
buf ( n7722 , n4728 );
xor ( n7723 , n7722 , n7720 );
and ( n7724 , n7723 , n6474 );
or ( n7725 , n7721 , n7724 );
xor ( n7726 , n7718 , n7725 );
buf ( n7727 , n4729 );
xor ( n7728 , n7726 , n7727 );
buf ( n7729 , n4730 );
xor ( n7730 , n7728 , n7729 );
buf ( n7731 , n4731 );
xor ( n7732 , n7730 , n7731 );
xor ( n7733 , n7711 , n7732 );
not ( n7734 , n7733 );
not ( n7735 , n6474 );
buf ( n7736 , n4732 );
and ( n7737 , n7735 , n7736 );
buf ( n7738 , n4733 );
xor ( n7739 , n7738 , n7736 );
and ( n7740 , n7739 , n6474 );
or ( n7741 , n7737 , n7740 );
xor ( n7742 , n7741 , n7030 );
xor ( n7743 , n7742 , n7046 );
and ( n7744 , n7734 , n7743 );
xor ( n7745 , n7682 , n7744 );
xor ( n7746 , n7638 , n7745 );
xor ( n7747 , n7186 , n7746 );
buf ( n7748 , n4734 );
not ( n7749 , n6474 );
buf ( n7750 , n4735 );
and ( n7751 , n7749 , n7750 );
buf ( n7752 , n4736 );
xor ( n7753 , n7752 , n7750 );
and ( n7754 , n7753 , n6474 );
or ( n7755 , n7751 , n7754 );
not ( n7756 , n6474 );
buf ( n7757 , n4737 );
and ( n7758 , n7756 , n7757 );
buf ( n7759 , n4738 );
xor ( n7760 , n7759 , n7757 );
and ( n7761 , n7760 , n6474 );
or ( n7762 , n7758 , n7761 );
xor ( n7763 , n7755 , n7762 );
buf ( n7764 , n4739 );
xor ( n7765 , n7763 , n7764 );
not ( n7766 , n4740 );
buf ( n7767 , n7766 );
buf ( n7768 , n7767 );
xor ( n7769 , n7765 , n7768 );
buf ( n7770 , n4741 );
xor ( n7771 , n7769 , n7770 );
xor ( n7772 , n7748 , n7771 );
not ( n7773 , n6474 );
buf ( n7774 , n4742 );
and ( n7775 , n7773 , n7774 );
buf ( n7776 , n4743 );
xor ( n7777 , n7776 , n7774 );
and ( n7778 , n7777 , n6474 );
or ( n7779 , n7775 , n7778 );
not ( n7780 , n6474 );
buf ( n7781 , n4744 );
and ( n7782 , n7780 , n7781 );
buf ( n7783 , n4745 );
xor ( n7784 , n7783 , n7781 );
and ( n7785 , n7784 , n6474 );
or ( n7786 , n7782 , n7785 );
xor ( n7787 , n7779 , n7786 );
buf ( n7788 , n4746 );
xor ( n7789 , n7787 , n7788 );
buf ( n7790 , n4747 );
xor ( n7791 , n7789 , n7790 );
buf ( n7792 , n4748 );
xor ( n7793 , n7791 , n7792 );
xor ( n7794 , n7772 , n7793 );
not ( n7795 , n6474 );
buf ( n7796 , n4749 );
and ( n7797 , n7795 , n7796 );
buf ( n7798 , n4750 );
xor ( n7799 , n7798 , n7796 );
and ( n7800 , n7799 , n6474 );
or ( n7801 , n7797 , n7800 );
not ( n7802 , n6474 );
buf ( n7803 , n4751 );
and ( n7804 , n7802 , n7803 );
buf ( n7805 , n4752 );
xor ( n7806 , n7805 , n7803 );
and ( n7807 , n7806 , n6474 );
or ( n7808 , n7804 , n7807 );
not ( n7809 , n6474 );
buf ( n7810 , n4753 );
and ( n7811 , n7809 , n7810 );
buf ( n7812 , n4754 );
xor ( n7813 , n7812 , n7810 );
and ( n7814 , n7813 , n6474 );
or ( n7815 , n7811 , n7814 );
xor ( n7816 , n7808 , n7815 );
buf ( n7817 , n4755 );
xor ( n7818 , n7816 , n7817 );
buf ( n7819 , n4756 );
xor ( n7820 , n7818 , n7819 );
buf ( n7821 , n4757 );
xor ( n7822 , n7820 , n7821 );
xor ( n7823 , n7801 , n7822 );
not ( n7824 , n6474 );
buf ( n7825 , n4758 );
and ( n7826 , n7824 , n7825 );
buf ( n7827 , n4759 );
xor ( n7828 , n7827 , n7825 );
and ( n7829 , n7828 , n6474 );
or ( n7830 , n7826 , n7829 );
xor ( n7831 , n7830 , n7379 );
buf ( n7832 , n4760 );
xor ( n7833 , n7831 , n7832 );
buf ( n7834 , n4761 );
xor ( n7835 , n7833 , n7834 );
buf ( n7836 , n4762 );
xor ( n7837 , n7835 , n7836 );
xor ( n7838 , n7823 , n7837 );
not ( n7839 , n7838 );
buf ( n7840 , n4763 );
not ( n7841 , n6474 );
buf ( n7842 , n4764 );
and ( n7843 , n7841 , n7842 );
buf ( n7844 , n4765 );
xor ( n7845 , n7844 , n7842 );
and ( n7846 , n7845 , n6474 );
or ( n7847 , n7843 , n7846 );
not ( n7848 , n6474 );
buf ( n7849 , n4766 );
and ( n7850 , n7848 , n7849 );
buf ( n7851 , n4767 );
xor ( n7852 , n7851 , n7849 );
and ( n7853 , n7852 , n6474 );
or ( n7854 , n7850 , n7853 );
xor ( n7855 , n7847 , n7854 );
buf ( n7856 , n4768 );
xor ( n7857 , n7855 , n7856 );
buf ( n7858 , n4769 );
xor ( n7859 , n7857 , n7858 );
buf ( n7860 , n4770 );
xor ( n7861 , n7859 , n7860 );
xor ( n7862 , n7840 , n7861 );
not ( n7863 , n6474 );
buf ( n7864 , n4771 );
and ( n7865 , n7863 , n7864 );
buf ( n7866 , n4772 );
xor ( n7867 , n7866 , n7864 );
and ( n7868 , n7867 , n6474 );
or ( n7869 , n7865 , n7868 );
not ( n7870 , n6474 );
buf ( n7871 , n4773 );
and ( n7872 , n7870 , n7871 );
buf ( n7873 , n4774 );
xor ( n7874 , n7873 , n7871 );
and ( n7875 , n7874 , n6474 );
or ( n7876 , n7872 , n7875 );
xor ( n7877 , n7869 , n7876 );
buf ( n7878 , n4775 );
xor ( n7879 , n7877 , n7878 );
buf ( n7880 , n4776 );
xor ( n7881 , n7879 , n7880 );
buf ( n7882 , n4777 );
xor ( n7883 , n7881 , n7882 );
xor ( n7884 , n7862 , n7883 );
and ( n7885 , n7839 , n7884 );
xor ( n7886 , n7794 , n7885 );
not ( n7887 , n4780 );
buf ( n7888 , n7887 );
buf ( n7889 , n7888 );
not ( n7890 , n6474 );
buf ( n7891 , n4778 );
and ( n7892 , n7890 , n7891 );
buf ( n7893 , n4779 );
xor ( n7894 , n7893 , n7891 );
and ( n7895 , n7894 , n6474 );
or ( n7896 , n7892 , n7895 );
not ( n7897 , n6474 );
buf ( n7898 , n4780 );
and ( n7899 , n7897 , n7898 );
buf ( n7900 , n4781 );
xor ( n7901 , n7900 , n7898 );
and ( n7902 , n7901 , n6474 );
or ( n7903 , n7899 , n7902 );
xor ( n7904 , n7896 , n7903 );
buf ( n7905 , n4782 );
xor ( n7906 , n7904 , n7905 );
buf ( n7907 , n4783 );
xor ( n7908 , n7906 , n7907 );
buf ( n7909 , n4784 );
xor ( n7910 , n7908 , n7909 );
xor ( n7911 , n7889 , n7910 );
not ( n7912 , n6474 );
buf ( n7913 , n4785 );
and ( n7914 , n7912 , n7913 );
buf ( n7915 , n4786 );
xor ( n7916 , n7915 , n7913 );
and ( n7917 , n7916 , n6474 );
or ( n7918 , n7914 , n7917 );
buf ( n7919 , n4787 );
xor ( n7920 , n7918 , n7919 );
buf ( n7921 , n4788 );
xor ( n7922 , n7920 , n7921 );
buf ( n7923 , n4789 );
xor ( n7924 , n7922 , n7923 );
xor ( n7925 , n7924 , n6518 );
xor ( n7926 , n7911 , n7925 );
buf ( n7927 , n4790 );
not ( n7928 , n6474 );
buf ( n7929 , n4791 );
and ( n7930 , n7928 , n7929 );
buf ( n7931 , n4792 );
xor ( n7932 , n7931 , n7929 );
and ( n7933 , n7932 , n6474 );
or ( n7934 , n7930 , n7933 );
not ( n7935 , n6474 );
buf ( n7936 , n4793 );
and ( n7937 , n7935 , n7936 );
buf ( n7938 , n4794 );
xor ( n7939 , n7938 , n7936 );
and ( n7940 , n7939 , n6474 );
or ( n7941 , n7937 , n7940 );
xor ( n7942 , n7934 , n7941 );
buf ( n7943 , n4795 );
xor ( n7944 , n7942 , n7943 );
buf ( n7945 , n4796 );
xor ( n7946 , n7944 , n7945 );
buf ( n7947 , n4797 );
xor ( n7948 , n7946 , n7947 );
xor ( n7949 , n7927 , n7948 );
not ( n7950 , n6474 );
buf ( n7951 , n4798 );
and ( n7952 , n7950 , n7951 );
buf ( n7953 , n4799 );
xor ( n7954 , n7953 , n7951 );
and ( n7955 , n7954 , n6474 );
or ( n7956 , n7952 , n7955 );
not ( n7957 , n6474 );
buf ( n7958 , n4800 );
and ( n7959 , n7957 , n7958 );
buf ( n7960 , n4801 );
xor ( n7961 , n7960 , n7958 );
and ( n7962 , n7961 , n6474 );
or ( n7963 , n7959 , n7962 );
xor ( n7964 , n7956 , n7963 );
buf ( n7965 , n4802 );
xor ( n7966 , n7964 , n7965 );
buf ( n7967 , n4803 );
xor ( n7968 , n7966 , n7967 );
buf ( n7969 , n4804 );
xor ( n7970 , n7968 , n7969 );
xor ( n7971 , n7949 , n7970 );
not ( n7972 , n7971 );
not ( n7973 , n6474 );
buf ( n7974 , n4805 );
and ( n7975 , n7973 , n7974 );
buf ( n7976 , n4806 );
xor ( n7977 , n7976 , n7974 );
and ( n7978 , n7977 , n6474 );
or ( n7979 , n7975 , n7978 );
not ( n7980 , n6474 );
buf ( n7981 , n4807 );
and ( n7982 , n7980 , n7981 );
buf ( n7983 , n4808 );
xor ( n7984 , n7983 , n7981 );
and ( n7985 , n7984 , n6474 );
or ( n7986 , n7982 , n7985 );
buf ( n7987 , n4809 );
xor ( n7988 , n7986 , n7987 );
buf ( n7989 , n4810 );
xor ( n7990 , n7988 , n7989 );
buf ( n7991 , n4811 );
xor ( n7992 , n7990 , n7991 );
buf ( n7993 , n4812 );
xor ( n7994 , n7992 , n7993 );
xor ( n7995 , n7979 , n7994 );
not ( n7996 , n6474 );
buf ( n7997 , n4813 );
and ( n7998 , n7996 , n7997 );
buf ( n7999 , n4814 );
xor ( n8000 , n7999 , n7997 );
and ( n8001 , n8000 , n6474 );
or ( n8002 , n7998 , n8001 );
not ( n8003 , n6474 );
buf ( n8004 , n4815 );
and ( n8005 , n8003 , n8004 );
buf ( n8006 , n4816 );
xor ( n8007 , n8006 , n8004 );
and ( n8008 , n8007 , n6474 );
or ( n8009 , n8005 , n8008 );
xor ( n8010 , n8002 , n8009 );
buf ( n8011 , n4817 );
xor ( n8012 , n8010 , n8011 );
buf ( n8013 , n4818 );
xor ( n8014 , n8012 , n8013 );
buf ( n8015 , n4819 );
xor ( n8016 , n8014 , n8015 );
xor ( n8017 , n7995 , n8016 );
and ( n8018 , n7972 , n8017 );
xor ( n8019 , n7926 , n8018 );
buf ( n8020 , n4820 );
not ( n8021 , n6474 );
buf ( n8022 , n4821 );
and ( n8023 , n8021 , n8022 );
buf ( n8024 , n4822 );
xor ( n8025 , n8024 , n8022 );
and ( n8026 , n8025 , n6474 );
or ( n8027 , n8023 , n8026 );
xor ( n8028 , n8027 , n7597 );
buf ( n8029 , n4823 );
xor ( n8030 , n8028 , n8029 );
buf ( n8031 , n4824 );
xor ( n8032 , n8030 , n8031 );
buf ( n8033 , n4825 );
xor ( n8034 , n8032 , n8033 );
xor ( n8035 , n8020 , n8034 );
not ( n8036 , n6474 );
buf ( n8037 , n4826 );
and ( n8038 , n8036 , n8037 );
buf ( n8039 , n4827 );
xor ( n8040 , n8039 , n8037 );
and ( n8041 , n8040 , n6474 );
or ( n8042 , n8038 , n8041 );
not ( n8043 , n6474 );
buf ( n8044 , n4828 );
and ( n8045 , n8043 , n8044 );
buf ( n8046 , n4829 );
xor ( n8047 , n8046 , n8044 );
and ( n8048 , n8047 , n6474 );
or ( n8049 , n8045 , n8048 );
xor ( n8050 , n8042 , n8049 );
buf ( n8051 , n4830 );
xor ( n8052 , n8050 , n8051 );
buf ( n8053 , n4831 );
xor ( n8054 , n8052 , n8053 );
buf ( n8055 , n4832 );
xor ( n8056 , n8054 , n8055 );
xor ( n8057 , n8035 , n8056 );
not ( n8058 , n7794 );
and ( n8059 , n8058 , n7838 );
xor ( n8060 , n8057 , n8059 );
xor ( n8061 , n8019 , n8060 );
xor ( n8062 , n6581 , n7732 );
not ( n8063 , n6474 );
buf ( n8064 , n4833 );
and ( n8065 , n8063 , n8064 );
buf ( n8066 , n4834 );
xor ( n8067 , n8066 , n8064 );
and ( n8068 , n8067 , n6474 );
or ( n8069 , n8065 , n8068 );
xor ( n8070 , n7238 , n8069 );
buf ( n8071 , n4835 );
xor ( n8072 , n8070 , n8071 );
buf ( n8073 , n4836 );
xor ( n8074 , n8072 , n8073 );
buf ( n8075 , n4837 );
xor ( n8076 , n8074 , n8075 );
xor ( n8077 , n8062 , n8076 );
not ( n8078 , n6474 );
buf ( n8079 , n4838 );
and ( n8080 , n8078 , n8079 );
buf ( n8081 , n4839 );
xor ( n8082 , n8081 , n8079 );
and ( n8083 , n8082 , n6474 );
or ( n8084 , n8080 , n8083 );
buf ( n8085 , n4840 );
xor ( n8086 , n8084 , n8085 );
buf ( n8087 , n4841 );
xor ( n8088 , n8086 , n8087 );
buf ( n8089 , n4842 );
xor ( n8090 , n8088 , n8089 );
buf ( n8091 , n4843 );
xor ( n8092 , n8090 , n8091 );
xor ( n8093 , n6938 , n8092 );
not ( n8094 , n6474 );
buf ( n8095 , n4844 );
and ( n8096 , n8094 , n8095 );
buf ( n8097 , n4845 );
xor ( n8098 , n8097 , n8095 );
and ( n8099 , n8098 , n6474 );
or ( n8100 , n8096 , n8099 );
not ( n8101 , n6474 );
buf ( n8102 , n4846 );
and ( n8103 , n8101 , n8102 );
buf ( n8104 , n4847 );
xor ( n8105 , n8104 , n8102 );
and ( n8106 , n8105 , n6474 );
or ( n8107 , n8103 , n8106 );
xor ( n8108 , n8100 , n8107 );
buf ( n8109 , n4848 );
xor ( n8110 , n8108 , n8109 );
buf ( n8111 , n4849 );
xor ( n8112 , n8110 , n8111 );
buf ( n8113 , n4850 );
xor ( n8114 , n8112 , n8113 );
xor ( n8115 , n8093 , n8114 );
not ( n8116 , n8115 );
not ( n8117 , n6474 );
buf ( n8118 , n4851 );
and ( n8119 , n8117 , n8118 );
buf ( n8120 , n4852 );
xor ( n8121 , n8120 , n8118 );
and ( n8122 , n8121 , n6474 );
or ( n8123 , n8119 , n8122 );
not ( n8124 , n6474 );
buf ( n8125 , n4853 );
and ( n8126 , n8124 , n8125 );
buf ( n8127 , n4854 );
xor ( n8128 , n8127 , n8125 );
and ( n8129 , n8128 , n6474 );
or ( n8130 , n8126 , n8129 );
xor ( n8131 , n8123 , n8130 );
buf ( n8132 , n4855 );
xor ( n8133 , n8131 , n8132 );
buf ( n8134 , n4856 );
xor ( n8135 , n8133 , n8134 );
buf ( n8136 , n4857 );
xor ( n8137 , n8135 , n8136 );
xor ( n8138 , n8002 , n8137 );
not ( n8139 , n6474 );
buf ( n8140 , n4858 );
and ( n8141 , n8139 , n8140 );
buf ( n8142 , n4859 );
xor ( n8143 , n8142 , n8140 );
and ( n8144 , n8143 , n6474 );
or ( n8145 , n8141 , n8144 );
not ( n8146 , n6474 );
buf ( n8147 , n4860 );
and ( n8148 , n8146 , n8147 );
buf ( n8149 , n4861 );
xor ( n8150 , n8149 , n8147 );
and ( n8151 , n8150 , n6474 );
or ( n8152 , n8148 , n8151 );
xor ( n8153 , n8145 , n8152 );
buf ( n8154 , n4862 );
xor ( n8155 , n8153 , n8154 );
buf ( n8156 , n4863 );
xor ( n8157 , n8155 , n8156 );
buf ( n8158 , n4864 );
xor ( n8159 , n8157 , n8158 );
xor ( n8160 , n8138 , n8159 );
and ( n8161 , n8116 , n8160 );
xor ( n8162 , n8077 , n8161 );
xor ( n8163 , n8061 , n8162 );
buf ( n8164 , n4865 );
xor ( n8165 , n8164 , n7494 );
xor ( n8166 , n8165 , n6850 );
buf ( n8167 , n4866 );
not ( n8168 , n6474 );
buf ( n8169 , n4867 );
and ( n8170 , n8168 , n8169 );
buf ( n8171 , n4868 );
xor ( n8172 , n8171 , n8169 );
and ( n8173 , n8172 , n6474 );
or ( n8174 , n8170 , n8173 );
not ( n8175 , n6474 );
buf ( n8176 , n4869 );
and ( n8177 , n8175 , n8176 );
buf ( n8178 , n4870 );
xor ( n8179 , n8178 , n8176 );
and ( n8180 , n8179 , n6474 );
or ( n8181 , n8177 , n8180 );
xor ( n8182 , n8174 , n8181 );
buf ( n8183 , n4871 );
xor ( n8184 , n8182 , n8183 );
buf ( n8185 , n4872 );
xor ( n8186 , n8184 , n8185 );
buf ( n8187 , n4873 );
xor ( n8188 , n8186 , n8187 );
xor ( n8189 , n8167 , n8188 );
not ( n8190 , n6474 );
buf ( n8191 , n4874 );
and ( n8192 , n8190 , n8191 );
buf ( n8193 , n4875 );
xor ( n8194 , n8193 , n8191 );
and ( n8195 , n8194 , n6474 );
or ( n8196 , n8192 , n8195 );
buf ( n8197 , n4876 );
xor ( n8198 , n8196 , n8197 );
buf ( n8199 , n4877 );
xor ( n8200 , n8198 , n8199 );
buf ( n8201 , n4878 );
xor ( n8202 , n8200 , n8201 );
buf ( n8203 , n4879 );
xor ( n8204 , n8202 , n8203 );
xor ( n8205 , n8189 , n8204 );
not ( n8206 , n8205 );
not ( n8207 , n6474 );
buf ( n8208 , n4880 );
and ( n8209 , n8207 , n8208 );
buf ( n8210 , n4881 );
xor ( n8211 , n8210 , n8208 );
and ( n8212 , n8211 , n6474 );
or ( n8213 , n8209 , n8212 );
not ( n8214 , n6474 );
buf ( n8215 , n4882 );
and ( n8216 , n8214 , n8215 );
buf ( n8217 , n4883 );
xor ( n8218 , n8217 , n8215 );
and ( n8219 , n8218 , n6474 );
or ( n8220 , n8216 , n8219 );
xor ( n8221 , n8213 , n8220 );
buf ( n8222 , n4884 );
xor ( n8223 , n8221 , n8222 );
buf ( n8224 , n4885 );
xor ( n8225 , n8223 , n8224 );
buf ( n8226 , n4886 );
xor ( n8227 , n8225 , n8226 );
xor ( n8228 , n7433 , n8227 );
not ( n8229 , n6474 );
buf ( n8230 , n4887 );
and ( n8231 , n8229 , n8230 );
buf ( n8232 , n4888 );
xor ( n8233 , n8232 , n8230 );
and ( n8234 , n8233 , n6474 );
or ( n8235 , n8231 , n8234 );
not ( n8236 , n6474 );
buf ( n8237 , n4889 );
and ( n8238 , n8236 , n8237 );
buf ( n8239 , n4890 );
xor ( n8240 , n8239 , n8237 );
and ( n8241 , n8240 , n6474 );
or ( n8242 , n8238 , n8241 );
xor ( n8243 , n8235 , n8242 );
buf ( n8244 , n4891 );
xor ( n8245 , n8243 , n8244 );
buf ( n8246 , n4892 );
xor ( n8247 , n8245 , n8246 );
buf ( n8248 , n4893 );
xor ( n8249 , n8247 , n8248 );
xor ( n8250 , n8228 , n8249 );
and ( n8251 , n8206 , n8250 );
xor ( n8252 , n8166 , n8251 );
xor ( n8253 , n8163 , n8252 );
buf ( n8254 , n4894 );
not ( n8255 , n6474 );
buf ( n8256 , n4895 );
and ( n8257 , n8255 , n8256 );
buf ( n8258 , n4896 );
xor ( n8259 , n8258 , n8256 );
and ( n8260 , n8259 , n6474 );
or ( n8261 , n8257 , n8260 );
buf ( n8262 , n4897 );
xor ( n8263 , n8261 , n8262 );
buf ( n8264 , n4898 );
xor ( n8265 , n8263 , n8264 );
buf ( n8266 , n4899 );
xor ( n8267 , n8265 , n8266 );
buf ( n8268 , n4900 );
xor ( n8269 , n8267 , n8268 );
xor ( n8270 , n8254 , n8269 );
not ( n8271 , n6474 );
buf ( n8272 , n4901 );
and ( n8273 , n8271 , n8272 );
buf ( n8274 , n4902 );
xor ( n8275 , n8274 , n8272 );
and ( n8276 , n8275 , n6474 );
or ( n8277 , n8273 , n8276 );
not ( n8278 , n6474 );
buf ( n8279 , n4903 );
and ( n8280 , n8278 , n8279 );
buf ( n8281 , n4904 );
xor ( n8282 , n8281 , n8279 );
and ( n8283 , n8282 , n6474 );
or ( n8284 , n8280 , n8283 );
xor ( n8285 , n8277 , n8284 );
buf ( n8286 , n4905 );
xor ( n8287 , n8285 , n8286 );
buf ( n8288 , n4906 );
xor ( n8289 , n8287 , n8288 );
buf ( n8290 , n4907 );
xor ( n8291 , n8289 , n8290 );
xor ( n8292 , n8270 , n8291 );
buf ( n8293 , n4908 );
not ( n8294 , n6474 );
buf ( n8295 , n4909 );
and ( n8296 , n8294 , n8295 );
buf ( n8297 , n4910 );
xor ( n8298 , n8297 , n8295 );
and ( n8299 , n8298 , n6474 );
or ( n8300 , n8296 , n8299 );
not ( n8301 , n6474 );
buf ( n8302 , n4911 );
and ( n8303 , n8301 , n8302 );
buf ( n8304 , n4912 );
xor ( n8305 , n8304 , n8302 );
and ( n8306 , n8305 , n6474 );
or ( n8307 , n8303 , n8306 );
xor ( n8308 , n8300 , n8307 );
buf ( n8309 , n4913 );
xor ( n8310 , n8308 , n8309 );
buf ( n8311 , n4914 );
xor ( n8312 , n8310 , n8311 );
buf ( n8313 , n4915 );
xor ( n8314 , n8312 , n8313 );
xor ( n8315 , n8293 , n8314 );
not ( n8316 , n6474 );
buf ( n8317 , n4916 );
and ( n8318 , n8316 , n8317 );
buf ( n8319 , n4917 );
xor ( n8320 , n8319 , n8317 );
and ( n8321 , n8320 , n6474 );
or ( n8322 , n8318 , n8321 );
not ( n8323 , n6474 );
buf ( n8324 , n4918 );
and ( n8325 , n8323 , n8324 );
buf ( n8326 , n4919 );
xor ( n8327 , n8326 , n8324 );
and ( n8328 , n8327 , n6474 );
or ( n8329 , n8325 , n8328 );
xor ( n8330 , n8322 , n8329 );
buf ( n8331 , n4920 );
xor ( n8332 , n8330 , n8331 );
buf ( n8333 , n4921 );
xor ( n8334 , n8332 , n8333 );
buf ( n8335 , n4922 );
xor ( n8336 , n8334 , n8335 );
xor ( n8337 , n8315 , n8336 );
not ( n8338 , n8337 );
not ( n8339 , n6474 );
buf ( n8340 , n4923 );
and ( n8341 , n8339 , n8340 );
buf ( n8342 , n4924 );
xor ( n8343 , n8342 , n8340 );
and ( n8344 , n8343 , n6474 );
or ( n8345 , n8341 , n8344 );
not ( n8346 , n6474 );
buf ( n8347 , n4925 );
and ( n8348 , n8346 , n8347 );
buf ( n8349 , n4926 );
xor ( n8350 , n8349 , n8347 );
and ( n8351 , n8350 , n6474 );
or ( n8352 , n8348 , n8351 );
not ( n8353 , n6474 );
buf ( n8354 , n4927 );
and ( n8355 , n8353 , n8354 );
buf ( n8356 , n4928 );
xor ( n8357 , n8356 , n8354 );
and ( n8358 , n8357 , n6474 );
or ( n8359 , n8355 , n8358 );
xor ( n8360 , n8352 , n8359 );
buf ( n8361 , n4929 );
xor ( n8362 , n8360 , n8361 );
buf ( n8363 , n4930 );
xor ( n8364 , n8362 , n8363 );
buf ( n8365 , n4931 );
xor ( n8366 , n8364 , n8365 );
xor ( n8367 , n8345 , n8366 );
not ( n8368 , n6474 );
buf ( n8369 , n4932 );
and ( n8370 , n8368 , n8369 );
buf ( n8371 , n4933 );
xor ( n8372 , n8371 , n8369 );
and ( n8373 , n8372 , n6474 );
or ( n8374 , n8370 , n8373 );
not ( n8375 , n6474 );
buf ( n8376 , n4934 );
and ( n8377 , n8375 , n8376 );
buf ( n8378 , n4935 );
xor ( n8379 , n8378 , n8376 );
and ( n8380 , n8379 , n6474 );
or ( n8381 , n8377 , n8380 );
xor ( n8382 , n8374 , n8381 );
buf ( n8383 , n4936 );
xor ( n8384 , n8382 , n8383 );
buf ( n8385 , n4937 );
xor ( n8386 , n8384 , n8385 );
buf ( n8387 , n4938 );
xor ( n8388 , n8386 , n8387 );
xor ( n8389 , n8367 , n8388 );
and ( n8390 , n8338 , n8389 );
xor ( n8391 , n8292 , n8390 );
xor ( n8392 , n8253 , n8391 );
xor ( n8393 , n7886 , n8392 );
xor ( n8394 , n8123 , n7046 );
not ( n8395 , n6474 );
buf ( n8396 , n4939 );
and ( n8397 , n8395 , n8396 );
buf ( n8398 , n4940 );
xor ( n8399 , n8398 , n8396 );
and ( n8400 , n8399 , n6474 );
or ( n8401 , n8397 , n8400 );
not ( n8402 , n6474 );
buf ( n8403 , n4941 );
and ( n8404 , n8402 , n8403 );
buf ( n8405 , n4942 );
xor ( n8406 , n8405 , n8403 );
and ( n8407 , n8406 , n6474 );
or ( n8408 , n8404 , n8407 );
xor ( n8409 , n8401 , n8408 );
buf ( n8410 , n4943 );
xor ( n8411 , n8409 , n8410 );
buf ( n8412 , n4944 );
xor ( n8413 , n8411 , n8412 );
xor ( n8414 , n8413 , n8293 );
xor ( n8415 , n8394 , n8414 );
not ( n8416 , n6474 );
buf ( n8417 , n4945 );
and ( n8418 , n8416 , n8417 );
buf ( n8419 , n4946 );
xor ( n8420 , n8419 , n8417 );
and ( n8421 , n8420 , n6474 );
or ( n8422 , n8418 , n8421 );
xor ( n8423 , n8422 , n8034 );
xor ( n8424 , n8423 , n8056 );
not ( n8425 , n8424 );
buf ( n8426 , n4947 );
not ( n8427 , n6474 );
buf ( n8428 , n4948 );
and ( n8429 , n8427 , n8428 );
buf ( n8430 , n4949 );
xor ( n8431 , n8430 , n8428 );
and ( n8432 , n8431 , n6474 );
or ( n8433 , n8429 , n8432 );
not ( n8434 , n6474 );
buf ( n8435 , n4950 );
and ( n8436 , n8434 , n8435 );
buf ( n8437 , n4951 );
xor ( n8438 , n8437 , n8435 );
and ( n8439 , n8438 , n6474 );
or ( n8440 , n8436 , n8439 );
xor ( n8441 , n8433 , n8440 );
buf ( n8442 , n4952 );
xor ( n8443 , n8441 , n8442 );
buf ( n8444 , n4953 );
xor ( n8445 , n8443 , n8444 );
buf ( n8446 , n4954 );
xor ( n8447 , n8445 , n8446 );
xor ( n8448 , n8426 , n8447 );
not ( n8449 , n6474 );
buf ( n8450 , n4955 );
and ( n8451 , n8449 , n8450 );
buf ( n8452 , n4956 );
xor ( n8453 , n8452 , n8450 );
and ( n8454 , n8453 , n6474 );
or ( n8455 , n8451 , n8454 );
not ( n8456 , n6474 );
buf ( n8457 , n4957 );
and ( n8458 , n8456 , n8457 );
buf ( n8459 , n4958 );
xor ( n8460 , n8459 , n8457 );
and ( n8461 , n8460 , n6474 );
or ( n8462 , n8458 , n8461 );
xor ( n8463 , n8455 , n8462 );
buf ( n8464 , n4959 );
xor ( n8465 , n8463 , n8464 );
buf ( n8466 , n4960 );
xor ( n8467 , n8465 , n8466 );
buf ( n8468 , n4961 );
xor ( n8469 , n8467 , n8468 );
xor ( n8470 , n8448 , n8469 );
and ( n8471 , n8425 , n8470 );
xor ( n8472 , n8415 , n8471 );
xor ( n8473 , n7386 , n6500 );
xor ( n8474 , n8473 , n6516 );
buf ( n8475 , n4962 );
not ( n8476 , n6474 );
buf ( n8477 , n4963 );
and ( n8478 , n8476 , n8477 );
buf ( n8479 , n4964 );
xor ( n8480 , n8479 , n8477 );
and ( n8481 , n8480 , n6474 );
or ( n8482 , n8478 , n8481 );
not ( n8483 , n6474 );
buf ( n8484 , n4965 );
and ( n8485 , n8483 , n8484 );
buf ( n8486 , n4966 );
xor ( n8487 , n8486 , n8484 );
and ( n8488 , n8487 , n6474 );
or ( n8489 , n8485 , n8488 );
xor ( n8490 , n8482 , n8489 );
buf ( n8491 , n4967 );
xor ( n8492 , n8490 , n8491 );
xor ( n8493 , n8492 , n7889 );
buf ( n8494 , n4968 );
xor ( n8495 , n8493 , n8494 );
xor ( n8496 , n8475 , n8495 );
not ( n8497 , n6474 );
buf ( n8498 , n4969 );
and ( n8499 , n8497 , n8498 );
buf ( n8500 , n4970 );
xor ( n8501 , n8500 , n8498 );
and ( n8502 , n8501 , n6474 );
or ( n8503 , n8499 , n8502 );
not ( n8504 , n6474 );
buf ( n8505 , n4971 );
and ( n8506 , n8504 , n8505 );
buf ( n8507 , n4972 );
xor ( n8508 , n8507 , n8505 );
and ( n8509 , n8508 , n6474 );
or ( n8510 , n8506 , n8509 );
xor ( n8511 , n8503 , n8510 );
buf ( n8512 , n4973 );
xor ( n8513 , n8511 , n8512 );
buf ( n8514 , n4974 );
xor ( n8515 , n8513 , n8514 );
buf ( n8516 , n4975 );
xor ( n8517 , n8515 , n8516 );
xor ( n8518 , n8496 , n8517 );
not ( n8519 , n8518 );
buf ( n8520 , n4976 );
not ( n8521 , n6474 );
buf ( n8522 , n4977 );
and ( n8523 , n8521 , n8522 );
buf ( n8524 , n4978 );
xor ( n8525 , n8524 , n8522 );
and ( n8526 , n8525 , n6474 );
or ( n8527 , n8523 , n8526 );
buf ( n8528 , n4979 );
xor ( n8529 , n8527 , n8528 );
buf ( n8530 , n4980 );
xor ( n8531 , n8529 , n8530 );
buf ( n8532 , n4981 );
xor ( n8533 , n8531 , n8532 );
buf ( n8534 , n4982 );
xor ( n8535 , n8533 , n8534 );
xor ( n8536 , n8520 , n8535 );
xor ( n8537 , n8536 , n6763 );
and ( n8538 , n8519 , n8537 );
xor ( n8539 , n8474 , n8538 );
xor ( n8540 , n8472 , n8539 );
xor ( n8541 , n8401 , n8314 );
xor ( n8542 , n8541 , n8336 );
not ( n8543 , n6474 );
buf ( n8544 , n4983 );
and ( n8545 , n8543 , n8544 );
buf ( n8546 , n4984 );
xor ( n8547 , n8546 , n8544 );
and ( n8548 , n8547 , n6474 );
or ( n8549 , n8545 , n8548 );
xor ( n8550 , n8549 , n7710 );
xor ( n8551 , n8550 , n7732 );
not ( n8552 , n8551 );
buf ( n8553 , n4985 );
not ( n8554 , n6474 );
buf ( n8555 , n4986 );
and ( n8556 , n8554 , n8555 );
buf ( n8557 , n4987 );
xor ( n8558 , n8557 , n8555 );
and ( n8559 , n8558 , n6474 );
or ( n8560 , n8556 , n8559 );
not ( n8561 , n6474 );
buf ( n8562 , n4988 );
and ( n8563 , n8561 , n8562 );
buf ( n8564 , n4989 );
xor ( n8565 , n8564 , n8562 );
and ( n8566 , n8565 , n6474 );
or ( n8567 , n8563 , n8566 );
xor ( n8568 , n8560 , n8567 );
buf ( n8569 , n4990 );
xor ( n8570 , n8568 , n8569 );
buf ( n8571 , n4991 );
xor ( n8572 , n8570 , n8571 );
buf ( n8573 , n4992 );
xor ( n8574 , n8572 , n8573 );
xor ( n8575 , n8553 , n8574 );
xor ( n8576 , n8575 , n7441 );
and ( n8577 , n8552 , n8576 );
xor ( n8578 , n8542 , n8577 );
xor ( n8579 , n8540 , n8578 );
not ( n8580 , n6474 );
buf ( n8581 , n4993 );
and ( n8582 , n8580 , n8581 );
buf ( n8583 , n4994 );
xor ( n8584 , n8583 , n8581 );
and ( n8585 , n8584 , n6474 );
or ( n8586 , n8582 , n8585 );
not ( n8587 , n6474 );
buf ( n8588 , n4995 );
and ( n8589 , n8587 , n8588 );
buf ( n8590 , n4996 );
xor ( n8591 , n8590 , n8588 );
and ( n8592 , n8591 , n6474 );
or ( n8593 , n8589 , n8592 );
xor ( n8594 , n7801 , n8593 );
buf ( n8595 , n4997 );
xor ( n8596 , n8594 , n8595 );
buf ( n8597 , n4998 );
xor ( n8598 , n8596 , n8597 );
buf ( n8599 , n4999 );
xor ( n8600 , n8598 , n8599 );
xor ( n8601 , n8586 , n8600 );
not ( n8602 , n6474 );
buf ( n8603 , n5000 );
and ( n8604 , n8602 , n8603 );
buf ( n8605 , n5001 );
xor ( n8606 , n8605 , n8603 );
and ( n8607 , n8606 , n6474 );
or ( n8608 , n8604 , n8607 );
not ( n8609 , n6474 );
buf ( n8610 , n5002 );
and ( n8611 , n8609 , n8610 );
buf ( n8612 , n5003 );
xor ( n8613 , n8612 , n8610 );
and ( n8614 , n8613 , n6474 );
or ( n8615 , n8611 , n8614 );
xor ( n8616 , n8608 , n8615 );
buf ( n8617 , n5004 );
xor ( n8618 , n8616 , n8617 );
buf ( n8619 , n5005 );
xor ( n8620 , n8618 , n8619 );
buf ( n8621 , n5006 );
xor ( n8622 , n8620 , n8621 );
xor ( n8623 , n8601 , n8622 );
not ( n8624 , n6474 );
buf ( n8625 , n5007 );
and ( n8626 , n8624 , n8625 );
buf ( n8627 , n5008 );
xor ( n8628 , n8627 , n8625 );
and ( n8629 , n8628 , n6474 );
or ( n8630 , n8626 , n8629 );
buf ( n8631 , n5009 );
xor ( n8632 , n8630 , n8631 );
buf ( n8633 , n5010 );
xor ( n8634 , n8632 , n8633 );
buf ( n8635 , n5011 );
xor ( n8636 , n8634 , n8635 );
buf ( n8637 , n5012 );
xor ( n8638 , n8636 , n8637 );
xor ( n8639 , n7581 , n8638 );
not ( n8640 , n6474 );
buf ( n8641 , n5013 );
and ( n8642 , n8640 , n8641 );
buf ( n8643 , n5014 );
xor ( n8644 , n8643 , n8641 );
and ( n8645 , n8644 , n6474 );
or ( n8646 , n8642 , n8645 );
not ( n8647 , n6474 );
buf ( n8648 , n5015 );
and ( n8649 , n8647 , n8648 );
buf ( n8650 , n5016 );
xor ( n8651 , n8650 , n8648 );
and ( n8652 , n8651 , n6474 );
or ( n8653 , n8649 , n8652 );
xor ( n8654 , n8646 , n8653 );
buf ( n8655 , n5017 );
xor ( n8656 , n8654 , n8655 );
buf ( n8657 , n5018 );
xor ( n8658 , n8656 , n8657 );
buf ( n8659 , n5019 );
xor ( n8660 , n8658 , n8659 );
xor ( n8661 , n8639 , n8660 );
not ( n8662 , n8661 );
buf ( n8663 , n5020 );
xor ( n8664 , n8663 , n7659 );
xor ( n8665 , n8664 , n7681 );
and ( n8666 , n8662 , n8665 );
xor ( n8667 , n8623 , n8666 );
xor ( n8668 , n8579 , n8667 );
not ( n8669 , n6474 );
buf ( n8670 , n5021 );
and ( n8671 , n8669 , n8670 );
buf ( n8672 , n5022 );
xor ( n8673 , n8672 , n8670 );
and ( n8674 , n8673 , n6474 );
or ( n8675 , n8671 , n8674 );
not ( n8676 , n6474 );
buf ( n8677 , n5023 );
and ( n8678 , n8676 , n8677 );
buf ( n8679 , n5024 );
xor ( n8680 , n8679 , n8677 );
and ( n8681 , n8680 , n6474 );
or ( n8682 , n8678 , n8681 );
not ( n8683 , n6474 );
buf ( n8684 , n5025 );
and ( n8685 , n8683 , n8684 );
buf ( n8686 , n5026 );
xor ( n8687 , n8686 , n8684 );
and ( n8688 , n8687 , n6474 );
or ( n8689 , n8685 , n8688 );
xor ( n8690 , n8682 , n8689 );
buf ( n8691 , n5027 );
xor ( n8692 , n8690 , n8691 );
buf ( n8693 , n5028 );
xor ( n8694 , n8692 , n8693 );
buf ( n8695 , n5029 );
xor ( n8696 , n8694 , n8695 );
xor ( n8697 , n8675 , n8696 );
not ( n8698 , n6474 );
buf ( n8699 , n5030 );
and ( n8700 , n8698 , n8699 );
buf ( n8701 , n5031 );
xor ( n8702 , n8701 , n8699 );
and ( n8703 , n8702 , n6474 );
or ( n8704 , n8700 , n8703 );
xor ( n8705 , n8704 , n7741 );
buf ( n8706 , n5032 );
xor ( n8707 , n8705 , n8706 );
buf ( n8708 , n5033 );
xor ( n8709 , n8707 , n8708 );
xor ( n8710 , n8709 , n7009 );
xor ( n8711 , n8697 , n8710 );
not ( n8712 , n6474 );
buf ( n8713 , n5034 );
and ( n8714 , n8712 , n8713 );
buf ( n8715 , n5035 );
xor ( n8716 , n8715 , n8713 );
and ( n8717 , n8716 , n6474 );
or ( n8718 , n8714 , n8717 );
xor ( n8719 , n8718 , n8188 );
xor ( n8720 , n8719 , n8204 );
not ( n8721 , n8720 );
buf ( n8722 , n5036 );
not ( n8723 , n6474 );
buf ( n8724 , n5037 );
and ( n8725 , n8723 , n8724 );
buf ( n8726 , n5038 );
xor ( n8727 , n8726 , n8724 );
and ( n8728 , n8727 , n6474 );
or ( n8729 , n8725 , n8728 );
not ( n8730 , n6474 );
buf ( n8731 , n5039 );
and ( n8732 , n8730 , n8731 );
buf ( n8733 , n5040 );
xor ( n8734 , n8733 , n8731 );
and ( n8735 , n8734 , n6474 );
or ( n8736 , n8732 , n8735 );
xor ( n8737 , n8729 , n8736 );
buf ( n8738 , n5041 );
xor ( n8739 , n8737 , n8738 );
buf ( n8740 , n5042 );
xor ( n8741 , n8739 , n8740 );
buf ( n8742 , n5043 );
xor ( n8743 , n8741 , n8742 );
xor ( n8744 , n8722 , n8743 );
not ( n8745 , n6474 );
buf ( n8746 , n5044 );
and ( n8747 , n8745 , n8746 );
buf ( n8748 , n5045 );
xor ( n8749 , n8748 , n8746 );
and ( n8750 , n8749 , n6474 );
or ( n8751 , n8747 , n8750 );
not ( n8752 , n6474 );
buf ( n8753 , n5046 );
and ( n8754 , n8752 , n8753 );
buf ( n8755 , n5047 );
xor ( n8756 , n8755 , n8753 );
and ( n8757 , n8756 , n6474 );
or ( n8758 , n8754 , n8757 );
xor ( n8759 , n8751 , n8758 );
buf ( n8760 , n5048 );
xor ( n8761 , n8759 , n8760 );
xor ( n8762 , n8761 , n8254 );
buf ( n8763 , n5049 );
xor ( n8764 , n8762 , n8763 );
xor ( n8765 , n8744 , n8764 );
and ( n8766 , n8721 , n8765 );
xor ( n8767 , n8711 , n8766 );
xor ( n8768 , n8668 , n8767 );
xor ( n8769 , n8393 , n8768 );
not ( n8770 , n8769 );
not ( n8771 , n6474 );
buf ( n8772 , n5050 );
and ( n8773 , n8771 , n8772 );
buf ( n8774 , n5051 );
xor ( n8775 , n8774 , n8772 );
and ( n8776 , n8775 , n6474 );
or ( n8777 , n8773 , n8776 );
xor ( n8778 , n8777 , n7095 );
not ( n8779 , n6474 );
buf ( n8780 , n5052 );
and ( n8781 , n8779 , n8780 );
buf ( n8782 , n5053 );
xor ( n8783 , n8782 , n8780 );
and ( n8784 , n8783 , n6474 );
or ( n8785 , n8781 , n8784 );
not ( n8786 , n6474 );
buf ( n8787 , n5054 );
and ( n8788 , n8786 , n8787 );
buf ( n8789 , n5055 );
xor ( n8790 , n8789 , n8787 );
and ( n8791 , n8790 , n6474 );
or ( n8792 , n8788 , n8791 );
xor ( n8793 , n8785 , n8792 );
buf ( n8794 , n5056 );
xor ( n8795 , n8793 , n8794 );
buf ( n8796 , n5057 );
xor ( n8797 , n8795 , n8796 );
buf ( n8798 , n5058 );
xor ( n8799 , n8797 , n8798 );
xor ( n8800 , n8778 , n8799 );
not ( n8801 , n6474 );
buf ( n8802 , n5059 );
and ( n8803 , n8801 , n8802 );
buf ( n8804 , n5060 );
xor ( n8805 , n8804 , n8802 );
and ( n8806 , n8805 , n6474 );
or ( n8807 , n8803 , n8806 );
not ( n8808 , n6474 );
buf ( n8809 , n5061 );
and ( n8810 , n8808 , n8809 );
buf ( n8811 , n5062 );
xor ( n8812 , n8811 , n8809 );
and ( n8813 , n8812 , n6474 );
or ( n8814 , n8810 , n8813 );
xor ( n8815 , n8814 , n7283 );
buf ( n8816 , n5063 );
xor ( n8817 , n8815 , n8816 );
xor ( n8818 , n8817 , n6697 );
buf ( n8819 , n5064 );
xor ( n8820 , n8818 , n8819 );
xor ( n8821 , n8807 , n8820 );
not ( n8822 , n6474 );
buf ( n8823 , n5065 );
and ( n8824 , n8822 , n8823 );
buf ( n8825 , n5066 );
xor ( n8826 , n8825 , n8823 );
and ( n8827 , n8826 , n6474 );
or ( n8828 , n8824 , n8827 );
not ( n8829 , n6474 );
buf ( n8830 , n5067 );
and ( n8831 , n8829 , n8830 );
buf ( n8832 , n5068 );
xor ( n8833 , n8832 , n8830 );
and ( n8834 , n8833 , n6474 );
or ( n8835 , n8831 , n8834 );
xor ( n8836 , n8828 , n8835 );
buf ( n8837 , n5069 );
xor ( n8838 , n8836 , n8837 );
buf ( n8839 , n5070 );
xor ( n8840 , n8838 , n8839 );
buf ( n8841 , n5071 );
xor ( n8842 , n8840 , n8841 );
xor ( n8843 , n8821 , n8842 );
not ( n8844 , n8843 );
not ( n8845 , n6474 );
buf ( n8846 , n5072 );
and ( n8847 , n8845 , n8846 );
buf ( n8848 , n5073 );
xor ( n8849 , n8848 , n8846 );
and ( n8850 , n8849 , n6474 );
or ( n8851 , n8847 , n8850 );
not ( n8852 , n6474 );
buf ( n8853 , n5074 );
and ( n8854 , n8852 , n8853 );
buf ( n8855 , n5075 );
xor ( n8856 , n8855 , n8853 );
and ( n8857 , n8856 , n6474 );
or ( n8858 , n8854 , n8857 );
xor ( n8859 , n8851 , n8858 );
buf ( n8860 , n5076 );
xor ( n8861 , n8859 , n8860 );
buf ( n8862 , n5077 );
xor ( n8863 , n8861 , n8862 );
buf ( n8864 , n5078 );
xor ( n8865 , n8863 , n8864 );
xor ( n8866 , n7727 , n8865 );
xor ( n8867 , n8866 , n7253 );
and ( n8868 , n8844 , n8867 );
xor ( n8869 , n8800 , n8868 );
buf ( n8870 , n5079 );
not ( n8871 , n6474 );
buf ( n8872 , n5080 );
and ( n8873 , n8871 , n8872 );
buf ( n8874 , n5081 );
xor ( n8875 , n8874 , n8872 );
and ( n8876 , n8875 , n6474 );
or ( n8877 , n8873 , n8876 );
not ( n8878 , n6474 );
buf ( n8879 , n5082 );
and ( n8880 , n8878 , n8879 );
buf ( n8881 , n5083 );
xor ( n8882 , n8881 , n8879 );
and ( n8883 , n8882 , n6474 );
or ( n8884 , n8880 , n8883 );
xor ( n8885 , n8877 , n8884 );
buf ( n8886 , n5084 );
xor ( n8887 , n8885 , n8886 );
buf ( n8888 , n5085 );
xor ( n8889 , n8887 , n8888 );
buf ( n8890 , n5086 );
xor ( n8891 , n8889 , n8890 );
xor ( n8892 , n8870 , n8891 );
not ( n8893 , n6474 );
buf ( n8894 , n5087 );
and ( n8895 , n8893 , n8894 );
buf ( n8896 , n5088 );
xor ( n8897 , n8896 , n8894 );
and ( n8898 , n8897 , n6474 );
or ( n8899 , n8895 , n8898 );
not ( n8900 , n6474 );
buf ( n8901 , n5089 );
and ( n8902 , n8900 , n8901 );
buf ( n8903 , n5090 );
xor ( n8904 , n8903 , n8901 );
and ( n8905 , n8904 , n6474 );
or ( n8906 , n8902 , n8905 );
xor ( n8907 , n8899 , n8906 );
buf ( n8908 , n5091 );
xor ( n8909 , n8907 , n8908 );
buf ( n8910 , n5092 );
xor ( n8911 , n8909 , n8910 );
buf ( n8912 , n5093 );
xor ( n8913 , n8911 , n8912 );
xor ( n8914 , n8892 , n8913 );
not ( n8915 , n6474 );
buf ( n8916 , n5094 );
and ( n8917 , n8915 , n8916 );
buf ( n8918 , n5095 );
xor ( n8919 , n8918 , n8916 );
and ( n8920 , n8919 , n6474 );
or ( n8921 , n8917 , n8920 );
not ( n8922 , n6474 );
buf ( n8923 , n5096 );
and ( n8924 , n8922 , n8923 );
buf ( n8925 , n5097 );
xor ( n8926 , n8925 , n8923 );
and ( n8927 , n8926 , n6474 );
or ( n8928 , n8924 , n8927 );
buf ( n8929 , n5098 );
xor ( n8930 , n8928 , n8929 );
xor ( n8931 , n8930 , n7051 );
buf ( n8932 , n5099 );
xor ( n8933 , n8931 , n8932 );
buf ( n8934 , n5100 );
xor ( n8935 , n8933 , n8934 );
xor ( n8936 , n8921 , n8935 );
not ( n8937 , n6474 );
buf ( n8938 , n5101 );
and ( n8939 , n8937 , n8938 );
buf ( n8940 , n5102 );
xor ( n8941 , n8940 , n8938 );
and ( n8942 , n8941 , n6474 );
or ( n8943 , n8939 , n8942 );
xor ( n8944 , n8777 , n8943 );
buf ( n8945 , n5103 );
xor ( n8946 , n8944 , n8945 );
buf ( n8947 , n5104 );
xor ( n8948 , n8946 , n8947 );
buf ( n8949 , n5105 );
xor ( n8950 , n8948 , n8949 );
xor ( n8951 , n8936 , n8950 );
not ( n8952 , n8951 );
not ( n8953 , n6474 );
buf ( n8954 , n5106 );
and ( n8955 , n8953 , n8954 );
buf ( n8956 , n5107 );
xor ( n8957 , n8956 , n8954 );
and ( n8958 , n8957 , n6474 );
or ( n8959 , n8955 , n8958 );
not ( n8960 , n6474 );
buf ( n8961 , n5108 );
and ( n8962 , n8960 , n8961 );
buf ( n8963 , n5109 );
xor ( n8964 , n8963 , n8961 );
and ( n8965 , n8964 , n6474 );
or ( n8966 , n8962 , n8965 );
xor ( n8967 , n8959 , n8966 );
buf ( n8968 , n5110 );
xor ( n8969 , n8967 , n8968 );
buf ( n8970 , n5111 );
xor ( n8971 , n8969 , n8970 );
xor ( n8972 , n8971 , n7426 );
xor ( n8973 , n6906 , n8972 );
xor ( n8974 , n8973 , n7822 );
and ( n8975 , n8952 , n8974 );
xor ( n8976 , n8914 , n8975 );
buf ( n8977 , n5112 );
xor ( n8978 , n8977 , n8447 );
xor ( n8979 , n8978 , n8469 );
not ( n8980 , n6474 );
buf ( n8981 , n5113 );
and ( n8982 , n8980 , n8981 );
buf ( n8983 , n5114 );
xor ( n8984 , n8983 , n8981 );
and ( n8985 , n8984 , n6474 );
or ( n8986 , n8982 , n8985 );
xor ( n8987 , n8986 , n7181 );
not ( n8988 , n6474 );
buf ( n8989 , n5115 );
and ( n8990 , n8988 , n8989 );
buf ( n8991 , n5116 );
xor ( n8992 , n8991 , n8989 );
and ( n8993 , n8992 , n6474 );
or ( n8994 , n8990 , n8993 );
buf ( n8995 , n5117 );
xor ( n8996 , n8994 , n8995 );
buf ( n8997 , n5118 );
xor ( n8998 , n8996 , n8997 );
buf ( n8999 , n5119 );
xor ( n9000 , n8998 , n8999 );
buf ( n9001 , n5120 );
xor ( n9002 , n9000 , n9001 );
xor ( n9003 , n8987 , n9002 );
not ( n9004 , n9003 );
buf ( n9005 , n5121 );
not ( n9006 , n6474 );
buf ( n9007 , n5122 );
and ( n9008 , n9006 , n9007 );
buf ( n9009 , n5123 );
xor ( n9010 , n9009 , n9007 );
and ( n9011 , n9010 , n6474 );
or ( n9012 , n9008 , n9011 );
not ( n9013 , n6474 );
buf ( n9014 , n5124 );
and ( n9015 , n9013 , n9014 );
buf ( n9016 , n5125 );
xor ( n9017 , n9016 , n9014 );
and ( n9018 , n9017 , n6474 );
or ( n9019 , n9015 , n9018 );
xor ( n9020 , n9012 , n9019 );
buf ( n9021 , n5126 );
xor ( n9022 , n9020 , n9021 );
buf ( n9023 , n5127 );
xor ( n9024 , n9022 , n9023 );
buf ( n9025 , n5128 );
xor ( n9026 , n9024 , n9025 );
xor ( n9027 , n9005 , n9026 );
not ( n9028 , n6474 );
buf ( n9029 , n5129 );
and ( n9030 , n9028 , n9029 );
buf ( n9031 , n5130 );
xor ( n9032 , n9031 , n9029 );
and ( n9033 , n9032 , n6474 );
or ( n9034 , n9030 , n9033 );
not ( n9035 , n6474 );
buf ( n9036 , n5131 );
and ( n9037 , n9035 , n9036 );
buf ( n9038 , n5132 );
xor ( n9039 , n9038 , n9036 );
and ( n9040 , n9039 , n6474 );
or ( n9041 , n9037 , n9040 );
xor ( n9042 , n9034 , n9041 );
xor ( n9043 , n9042 , n8520 );
buf ( n9044 , n5133 );
xor ( n9045 , n9043 , n9044 );
buf ( n9046 , n5134 );
xor ( n9047 , n9045 , n9046 );
xor ( n9048 , n9027 , n9047 );
and ( n9049 , n9004 , n9048 );
xor ( n9050 , n8979 , n9049 );
xor ( n9051 , n8976 , n9050 );
xor ( n9052 , n8136 , n7046 );
xor ( n9053 , n9052 , n8414 );
not ( n9054 , n8800 );
and ( n9055 , n9054 , n8843 );
xor ( n9056 , n9053 , n9055 );
xor ( n9057 , n9051 , n9056 );
buf ( n9058 , n5135 );
not ( n9059 , n6474 );
buf ( n9060 , n5136 );
and ( n9061 , n9059 , n9060 );
buf ( n9062 , n5137 );
xor ( n9063 , n9062 , n9060 );
and ( n9064 , n9063 , n6474 );
or ( n9065 , n9061 , n9064 );
not ( n9066 , n6474 );
buf ( n9067 , n5138 );
and ( n9068 , n9066 , n9067 );
buf ( n9069 , n5139 );
xor ( n9070 , n9069 , n9067 );
and ( n9071 , n9070 , n6474 );
or ( n9072 , n9068 , n9071 );
xor ( n9073 , n9065 , n9072 );
buf ( n9074 , n5140 );
xor ( n9075 , n9073 , n9074 );
buf ( n9076 , n5141 );
xor ( n9077 , n9075 , n9076 );
buf ( n9078 , n5142 );
xor ( n9079 , n9077 , n9078 );
xor ( n9080 , n9058 , n9079 );
not ( n9081 , n6474 );
buf ( n9082 , n5143 );
and ( n9083 , n9081 , n9082 );
buf ( n9084 , n5144 );
xor ( n9085 , n9084 , n9082 );
and ( n9086 , n9085 , n6474 );
or ( n9087 , n9083 , n9086 );
buf ( n9088 , n5145 );
xor ( n9089 , n9087 , n9088 );
xor ( n9090 , n9089 , n8722 );
buf ( n9091 , n5146 );
xor ( n9092 , n9090 , n9091 );
buf ( n9093 , n5147 );
xor ( n9094 , n9092 , n9093 );
xor ( n9095 , n9080 , n9094 );
not ( n9096 , n6474 );
buf ( n9097 , n5148 );
and ( n9098 , n9096 , n9097 );
buf ( n9099 , n5149 );
xor ( n9100 , n9099 , n9097 );
and ( n9101 , n9100 , n6474 );
or ( n9102 , n9098 , n9101 );
not ( n9103 , n6474 );
buf ( n9104 , n5150 );
and ( n9105 , n9103 , n9104 );
buf ( n9106 , n5151 );
xor ( n9107 , n9106 , n9104 );
and ( n9108 , n9107 , n6474 );
or ( n9109 , n9105 , n9108 );
not ( n9110 , n6474 );
buf ( n9111 , n5152 );
and ( n9112 , n9110 , n9111 );
buf ( n9113 , n5153 );
xor ( n9114 , n9113 , n9111 );
and ( n9115 , n9114 , n6474 );
or ( n9116 , n9112 , n9115 );
xor ( n9117 , n9109 , n9116 );
buf ( n9118 , n5154 );
xor ( n9119 , n9117 , n9118 );
buf ( n9120 , n5155 );
xor ( n9121 , n9119 , n9120 );
buf ( n9122 , n5156 );
xor ( n9123 , n9121 , n9122 );
xor ( n9124 , n9102 , n9123 );
xor ( n9125 , n9124 , n7659 );
not ( n9126 , n9125 );
not ( n9127 , n6474 );
buf ( n9128 , n5157 );
and ( n9129 , n9127 , n9128 );
buf ( n9130 , n5158 );
xor ( n9131 , n9130 , n9128 );
and ( n9132 , n9131 , n6474 );
or ( n9133 , n9129 , n9132 );
not ( n9134 , n6474 );
buf ( n9135 , n5159 );
and ( n9136 , n9134 , n9135 );
buf ( n9137 , n5160 );
xor ( n9138 , n9137 , n9135 );
and ( n9139 , n9138 , n6474 );
or ( n9140 , n9136 , n9139 );
buf ( n9141 , n5161 );
xor ( n9142 , n9140 , n9141 );
buf ( n9143 , n5162 );
xor ( n9144 , n9142 , n9143 );
buf ( n9145 , n5163 );
xor ( n9146 , n9144 , n9145 );
buf ( n9147 , n5164 );
xor ( n9148 , n9146 , n9147 );
xor ( n9149 , n9133 , n9148 );
not ( n9150 , n6474 );
buf ( n9151 , n5165 );
and ( n9152 , n9150 , n9151 );
buf ( n9153 , n5166 );
xor ( n9154 , n9153 , n9151 );
and ( n9155 , n9154 , n6474 );
or ( n9156 , n9152 , n9155 );
not ( n9157 , n6474 );
buf ( n9158 , n5167 );
and ( n9159 , n9157 , n9158 );
buf ( n9160 , n5168 );
xor ( n9161 , n9160 , n9158 );
and ( n9162 , n9161 , n6474 );
or ( n9163 , n9159 , n9162 );
xor ( n9164 , n9156 , n9163 );
buf ( n9165 , n5169 );
xor ( n9166 , n9164 , n9165 );
buf ( n9167 , n5170 );
xor ( n9168 , n9166 , n9167 );
buf ( n9169 , n5171 );
xor ( n9170 , n9168 , n9169 );
xor ( n9171 , n9149 , n9170 );
and ( n9172 , n9126 , n9171 );
xor ( n9173 , n9095 , n9172 );
xor ( n9174 , n9057 , n9173 );
buf ( n9175 , n5172 );
not ( n9176 , n6474 );
buf ( n9177 , n5173 );
and ( n9178 , n9176 , n9177 );
buf ( n9179 , n5174 );
xor ( n9180 , n9179 , n9177 );
and ( n9181 , n9180 , n6474 );
or ( n9182 , n9178 , n9181 );
not ( n9183 , n6474 );
buf ( n9184 , n5175 );
and ( n9185 , n9183 , n9184 );
buf ( n9186 , n5176 );
xor ( n9187 , n9186 , n9184 );
and ( n9188 , n9187 , n6474 );
or ( n9189 , n9185 , n9188 );
xor ( n9190 , n9182 , n9189 );
buf ( n9191 , n5177 );
xor ( n9192 , n9190 , n9191 );
xor ( n9193 , n9192 , n7097 );
buf ( n9194 , n5178 );
xor ( n9195 , n9193 , n9194 );
xor ( n9196 , n9175 , n9195 );
not ( n9197 , n6474 );
buf ( n9198 , n5179 );
and ( n9199 , n9197 , n9198 );
buf ( n9200 , n5180 );
xor ( n9201 , n9200 , n9198 );
and ( n9202 , n9201 , n6474 );
or ( n9203 , n9199 , n9202 );
not ( n9204 , n6474 );
buf ( n9205 , n5181 );
and ( n9206 , n9204 , n9205 );
buf ( n9207 , n5182 );
xor ( n9208 , n9207 , n9205 );
and ( n9209 , n9208 , n6474 );
or ( n9210 , n9206 , n9209 );
xor ( n9211 , n9203 , n9210 );
buf ( n9212 , n5183 );
xor ( n9213 , n9211 , n9212 );
buf ( n9214 , n5184 );
xor ( n9215 , n9213 , n9214 );
buf ( n9216 , n5185 );
xor ( n9217 , n9215 , n9216 );
xor ( n9218 , n9196 , n9217 );
not ( n9219 , n6474 );
buf ( n9220 , n5186 );
and ( n9221 , n9219 , n9220 );
buf ( n9222 , n5187 );
xor ( n9223 , n9222 , n9220 );
and ( n9224 , n9223 , n6474 );
or ( n9225 , n9221 , n9224 );
not ( n9226 , n6474 );
buf ( n9227 , n5188 );
and ( n9228 , n9226 , n9227 );
buf ( n9229 , n5189 );
xor ( n9230 , n9229 , n9227 );
and ( n9231 , n9230 , n6474 );
or ( n9232 , n9228 , n9231 );
xor ( n9233 , n9232 , n8422 );
buf ( n9234 , n5190 );
xor ( n9235 , n9233 , n9234 );
xor ( n9236 , n9235 , n8020 );
buf ( n9237 , n5191 );
xor ( n9238 , n9236 , n9237 );
xor ( n9239 , n9225 , n9238 );
not ( n9240 , n6474 );
buf ( n9241 , n5192 );
and ( n9242 , n9240 , n9241 );
buf ( n9243 , n5193 );
xor ( n9244 , n9243 , n9241 );
and ( n9245 , n9244 , n6474 );
or ( n9246 , n9242 , n9245 );
not ( n9247 , n6474 );
buf ( n9248 , n5194 );
and ( n9249 , n9247 , n9248 );
buf ( n9250 , n5195 );
xor ( n9251 , n9250 , n9248 );
and ( n9252 , n9251 , n6474 );
or ( n9253 , n9249 , n9252 );
xor ( n9254 , n9246 , n9253 );
buf ( n9255 , n5196 );
xor ( n9256 , n9254 , n9255 );
buf ( n9257 , n5197 );
xor ( n9258 , n9256 , n9257 );
buf ( n9259 , n5198 );
xor ( n9260 , n9258 , n9259 );
xor ( n9261 , n9239 , n9260 );
not ( n9262 , n9261 );
not ( n9263 , n6474 );
buf ( n9264 , n5199 );
and ( n9265 , n9263 , n9264 );
buf ( n9266 , n5200 );
xor ( n9267 , n9266 , n9264 );
and ( n9268 , n9267 , n6474 );
or ( n9269 , n9265 , n9268 );
not ( n9270 , n6474 );
buf ( n9271 , n5201 );
and ( n9272 , n9270 , n9271 );
buf ( n9273 , n5202 );
xor ( n9274 , n9273 , n9271 );
and ( n9275 , n9274 , n6474 );
or ( n9276 , n9272 , n9275 );
not ( n9277 , n6474 );
buf ( n9278 , n5203 );
and ( n9279 , n9277 , n9278 );
buf ( n9280 , n5204 );
xor ( n9281 , n9280 , n9278 );
and ( n9282 , n9281 , n6474 );
or ( n9283 , n9279 , n9282 );
xor ( n9284 , n9276 , n9283 );
buf ( n9285 , n5205 );
xor ( n9286 , n9284 , n9285 );
buf ( n9287 , n5206 );
xor ( n9288 , n9286 , n9287 );
buf ( n9289 , n5207 );
xor ( n9290 , n9288 , n9289 );
xor ( n9291 , n9269 , n9290 );
not ( n9292 , n6474 );
buf ( n9293 , n5208 );
and ( n9294 , n9292 , n9293 );
buf ( n9295 , n5209 );
xor ( n9296 , n9295 , n9293 );
and ( n9297 , n9296 , n6474 );
or ( n9298 , n9294 , n9297 );
buf ( n9299 , n5210 );
xor ( n9300 , n9298 , n9299 );
buf ( n9301 , n5211 );
xor ( n9302 , n9300 , n9301 );
buf ( n9303 , n5212 );
xor ( n9304 , n9302 , n9303 );
buf ( n9305 , n5213 );
xor ( n9306 , n9304 , n9305 );
xor ( n9307 , n9291 , n9306 );
and ( n9308 , n9262 , n9307 );
xor ( n9309 , n9218 , n9308 );
xor ( n9310 , n9174 , n9309 );
xor ( n9311 , n8869 , n9310 );
xor ( n9312 , n7456 , n8249 );
xor ( n9313 , n9312 , n6500 );
buf ( n9314 , n5214 );
xor ( n9315 , n9314 , n6913 );
xor ( n9316 , n9315 , n8600 );
not ( n9317 , n9316 );
buf ( n9318 , n5215 );
not ( n9319 , n6474 );
buf ( n9320 , n5215 );
and ( n9321 , n9319 , n9320 );
buf ( n9322 , n5216 );
xor ( n9323 , n9322 , n9320 );
and ( n9324 , n9323 , n6474 );
or ( n9325 , n9321 , n9324 );
not ( n9326 , n6474 );
buf ( n9327 , n5215 );
and ( n9328 , n9326 , n9327 );
buf ( n9329 , n5217 );
xor ( n9330 , n9329 , n9327 );
and ( n9331 , n9330 , n6474 );
or ( n9332 , n9328 , n9331 );
xor ( n9333 , n9325 , n9332 );
buf ( n9334 , n5218 );
xor ( n9335 , n9333 , n9334 );
buf ( n9336 , n5219 );
xor ( n9337 , n9335 , n9336 );
xor ( n9338 , n9337 , n6742 );
xor ( n9339 , n9318 , n9338 );
not ( n9340 , n6474 );
buf ( n9341 , n5220 );
and ( n9342 , n9340 , n9341 );
buf ( n9343 , n5221 );
xor ( n9344 , n9343 , n9341 );
and ( n9345 , n9344 , n6474 );
or ( n9346 , n9342 , n9345 );
buf ( n9347 , n5222 );
xor ( n9348 , n9346 , n9347 );
buf ( n9349 , n5223 );
xor ( n9350 , n9348 , n9349 );
buf ( n9351 , n5224 );
xor ( n9352 , n9350 , n9351 );
buf ( n9353 , n5225 );
xor ( n9354 , n9352 , n9353 );
xor ( n9355 , n9339 , n9354 );
and ( n9356 , n9317 , n9355 );
xor ( n9357 , n9313 , n9356 );
not ( n9358 , n6474 );
buf ( n9359 , n5226 );
and ( n9360 , n9358 , n9359 );
buf ( n9361 , n5227 );
xor ( n9362 , n9361 , n9359 );
and ( n9363 , n9362 , n6474 );
or ( n9364 , n9360 , n9363 );
not ( n9365 , n6474 );
buf ( n9366 , n5228 );
and ( n9367 , n9365 , n9366 );
buf ( n9368 , n5229 );
xor ( n9369 , n9368 , n9366 );
and ( n9370 , n9369 , n6474 );
or ( n9371 , n9367 , n9370 );
xor ( n9372 , n9364 , n9371 );
buf ( n9373 , n5230 );
xor ( n9374 , n9372 , n9373 );
buf ( n9375 , n5231 );
xor ( n9376 , n9374 , n9375 );
buf ( n9377 , n5232 );
xor ( n9378 , n9376 , n9377 );
xor ( n9379 , n8528 , n9378 );
not ( n9380 , n6474 );
buf ( n9381 , n5233 );
and ( n9382 , n9380 , n9381 );
buf ( n9383 , n5234 );
xor ( n9384 , n9383 , n9381 );
and ( n9385 , n9384 , n6474 );
or ( n9386 , n9382 , n9385 );
not ( n9387 , n6474 );
buf ( n9388 , n5235 );
and ( n9389 , n9387 , n9388 );
buf ( n9390 , n5236 );
xor ( n9391 , n9390 , n9388 );
and ( n9392 , n9391 , n6474 );
or ( n9393 , n9389 , n9392 );
xor ( n9394 , n9386 , n9393 );
buf ( n9395 , n5237 );
xor ( n9396 , n9394 , n9395 );
buf ( n9397 , n5238 );
xor ( n9398 , n9396 , n9397 );
buf ( n9399 , n5239 );
xor ( n9400 , n9398 , n9399 );
xor ( n9401 , n9379 , n9400 );
buf ( n9402 , n5240 );
not ( n9403 , n6474 );
buf ( n9404 , n5241 );
and ( n9405 , n9403 , n9404 );
buf ( n9406 , n5242 );
xor ( n9407 , n9406 , n9404 );
and ( n9408 , n9407 , n6474 );
or ( n9409 , n9405 , n9408 );
buf ( n9410 , n5243 );
xor ( n9411 , n9409 , n9410 );
buf ( n9412 , n5244 );
xor ( n9413 , n9411 , n9412 );
buf ( n9414 , n5245 );
xor ( n9415 , n9413 , n9414 );
buf ( n9416 , n5246 );
xor ( n9417 , n9415 , n9416 );
xor ( n9418 , n9402 , n9417 );
not ( n9419 , n6474 );
buf ( n9420 , n5247 );
and ( n9421 , n9419 , n9420 );
buf ( n9422 , n5248 );
xor ( n9423 , n9422 , n9420 );
and ( n9424 , n9423 , n6474 );
or ( n9425 , n9421 , n9424 );
not ( n9426 , n6474 );
buf ( n9427 , n5249 );
and ( n9428 , n9426 , n9427 );
buf ( n9429 , n5250 );
xor ( n9430 , n9429 , n9427 );
and ( n9431 , n9430 , n6474 );
or ( n9432 , n9428 , n9431 );
xor ( n9433 , n9425 , n9432 );
buf ( n9434 , n5251 );
xor ( n9435 , n9433 , n9434 );
buf ( n9436 , n5252 );
xor ( n9437 , n9435 , n9436 );
buf ( n9438 , n5253 );
xor ( n9439 , n9437 , n9438 );
xor ( n9440 , n9418 , n9439 );
not ( n9441 , n9440 );
buf ( n9442 , n5254 );
xor ( n9443 , n9442 , n8622 );
not ( n9444 , n6474 );
buf ( n9445 , n5255 );
and ( n9446 , n9444 , n9445 );
buf ( n9447 , n5256 );
xor ( n9448 , n9447 , n9445 );
and ( n9449 , n9448 , n6474 );
or ( n9450 , n9446 , n9449 );
not ( n9451 , n6474 );
buf ( n9452 , n5257 );
and ( n9453 , n9451 , n9452 );
buf ( n9454 , n5258 );
xor ( n9455 , n9454 , n9452 );
and ( n9456 , n9455 , n6474 );
or ( n9457 , n9453 , n9456 );
xor ( n9458 , n9450 , n9457 );
buf ( n9459 , n5259 );
xor ( n9460 , n9458 , n9459 );
buf ( n9461 , n5260 );
xor ( n9462 , n9460 , n9461 );
buf ( n9463 , n5261 );
xor ( n9464 , n9462 , n9463 );
xor ( n9465 , n9443 , n9464 );
and ( n9466 , n9441 , n9465 );
xor ( n9467 , n9401 , n9466 );
xor ( n9468 , n9357 , n9467 );
not ( n9469 , n6474 );
buf ( n9470 , n5262 );
and ( n9471 , n9469 , n9470 );
buf ( n9472 , n5263 );
xor ( n9473 , n9472 , n9470 );
and ( n9474 , n9473 , n6474 );
or ( n9475 , n9471 , n9474 );
not ( n9476 , n6474 );
buf ( n9477 , n5264 );
and ( n9478 , n9476 , n9477 );
buf ( n9479 , n5265 );
xor ( n9480 , n9479 , n9477 );
and ( n9481 , n9480 , n6474 );
or ( n9482 , n9478 , n9481 );
xor ( n9483 , n9475 , n9482 );
buf ( n9484 , n5266 );
xor ( n9485 , n9483 , n9484 );
buf ( n9486 , n5267 );
xor ( n9487 , n9485 , n9486 );
buf ( n9488 , n5268 );
xor ( n9489 , n9487 , n9488 );
xor ( n9490 , n6732 , n9489 );
not ( n9491 , n6474 );
buf ( n9492 , n5269 );
and ( n9493 , n9491 , n9492 );
buf ( n9494 , n5270 );
xor ( n9495 , n9494 , n9492 );
and ( n9496 , n9495 , n6474 );
or ( n9497 , n9493 , n9496 );
not ( n9498 , n6474 );
buf ( n9499 , n5271 );
and ( n9500 , n9498 , n9499 );
buf ( n9501 , n5272 );
xor ( n9502 , n9501 , n9499 );
and ( n9503 , n9502 , n6474 );
or ( n9504 , n9500 , n9503 );
xor ( n9505 , n9497 , n9504 );
buf ( n9506 , n5273 );
xor ( n9507 , n9505 , n9506 );
buf ( n9508 , n5274 );
xor ( n9509 , n9507 , n9508 );
buf ( n9510 , n5275 );
xor ( n9511 , n9509 , n9510 );
xor ( n9512 , n9490 , n9511 );
buf ( n9513 , n5276 );
not ( n9514 , n6474 );
buf ( n9515 , n5277 );
and ( n9516 , n9514 , n9515 );
buf ( n9517 , n5278 );
xor ( n9518 , n9517 , n9515 );
and ( n9519 , n9518 , n6474 );
or ( n9520 , n9516 , n9519 );
not ( n9521 , n6474 );
buf ( n9522 , n5279 );
and ( n9523 , n9521 , n9522 );
buf ( n9524 , n5280 );
xor ( n9525 , n9524 , n9522 );
and ( n9526 , n9525 , n6474 );
or ( n9527 , n9523 , n9526 );
xor ( n9528 , n9520 , n9527 );
buf ( n9529 , n5281 );
xor ( n9530 , n9528 , n9529 );
buf ( n9531 , n5282 );
xor ( n9532 , n9530 , n9531 );
buf ( n9533 , n5283 );
xor ( n9534 , n9532 , n9533 );
xor ( n9535 , n9513 , n9534 );
buf ( n9536 , n5284 );
xor ( n9537 , n9102 , n9536 );
buf ( n9538 , n5285 );
xor ( n9539 , n9537 , n9538 );
buf ( n9540 , n5286 );
xor ( n9541 , n9539 , n9540 );
buf ( n9542 , n5287 );
xor ( n9543 , n9541 , n9542 );
xor ( n9544 , n9535 , n9543 );
not ( n9545 , n9544 );
buf ( n9546 , n5288 );
not ( n9547 , n6474 );
buf ( n9548 , n5289 );
and ( n9549 , n9547 , n9548 );
buf ( n9550 , n5290 );
xor ( n9551 , n9550 , n9548 );
and ( n9552 , n9551 , n6474 );
or ( n9553 , n9549 , n9552 );
xor ( n9554 , n9553 , n8718 );
buf ( n9555 , n5291 );
xor ( n9556 , n9554 , n9555 );
buf ( n9557 , n5292 );
xor ( n9558 , n9556 , n9557 );
xor ( n9559 , n9558 , n8167 );
xor ( n9560 , n9546 , n9559 );
not ( n9561 , n6474 );
buf ( n9562 , n5293 );
and ( n9563 , n9561 , n9562 );
buf ( n9564 , n5294 );
xor ( n9565 , n9564 , n9562 );
and ( n9566 , n9565 , n6474 );
or ( n9567 , n9563 , n9566 );
not ( n9568 , n6474 );
buf ( n9569 , n5295 );
and ( n9570 , n9568 , n9569 );
buf ( n9571 , n5296 );
xor ( n9572 , n9571 , n9569 );
and ( n9573 , n9572 , n6474 );
or ( n9574 , n9570 , n9573 );
xor ( n9575 , n9567 , n9574 );
buf ( n9576 , n5297 );
xor ( n9577 , n9575 , n9576 );
buf ( n9578 , n5298 );
xor ( n9579 , n9577 , n9578 );
buf ( n9580 , n5299 );
xor ( n9581 , n9579 , n9580 );
xor ( n9582 , n9560 , n9581 );
and ( n9583 , n9545 , n9582 );
xor ( n9584 , n9512 , n9583 );
xor ( n9585 , n9468 , n9584 );
not ( n9586 , n6474 );
buf ( n9587 , n5300 );
and ( n9588 , n9586 , n9587 );
buf ( n9589 , n5301 );
xor ( n9590 , n9589 , n9587 );
and ( n9591 , n9590 , n6474 );
or ( n9592 , n9588 , n9591 );
not ( n9593 , n6474 );
buf ( n9594 , n5302 );
and ( n9595 , n9593 , n9594 );
buf ( n9596 , n5303 );
xor ( n9597 , n9596 , n9594 );
and ( n9598 , n9597 , n6474 );
or ( n9599 , n9595 , n9598 );
xor ( n9600 , n9599 , n7840 );
buf ( n9601 , n5304 );
xor ( n9602 , n9600 , n9601 );
buf ( n9603 , n5305 );
xor ( n9604 , n9602 , n9603 );
buf ( n9605 , n5306 );
xor ( n9606 , n9604 , n9605 );
xor ( n9607 , n9592 , n9606 );
not ( n9608 , n6474 );
buf ( n9609 , n5307 );
and ( n9610 , n9608 , n9609 );
buf ( n9611 , n5308 );
xor ( n9612 , n9611 , n9609 );
and ( n9613 , n9612 , n6474 );
or ( n9614 , n9610 , n9613 );
not ( n9615 , n6474 );
buf ( n9616 , n5309 );
and ( n9617 , n9615 , n9616 );
buf ( n9618 , n5310 );
xor ( n9619 , n9618 , n9616 );
and ( n9620 , n9619 , n6474 );
or ( n9621 , n9617 , n9620 );
xor ( n9622 , n9614 , n9621 );
buf ( n9623 , n5311 );
xor ( n9624 , n9622 , n9623 );
buf ( n9625 , n5312 );
xor ( n9626 , n9624 , n9625 );
buf ( n9627 , n5313 );
xor ( n9628 , n9626 , n9627 );
xor ( n9629 , n9607 , n9628 );
buf ( n9630 , n5314 );
not ( n9631 , n6474 );
buf ( n9632 , n5315 );
and ( n9633 , n9631 , n9632 );
buf ( n9634 , n5316 );
xor ( n9635 , n9634 , n9632 );
and ( n9636 , n9635 , n6474 );
or ( n9637 , n9633 , n9636 );
not ( n9638 , n6474 );
buf ( n9639 , n5317 );
and ( n9640 , n9638 , n9639 );
buf ( n9641 , n5318 );
xor ( n9642 , n9641 , n9639 );
and ( n9643 , n9642 , n6474 );
or ( n9644 , n9640 , n9643 );
xor ( n9645 , n9637 , n9644 );
buf ( n9646 , n5319 );
xor ( n9647 , n9645 , n9646 );
buf ( n9648 , n5320 );
xor ( n9649 , n9647 , n9648 );
buf ( n9650 , n5321 );
xor ( n9651 , n9649 , n9650 );
xor ( n9652 , n9630 , n9651 );
not ( n9653 , n6474 );
buf ( n9654 , n5322 );
and ( n9655 , n9653 , n9654 );
buf ( n9656 , n5323 );
xor ( n9657 , n9656 , n9654 );
and ( n9658 , n9657 , n6474 );
or ( n9659 , n9655 , n9658 );
not ( n9660 , n6474 );
buf ( n9661 , n5324 );
and ( n9662 , n9660 , n9661 );
buf ( n9663 , n5325 );
xor ( n9664 , n9663 , n9661 );
and ( n9665 , n9664 , n6474 );
or ( n9666 , n9662 , n9665 );
xor ( n9667 , n9659 , n9666 );
buf ( n9668 , n5326 );
xor ( n9669 , n9667 , n9668 );
buf ( n9670 , n5327 );
xor ( n9671 , n9669 , n9670 );
buf ( n9672 , n5328 );
xor ( n9673 , n9671 , n9672 );
xor ( n9674 , n9652 , n9673 );
not ( n9675 , n9674 );
buf ( n9676 , n5329 );
xor ( n9677 , n9676 , n8696 );
xor ( n9678 , n9677 , n8710 );
and ( n9679 , n9675 , n9678 );
xor ( n9680 , n9629 , n9679 );
xor ( n9681 , n9585 , n9680 );
not ( n9682 , n6474 );
buf ( n9683 , n5330 );
and ( n9684 , n9682 , n9683 );
buf ( n9685 , n5331 );
xor ( n9686 , n9685 , n9683 );
and ( n9687 , n9686 , n6474 );
or ( n9688 , n9684 , n9687 );
xor ( n9689 , n9688 , n9079 );
xor ( n9690 , n9689 , n9094 );
buf ( n9691 , n5332 );
xor ( n9692 , n9691 , n7208 );
xor ( n9693 , n9692 , n7230 );
not ( n9694 , n9693 );
buf ( n9695 , n5333 );
not ( n9696 , n6474 );
buf ( n9697 , n5334 );
and ( n9698 , n9696 , n9697 );
buf ( n9699 , n5335 );
xor ( n9700 , n9699 , n9697 );
and ( n9701 , n9700 , n6474 );
or ( n9702 , n9698 , n9701 );
buf ( n9703 , n5336 );
xor ( n9704 , n9702 , n9703 );
buf ( n9705 , n5337 );
xor ( n9706 , n9704 , n9705 );
buf ( n9707 , n5338 );
xor ( n9708 , n9706 , n9707 );
buf ( n9709 , n5339 );
xor ( n9710 , n9708 , n9709 );
xor ( n9711 , n9695 , n9710 );
not ( n9712 , n6474 );
buf ( n9713 , n5340 );
and ( n9714 , n9712 , n9713 );
buf ( n9715 , n5341 );
xor ( n9716 , n9715 , n9713 );
and ( n9717 , n9716 , n6474 );
or ( n9718 , n9714 , n9717 );
not ( n9719 , n6474 );
buf ( n9720 , n5342 );
and ( n9721 , n9719 , n9720 );
buf ( n9722 , n5343 );
xor ( n9723 , n9722 , n9720 );
and ( n9724 , n9723 , n6474 );
or ( n9725 , n9721 , n9724 );
xor ( n9726 , n9718 , n9725 );
buf ( n9727 , n5344 );
xor ( n9728 , n9726 , n9727 );
buf ( n9729 , n5345 );
xor ( n9730 , n9728 , n9729 );
buf ( n9731 , n5346 );
xor ( n9732 , n9730 , n9731 );
xor ( n9733 , n9711 , n9732 );
and ( n9734 , n9694 , n9733 );
xor ( n9735 , n9690 , n9734 );
xor ( n9736 , n9681 , n9735 );
xor ( n9737 , n9311 , n9736 );
and ( n9738 , n8770 , n9737 );
xor ( n9739 , n7747 , n9738 );
and ( n9740 , n9739 , n6475 );
or ( n9741 , n6478 , n9740 );
and ( n9742 , n6470 , n9741 );
buf ( n9743 , n9742 );
buf ( n9744 , n9743 );
not ( n9745 , n6469 );
not ( n9746 , n6475 );
buf ( n9747 , n5347 );
and ( n9748 , n9746 , n9747 );
buf ( n9749 , n5348 );
not ( n9750 , n6474 );
buf ( n9751 , n5349 );
and ( n9752 , n9750 , n9751 );
buf ( n9753 , n5350 );
xor ( n9754 , n9753 , n9751 );
and ( n9755 , n9754 , n6474 );
or ( n9756 , n9752 , n9755 );
not ( n9757 , n6474 );
buf ( n9758 , n5351 );
and ( n9759 , n9757 , n9758 );
buf ( n9760 , n5352 );
xor ( n9761 , n9760 , n9758 );
and ( n9762 , n9761 , n6474 );
or ( n9763 , n9759 , n9762 );
xor ( n9764 , n9756 , n9763 );
buf ( n9765 , n5353 );
xor ( n9766 , n9764 , n9765 );
buf ( n9767 , n5354 );
xor ( n9768 , n9766 , n9767 );
buf ( n9769 , n5355 );
xor ( n9770 , n9768 , n9769 );
xor ( n9771 , n9749 , n9770 );
xor ( n9772 , n9771 , n7112 );
buf ( n9773 , n5356 );
not ( n9774 , n6474 );
buf ( n9775 , n5357 );
and ( n9776 , n9774 , n9775 );
buf ( n9777 , n5358 );
xor ( n9778 , n9777 , n9775 );
and ( n9779 , n9778 , n6474 );
or ( n9780 , n9776 , n9779 );
not ( n9781 , n6474 );
buf ( n9782 , n5359 );
and ( n9783 , n9781 , n9782 );
buf ( n9784 , n5360 );
xor ( n9785 , n9784 , n9782 );
and ( n9786 , n9785 , n6474 );
or ( n9787 , n9783 , n9786 );
xor ( n9788 , n9780 , n9787 );
buf ( n9789 , n5361 );
xor ( n9790 , n9788 , n9789 );
buf ( n9791 , n5362 );
xor ( n9792 , n9790 , n9791 );
buf ( n9793 , n5363 );
xor ( n9794 , n9792 , n9793 );
xor ( n9795 , n9773 , n9794 );
not ( n9796 , n6474 );
buf ( n9797 , n5364 );
and ( n9798 , n9796 , n9797 );
buf ( n9799 , n5365 );
xor ( n9800 , n9799 , n9797 );
and ( n9801 , n9800 , n6474 );
or ( n9802 , n9798 , n9801 );
not ( n9803 , n6474 );
buf ( n9804 , n5366 );
and ( n9805 , n9803 , n9804 );
buf ( n9806 , n5367 );
xor ( n9807 , n9806 , n9804 );
and ( n9808 , n9807 , n6474 );
or ( n9809 , n9805 , n9808 );
xor ( n9810 , n9802 , n9809 );
buf ( n9811 , n5368 );
xor ( n9812 , n9810 , n9811 );
buf ( n9813 , n5369 );
xor ( n9814 , n9812 , n9813 );
buf ( n9815 , n5370 );
xor ( n9816 , n9814 , n9815 );
xor ( n9817 , n9795 , n9816 );
not ( n9818 , n9817 );
xor ( n9819 , n8763 , n8269 );
xor ( n9820 , n9819 , n8291 );
and ( n9821 , n9818 , n9820 );
xor ( n9822 , n9772 , n9821 );
not ( n9823 , n6474 );
buf ( n9824 , n5371 );
and ( n9825 , n9823 , n9824 );
buf ( n9826 , n5372 );
xor ( n9827 , n9826 , n9824 );
and ( n9828 , n9827 , n6474 );
or ( n9829 , n9825 , n9828 );
not ( n9830 , n6474 );
buf ( n9831 , n5373 );
and ( n9832 , n9830 , n9831 );
buf ( n9833 , n5374 );
xor ( n9834 , n9833 , n9831 );
and ( n9835 , n9834 , n6474 );
or ( n9836 , n9832 , n9835 );
not ( n9837 , n6474 );
buf ( n9838 , n5375 );
and ( n9839 , n9837 , n9838 );
buf ( n9840 , n5376 );
xor ( n9841 , n9840 , n9838 );
and ( n9842 , n9841 , n6474 );
or ( n9843 , n9839 , n9842 );
xor ( n9844 , n9836 , n9843 );
buf ( n9845 , n5377 );
xor ( n9846 , n9844 , n9845 );
buf ( n9847 , n5378 );
xor ( n9848 , n9846 , n9847 );
buf ( n9849 , n5379 );
xor ( n9850 , n9848 , n9849 );
xor ( n9851 , n9829 , n9850 );
not ( n9852 , n6474 );
buf ( n9853 , n5380 );
and ( n9854 , n9852 , n9853 );
buf ( n9855 , n5381 );
xor ( n9856 , n9855 , n9853 );
and ( n9857 , n9856 , n6474 );
or ( n9858 , n9854 , n9857 );
not ( n9859 , n6474 );
buf ( n9860 , n5382 );
and ( n9861 , n9859 , n9860 );
buf ( n9862 , n5383 );
xor ( n9863 , n9862 , n9860 );
and ( n9864 , n9863 , n6474 );
or ( n9865 , n9861 , n9864 );
xor ( n9866 , n9858 , n9865 );
buf ( n9867 , n5384 );
xor ( n9868 , n9866 , n9867 );
buf ( n9869 , n5385 );
xor ( n9870 , n9868 , n9869 );
buf ( n9871 , n5386 );
xor ( n9872 , n9870 , n9871 );
xor ( n9873 , n9851 , n9872 );
xor ( n9874 , n8154 , n8414 );
xor ( n9875 , n9874 , n9026 );
not ( n9876 , n9875 );
buf ( n9877 , n5387 );
not ( n9878 , n6474 );
and ( n9879 , n9878 , n9747 );
buf ( n9880 , n5388 );
xor ( n9881 , n9880 , n9747 );
and ( n9882 , n9881 , n6474 );
or ( n9883 , n9879 , n9882 );
not ( n9884 , n6474 );
buf ( n9885 , n5389 );
and ( n9886 , n9884 , n9885 );
buf ( n9887 , n5390 );
xor ( n9888 , n9887 , n9885 );
and ( n9889 , n9888 , n6474 );
or ( n9890 , n9886 , n9889 );
xor ( n9891 , n9883 , n9890 );
xor ( n9892 , n9891 , n8426 );
buf ( n9893 , n5391 );
xor ( n9894 , n9892 , n9893 );
xor ( n9895 , n9894 , n8977 );
xor ( n9896 , n9877 , n9895 );
xor ( n9897 , n9896 , n7612 );
and ( n9898 , n9876 , n9897 );
xor ( n9899 , n9873 , n9898 );
buf ( n9900 , n5392 );
not ( n9901 , n6474 );
buf ( n9902 , n5393 );
and ( n9903 , n9901 , n9902 );
buf ( n9904 , n5394 );
xor ( n9905 , n9904 , n9902 );
and ( n9906 , n9905 , n6474 );
or ( n9907 , n9903 , n9906 );
not ( n9908 , n6474 );
buf ( n9909 , n5395 );
and ( n9910 , n9908 , n9909 );
buf ( n9911 , n5396 );
xor ( n9912 , n9911 , n9909 );
and ( n9913 , n9912 , n6474 );
or ( n9914 , n9910 , n9913 );
xor ( n9915 , n9907 , n9914 );
buf ( n9916 , n5397 );
xor ( n9917 , n9915 , n9916 );
buf ( n9918 , n5398 );
xor ( n9919 , n9917 , n9918 );
buf ( n9920 , n5399 );
xor ( n9921 , n9919 , n9920 );
xor ( n9922 , n9900 , n9921 );
not ( n9923 , n6474 );
buf ( n9924 , n5400 );
and ( n9925 , n9923 , n9924 );
buf ( n9926 , n5401 );
xor ( n9927 , n9926 , n9924 );
and ( n9928 , n9927 , n6474 );
or ( n9929 , n9925 , n9928 );
not ( n9930 , n6474 );
and ( n9931 , n9930 , n6477 );
buf ( n9932 , n5402 );
xor ( n9933 , n9932 , n6477 );
and ( n9934 , n9933 , n6474 );
or ( n9935 , n9931 , n9934 );
xor ( n9936 , n9929 , n9935 );
buf ( n9937 , n5403 );
xor ( n9938 , n9936 , n9937 );
buf ( n9939 , n5404 );
xor ( n9940 , n9938 , n9939 );
buf ( n9941 , n5405 );
xor ( n9942 , n9940 , n9941 );
xor ( n9943 , n9922 , n9942 );
buf ( n9944 , n5406 );
xor ( n9945 , n9944 , n6891 );
xor ( n9946 , n9945 , n6913 );
not ( n9947 , n9946 );
buf ( n9948 , n5407 );
xor ( n9949 , n9948 , n9047 );
xor ( n9950 , n9949 , n9338 );
and ( n9951 , n9947 , n9950 );
xor ( n9952 , n9943 , n9951 );
xor ( n9953 , n9899 , n9952 );
not ( n9954 , n6474 );
buf ( n9955 , n5408 );
and ( n9956 , n9954 , n9955 );
buf ( n9957 , n5409 );
xor ( n9958 , n9957 , n9955 );
and ( n9959 , n9958 , n6474 );
or ( n9960 , n9956 , n9959 );
not ( n9961 , n6474 );
buf ( n9962 , n5410 );
and ( n9963 , n9961 , n9962 );
buf ( n9964 , n5411 );
xor ( n9965 , n9964 , n9962 );
and ( n9966 , n9965 , n6474 );
or ( n9967 , n9963 , n9966 );
xor ( n9968 , n9960 , n9967 );
buf ( n9969 , n5412 );
xor ( n9970 , n9968 , n9969 );
xor ( n9971 , n9970 , n9442 );
buf ( n9972 , n5413 );
xor ( n9973 , n9971 , n9972 );
xor ( n9974 , n6493 , n9973 );
not ( n9975 , n6474 );
buf ( n9976 , n5414 );
and ( n9977 , n9975 , n9976 );
buf ( n9978 , n5415 );
xor ( n9979 , n9978 , n9976 );
and ( n9980 , n9979 , n6474 );
or ( n9981 , n9977 , n9980 );
not ( n9982 , n6474 );
buf ( n9983 , n5416 );
and ( n9984 , n9982 , n9983 );
buf ( n9985 , n5417 );
xor ( n9986 , n9985 , n9983 );
and ( n9987 , n9986 , n6474 );
or ( n9988 , n9984 , n9987 );
xor ( n9989 , n9981 , n9988 );
buf ( n9990 , n5418 );
xor ( n9991 , n9989 , n9990 );
buf ( n9992 , n5419 );
xor ( n9993 , n9991 , n9992 );
buf ( n9994 , n5420 );
xor ( n9995 , n9993 , n9994 );
xor ( n9996 , n9974 , n9995 );
not ( n9997 , n9772 );
and ( n9998 , n9997 , n9817 );
xor ( n9999 , n9996 , n9998 );
xor ( n10000 , n9953 , n9999 );
not ( n10001 , n6474 );
buf ( n10002 , n5421 );
and ( n10003 , n10001 , n10002 );
buf ( n10004 , n5422 );
xor ( n10005 , n10004 , n10002 );
and ( n10006 , n10005 , n6474 );
or ( n10007 , n10003 , n10006 );
not ( n10008 , n6474 );
buf ( n10009 , n5423 );
and ( n10010 , n10008 , n10009 );
buf ( n10011 , n5424 );
xor ( n10012 , n10011 , n10009 );
and ( n10013 , n10012 , n6474 );
or ( n10014 , n10010 , n10013 );
buf ( n10015 , n5425 );
xor ( n10016 , n10014 , n10015 );
buf ( n10017 , n5426 );
xor ( n10018 , n10016 , n10017 );
buf ( n10019 , n5427 );
xor ( n10020 , n10018 , n10019 );
buf ( n10021 , n5428 );
xor ( n10022 , n10020 , n10021 );
xor ( n10023 , n10007 , n10022 );
not ( n10024 , n6474 );
buf ( n10025 , n5429 );
and ( n10026 , n10024 , n10025 );
buf ( n10027 , n5430 );
xor ( n10028 , n10027 , n10025 );
and ( n10029 , n10028 , n6474 );
or ( n10030 , n10026 , n10029 );
not ( n10031 , n6474 );
buf ( n10032 , n5431 );
and ( n10033 , n10031 , n10032 );
buf ( n10034 , n5432 );
xor ( n10035 , n10034 , n10032 );
and ( n10036 , n10035 , n6474 );
or ( n10037 , n10033 , n10036 );
xor ( n10038 , n10030 , n10037 );
buf ( n10039 , n5433 );
xor ( n10040 , n10038 , n10039 );
buf ( n10041 , n5434 );
xor ( n10042 , n10040 , n10041 );
buf ( n10043 , n5435 );
xor ( n10044 , n10042 , n10043 );
xor ( n10045 , n10023 , n10044 );
buf ( n10046 , n5436 );
not ( n10047 , n6474 );
buf ( n10048 , n5437 );
and ( n10049 , n10047 , n10048 );
buf ( n10050 , n5438 );
xor ( n10051 , n10050 , n10048 );
and ( n10052 , n10051 , n6474 );
or ( n10053 , n10049 , n10052 );
not ( n10054 , n6474 );
buf ( n10055 , n5439 );
and ( n10056 , n10054 , n10055 );
buf ( n10057 , n5440 );
xor ( n10058 , n10057 , n10055 );
and ( n10059 , n10058 , n6474 );
or ( n10060 , n10056 , n10059 );
xor ( n10061 , n10053 , n10060 );
buf ( n10062 , n5441 );
xor ( n10063 , n10061 , n10062 );
buf ( n10064 , n5442 );
xor ( n10065 , n10063 , n10064 );
buf ( n10066 , n5443 );
xor ( n10067 , n10065 , n10066 );
xor ( n10068 , n10046 , n10067 );
not ( n10069 , n6474 );
buf ( n10070 , n5444 );
and ( n10071 , n10069 , n10070 );
buf ( n10072 , n5445 );
xor ( n10073 , n10072 , n10070 );
and ( n10074 , n10073 , n6474 );
or ( n10075 , n10071 , n10074 );
not ( n10076 , n6474 );
buf ( n10077 , n5446 );
and ( n10078 , n10076 , n10077 );
buf ( n10079 , n5447 );
xor ( n10080 , n10079 , n10077 );
and ( n10081 , n10080 , n6474 );
or ( n10082 , n10078 , n10081 );
xor ( n10083 , n10075 , n10082 );
buf ( n10084 , n5448 );
xor ( n10085 , n10083 , n10084 );
buf ( n10086 , n5449 );
xor ( n10087 , n10085 , n10086 );
buf ( n10088 , n5450 );
xor ( n10089 , n10087 , n10088 );
xor ( n10090 , n10068 , n10089 );
not ( n10091 , n10090 );
xor ( n10092 , n9287 , n8660 );
not ( n10093 , n6474 );
buf ( n10094 , n5451 );
and ( n10095 , n10093 , n10094 );
buf ( n10096 , n5452 );
xor ( n10097 , n10096 , n10094 );
and ( n10098 , n10097 , n6474 );
or ( n10099 , n10095 , n10098 );
xor ( n10100 , n10099 , n9688 );
buf ( n10101 , n5453 );
xor ( n10102 , n10100 , n10101 );
buf ( n10103 , n5454 );
xor ( n10104 , n10102 , n10103 );
xor ( n10105 , n10104 , n9058 );
xor ( n10106 , n10092 , n10105 );
and ( n10107 , n10091 , n10106 );
xor ( n10108 , n10045 , n10107 );
xor ( n10109 , n10000 , n10108 );
not ( n10110 , n6474 );
buf ( n10111 , n5455 );
and ( n10112 , n10110 , n10111 );
buf ( n10113 , n5456 );
xor ( n10114 , n10113 , n10111 );
and ( n10115 , n10114 , n6474 );
or ( n10116 , n10112 , n10115 );
not ( n10117 , n6474 );
buf ( n10118 , n5457 );
and ( n10119 , n10117 , n10118 );
buf ( n10120 , n5458 );
xor ( n10121 , n10120 , n10118 );
and ( n10122 , n10121 , n6474 );
or ( n10123 , n10119 , n10122 );
xor ( n10124 , n10116 , n10123 );
buf ( n10125 , n5459 );
xor ( n10126 , n10124 , n10125 );
buf ( n10127 , n5460 );
xor ( n10128 , n10126 , n10127 );
buf ( n10129 , n5461 );
xor ( n10130 , n10128 , n10129 );
xor ( n10131 , n7941 , n10130 );
not ( n10132 , n6474 );
buf ( n10133 , n5462 );
and ( n10134 , n10132 , n10133 );
buf ( n10135 , n5463 );
xor ( n10136 , n10135 , n10133 );
and ( n10137 , n10136 , n6474 );
or ( n10138 , n10134 , n10137 );
buf ( n10139 , n5464 );
xor ( n10140 , n10138 , n10139 );
buf ( n10141 , n5465 );
xor ( n10142 , n10140 , n10141 );
buf ( n10143 , n5466 );
xor ( n10144 , n10142 , n10143 );
buf ( n10145 , n5467 );
xor ( n10146 , n10144 , n10145 );
xor ( n10147 , n10131 , n10146 );
buf ( n10148 , n5468 );
xor ( n10149 , n10148 , n7793 );
not ( n10150 , n6474 );
buf ( n10151 , n5469 );
and ( n10152 , n10150 , n10151 );
buf ( n10153 , n5470 );
xor ( n10154 , n10153 , n10151 );
and ( n10155 , n10154 , n6474 );
or ( n10156 , n10152 , n10155 );
not ( n10157 , n6474 );
buf ( n10158 , n5471 );
and ( n10159 , n10157 , n10158 );
buf ( n10160 , n5472 );
xor ( n10161 , n10160 , n10158 );
and ( n10162 , n10161 , n6474 );
or ( n10163 , n10159 , n10162 );
xor ( n10164 , n10156 , n10163 );
buf ( n10165 , n5473 );
xor ( n10166 , n10164 , n10165 );
buf ( n10167 , n5474 );
xor ( n10168 , n10166 , n10167 );
buf ( n10169 , n5475 );
xor ( n10170 , n10168 , n10169 );
xor ( n10171 , n10149 , n10170 );
not ( n10172 , n10171 );
buf ( n10173 , n5476 );
xor ( n10174 , n10173 , n7994 );
xor ( n10175 , n10174 , n8016 );
and ( n10176 , n10172 , n10175 );
xor ( n10177 , n10147 , n10176 );
xor ( n10178 , n10109 , n10177 );
xor ( n10179 , n9822 , n10178 );
not ( n10180 , n6474 );
buf ( n10181 , n5477 );
and ( n10182 , n10180 , n10181 );
buf ( n10183 , n5478 );
xor ( n10184 , n10183 , n10181 );
and ( n10185 , n10184 , n6474 );
or ( n10186 , n10182 , n10185 );
xor ( n10187 , n9225 , n10186 );
buf ( n10188 , n5479 );
xor ( n10189 , n10187 , n10188 );
buf ( n10190 , n5480 );
xor ( n10191 , n10189 , n10190 );
buf ( n10192 , n5481 );
xor ( n10193 , n10191 , n10192 );
xor ( n10194 , n8466 , n10193 );
not ( n10195 , n6474 );
buf ( n10196 , n5482 );
and ( n10197 , n10195 , n10196 );
buf ( n10198 , n5483 );
xor ( n10199 , n10198 , n10196 );
and ( n10200 , n10199 , n6474 );
or ( n10201 , n10197 , n10200 );
buf ( n10202 , n5484 );
xor ( n10203 , n10201 , n10202 );
buf ( n10204 , n5485 );
xor ( n10205 , n10203 , n10204 );
buf ( n10206 , n5486 );
xor ( n10207 , n10205 , n10206 );
buf ( n10208 , n5487 );
xor ( n10209 , n10207 , n10208 );
xor ( n10210 , n10194 , n10209 );
not ( n10211 , n6474 );
buf ( n10212 , n5488 );
and ( n10213 , n10211 , n10212 );
buf ( n10214 , n5489 );
xor ( n10215 , n10214 , n10212 );
and ( n10216 , n10215 , n6474 );
or ( n10217 , n10213 , n10216 );
xor ( n10218 , n10217 , n9269 );
buf ( n10219 , n5490 );
xor ( n10220 , n10218 , n10219 );
buf ( n10221 , n5491 );
xor ( n10222 , n10220 , n10221 );
buf ( n10223 , n5492 );
xor ( n10224 , n10222 , n10223 );
xor ( n10225 , n7375 , n10224 );
not ( n10226 , n6474 );
buf ( n10227 , n5493 );
and ( n10228 , n10226 , n10227 );
buf ( n10229 , n5494 );
xor ( n10230 , n10229 , n10227 );
and ( n10231 , n10230 , n6474 );
or ( n10232 , n10228 , n10231 );
not ( n10233 , n6474 );
buf ( n10234 , n5495 );
and ( n10235 , n10233 , n10234 );
buf ( n10236 , n5496 );
xor ( n10237 , n10236 , n10234 );
and ( n10238 , n10237 , n6474 );
or ( n10239 , n10235 , n10238 );
xor ( n10240 , n10232 , n10239 );
buf ( n10241 , n5497 );
xor ( n10242 , n10240 , n10241 );
buf ( n10243 , n5498 );
xor ( n10244 , n10242 , n10243 );
buf ( n10245 , n5499 );
xor ( n10246 , n10244 , n10245 );
xor ( n10247 , n10225 , n10246 );
not ( n10248 , n10247 );
not ( n10249 , n6474 );
buf ( n10250 , n5500 );
and ( n10251 , n10249 , n10250 );
buf ( n10252 , n5501 );
xor ( n10253 , n10252 , n10250 );
and ( n10254 , n10253 , n6474 );
or ( n10255 , n10251 , n10254 );
buf ( n10256 , n5502 );
xor ( n10257 , n10255 , n10256 );
buf ( n10258 , n5503 );
xor ( n10259 , n10257 , n10258 );
buf ( n10260 , n5504 );
xor ( n10261 , n10259 , n10260 );
buf ( n10262 , n5505 );
xor ( n10263 , n10261 , n10262 );
xor ( n10264 , n7216 , n10263 );
not ( n10265 , n6474 );
buf ( n10266 , n5506 );
and ( n10267 , n10265 , n10266 );
buf ( n10268 , n5507 );
xor ( n10269 , n10268 , n10266 );
and ( n10270 , n10269 , n6474 );
or ( n10271 , n10267 , n10270 );
not ( n10272 , n6474 );
buf ( n10273 , n5508 );
and ( n10274 , n10272 , n10273 );
buf ( n10275 , n5509 );
xor ( n10276 , n10275 , n10273 );
and ( n10277 , n10276 , n6474 );
or ( n10278 , n10274 , n10277 );
xor ( n10279 , n10271 , n10278 );
buf ( n10280 , n5510 );
xor ( n10281 , n10279 , n10280 );
buf ( n10282 , n5511 );
xor ( n10283 , n10281 , n10282 );
buf ( n10284 , n5512 );
xor ( n10285 , n10283 , n10284 );
xor ( n10286 , n10264 , n10285 );
and ( n10287 , n10248 , n10286 );
xor ( n10288 , n10210 , n10287 );
xor ( n10289 , n6760 , n9400 );
not ( n10290 , n6474 );
buf ( n10291 , n5513 );
and ( n10292 , n10290 , n10291 );
buf ( n10293 , n5514 );
xor ( n10294 , n10293 , n10291 );
and ( n10295 , n10294 , n6474 );
or ( n10296 , n10292 , n10295 );
not ( n10297 , n6474 );
buf ( n10298 , n5515 );
and ( n10299 , n10297 , n10298 );
buf ( n10300 , n5516 );
xor ( n10301 , n10300 , n10298 );
and ( n10302 , n10301 , n6474 );
or ( n10303 , n10299 , n10302 );
xor ( n10304 , n10296 , n10303 );
buf ( n10305 , n5517 );
xor ( n10306 , n10304 , n10305 );
buf ( n10307 , n5518 );
xor ( n10308 , n10306 , n10307 );
xor ( n10309 , n10308 , n7288 );
xor ( n10310 , n10289 , n10309 );
xor ( n10311 , n7909 , n9628 );
xor ( n10312 , n10311 , n6538 );
not ( n10313 , n10312 );
not ( n10314 , n6474 );
buf ( n10315 , n5519 );
and ( n10316 , n10314 , n10315 );
buf ( n10317 , n5520 );
xor ( n10318 , n10317 , n10315 );
and ( n10319 , n10318 , n6474 );
or ( n10320 , n10316 , n10319 );
not ( n10321 , n6474 );
buf ( n10322 , n5521 );
and ( n10323 , n10321 , n10322 );
buf ( n10324 , n5522 );
xor ( n10325 , n10324 , n10322 );
and ( n10326 , n10325 , n6474 );
or ( n10327 , n10323 , n10326 );
xor ( n10328 , n10320 , n10327 );
buf ( n10329 , n5523 );
xor ( n10330 , n10328 , n10329 );
buf ( n10331 , n5524 );
xor ( n10332 , n10330 , n10331 );
buf ( n10333 , n5525 );
xor ( n10334 , n10332 , n10333 );
xor ( n10335 , n6639 , n10334 );
not ( n10336 , n6474 );
buf ( n10337 , n5526 );
and ( n10338 , n10336 , n10337 );
buf ( n10339 , n5527 );
xor ( n10340 , n10339 , n10337 );
and ( n10341 , n10340 , n6474 );
or ( n10342 , n10338 , n10341 );
buf ( n10343 , n5528 );
xor ( n10344 , n10342 , n10343 );
buf ( n10345 , n5529 );
xor ( n10346 , n10344 , n10345 );
buf ( n10347 , n5530 );
xor ( n10348 , n10346 , n10347 );
buf ( n10349 , n5531 );
xor ( n10350 , n10348 , n10349 );
xor ( n10351 , n10335 , n10350 );
and ( n10352 , n10313 , n10351 );
xor ( n10353 , n10310 , n10352 );
xor ( n10354 , n10288 , n10353 );
buf ( n10355 , n5532 );
not ( n10356 , n6474 );
buf ( n10357 , n5533 );
and ( n10358 , n10356 , n10357 );
buf ( n10359 , n5534 );
xor ( n10360 , n10359 , n10357 );
and ( n10361 , n10360 , n6474 );
or ( n10362 , n10358 , n10361 );
not ( n10363 , n6474 );
buf ( n10364 , n5535 );
and ( n10365 , n10363 , n10364 );
buf ( n10366 , n5536 );
xor ( n10367 , n10366 , n10364 );
and ( n10368 , n10367 , n6474 );
or ( n10369 , n10365 , n10368 );
xor ( n10370 , n10362 , n10369 );
buf ( n10371 , n5537 );
xor ( n10372 , n10370 , n10371 );
buf ( n10373 , n5538 );
xor ( n10374 , n10372 , n10373 );
buf ( n10375 , n5539 );
xor ( n10376 , n10374 , n10375 );
xor ( n10377 , n10355 , n10376 );
xor ( n10378 , n10377 , n10067 );
buf ( n10379 , n5540 );
not ( n10380 , n6474 );
buf ( n10381 , n5541 );
and ( n10382 , n10380 , n10381 );
buf ( n10383 , n5542 );
xor ( n10384 , n10383 , n10381 );
and ( n10385 , n10384 , n6474 );
or ( n10386 , n10382 , n10385 );
buf ( n10387 , n5543 );
xor ( n10388 , n10386 , n10387 );
buf ( n10389 , n5544 );
xor ( n10390 , n10388 , n10389 );
buf ( n10391 , n5545 );
xor ( n10392 , n10390 , n10391 );
buf ( n10393 , n5546 );
xor ( n10394 , n10392 , n10393 );
xor ( n10395 , n10379 , n10394 );
not ( n10396 , n6474 );
buf ( n10397 , n5547 );
and ( n10398 , n10396 , n10397 );
buf ( n10399 , n5548 );
xor ( n10400 , n10399 , n10397 );
and ( n10401 , n10400 , n6474 );
or ( n10402 , n10398 , n10401 );
not ( n10403 , n6474 );
buf ( n10404 , n5549 );
and ( n10405 , n10403 , n10404 );
buf ( n10406 , n5550 );
xor ( n10407 , n10406 , n10404 );
and ( n10408 , n10407 , n6474 );
or ( n10409 , n10405 , n10408 );
xor ( n10410 , n10402 , n10409 );
buf ( n10411 , n5551 );
xor ( n10412 , n10410 , n10411 );
buf ( n10413 , n5552 );
xor ( n10414 , n10412 , n10413 );
buf ( n10415 , n5553 );
xor ( n10416 , n10414 , n10415 );
xor ( n10417 , n10395 , n10416 );
not ( n10418 , n10417 );
not ( n10419 , n6474 );
buf ( n10420 , n5554 );
and ( n10421 , n10419 , n10420 );
buf ( n10422 , n5555 );
xor ( n10423 , n10422 , n10420 );
and ( n10424 , n10423 , n6474 );
or ( n10425 , n10421 , n10424 );
not ( n10426 , n6474 );
buf ( n10427 , n5556 );
and ( n10428 , n10426 , n10427 );
buf ( n10429 , n5557 );
xor ( n10430 , n10429 , n10427 );
and ( n10431 , n10430 , n6474 );
or ( n10432 , n10428 , n10431 );
xor ( n10433 , n10425 , n10432 );
buf ( n10434 , n5558 );
xor ( n10435 , n10433 , n10434 );
xor ( n10436 , n10435 , n9695 );
buf ( n10437 , n5559 );
buf ( n10438 , n10437 );
xor ( n10439 , n10436 , n10438 );
xor ( n10440 , n10271 , n10439 );
xor ( n10441 , n10440 , n8574 );
and ( n10442 , n10418 , n10441 );
xor ( n10443 , n10378 , n10442 );
xor ( n10444 , n10354 , n10443 );
not ( n10445 , n6474 );
buf ( n10446 , n5560 );
and ( n10447 , n10445 , n10446 );
buf ( n10448 , n5561 );
xor ( n10449 , n10448 , n10446 );
and ( n10450 , n10449 , n6474 );
or ( n10451 , n10447 , n10450 );
not ( n10452 , n6474 );
buf ( n10453 , n5562 );
and ( n10454 , n10452 , n10453 );
buf ( n10455 , n5563 );
xor ( n10456 , n10455 , n10453 );
and ( n10457 , n10456 , n6474 );
or ( n10458 , n10454 , n10457 );
xor ( n10459 , n10451 , n10458 );
buf ( n10460 , n5564 );
xor ( n10461 , n10459 , n10460 );
buf ( n10462 , n5565 );
xor ( n10463 , n10461 , n10462 );
buf ( n10464 , n5566 );
xor ( n10465 , n10463 , n10464 );
xor ( n10466 , n9076 , n10465 );
xor ( n10467 , n10466 , n8743 );
not ( n10468 , n6474 );
buf ( n10469 , n5567 );
and ( n10470 , n10468 , n10469 );
buf ( n10471 , n5568 );
xor ( n10472 , n10471 , n10469 );
and ( n10473 , n10472 , n6474 );
or ( n10474 , n10470 , n10473 );
not ( n10475 , n6474 );
buf ( n10476 , n5569 );
and ( n10477 , n10475 , n10476 );
buf ( n10478 , n5570 );
xor ( n10479 , n10478 , n10476 );
and ( n10480 , n10479 , n6474 );
or ( n10481 , n10477 , n10480 );
xor ( n10482 , n10474 , n10481 );
buf ( n10483 , n5571 );
xor ( n10484 , n10482 , n10483 );
buf ( n10485 , n5572 );
xor ( n10486 , n10484 , n10485 );
buf ( n10487 , n5573 );
xor ( n10488 , n10486 , n10487 );
xor ( n10489 , n6849 , n10488 );
not ( n10490 , n6474 );
buf ( n10491 , n5574 );
and ( n10492 , n10490 , n10491 );
buf ( n10493 , n5575 );
xor ( n10494 , n10493 , n10491 );
and ( n10495 , n10494 , n6474 );
or ( n10496 , n10492 , n10495 );
buf ( n10497 , n5576 );
xor ( n10498 , n10496 , n10497 );
buf ( n10499 , n5577 );
xor ( n10500 , n10498 , n10499 );
buf ( n10501 , n5578 );
xor ( n10502 , n10500 , n10501 );
buf ( n10503 , n5579 );
xor ( n10504 , n10502 , n10503 );
xor ( n10505 , n10489 , n10504 );
not ( n10506 , n10505 );
not ( n10507 , n6474 );
buf ( n10508 , n5580 );
and ( n10509 , n10507 , n10508 );
buf ( n10510 , n5581 );
xor ( n10511 , n10510 , n10508 );
and ( n10512 , n10511 , n6474 );
or ( n10513 , n10509 , n10512 );
not ( n10514 , n6474 );
buf ( n10515 , n5582 );
and ( n10516 , n10514 , n10515 );
buf ( n10517 , n5583 );
xor ( n10518 , n10517 , n10515 );
and ( n10519 , n10518 , n6474 );
or ( n10520 , n10516 , n10519 );
xor ( n10521 , n10513 , n10520 );
buf ( n10522 , n5584 );
xor ( n10523 , n10521 , n10522 );
buf ( n10524 , n5585 );
xor ( n10525 , n10523 , n10524 );
buf ( n10526 , n5586 );
xor ( n10527 , n10525 , n10526 );
xor ( n10528 , n9409 , n10527 );
not ( n10529 , n6474 );
buf ( n10530 , n5587 );
and ( n10531 , n10529 , n10530 );
buf ( n10532 , n5588 );
xor ( n10533 , n10532 , n10530 );
and ( n10534 , n10533 , n6474 );
or ( n10535 , n10531 , n10534 );
not ( n10536 , n6474 );
buf ( n10537 , n5589 );
and ( n10538 , n10536 , n10537 );
buf ( n10539 , n5590 );
xor ( n10540 , n10539 , n10537 );
and ( n10541 , n10540 , n6474 );
or ( n10542 , n10538 , n10541 );
xor ( n10543 , n10535 , n10542 );
buf ( n10544 , n5591 );
xor ( n10545 , n10543 , n10544 );
buf ( n10546 , n5592 );
xor ( n10547 , n10545 , n10546 );
buf ( n10548 , n5593 );
xor ( n10549 , n10547 , n10548 );
xor ( n10550 , n10528 , n10549 );
and ( n10551 , n10506 , n10550 );
xor ( n10552 , n10467 , n10551 );
xor ( n10553 , n10444 , n10552 );
xor ( n10554 , n8134 , n7046 );
xor ( n10555 , n10554 , n8414 );
not ( n10556 , n6474 );
buf ( n10557 , n5594 );
and ( n10558 , n10556 , n10557 );
buf ( n10559 , n5595 );
xor ( n10560 , n10559 , n10557 );
and ( n10561 , n10560 , n6474 );
or ( n10562 , n10558 , n10561 );
not ( n10563 , n6474 );
buf ( n10564 , n5596 );
and ( n10565 , n10563 , n10564 );
buf ( n10566 , n5597 );
xor ( n10567 , n10566 , n10564 );
and ( n10568 , n10567 , n6474 );
or ( n10569 , n10565 , n10568 );
xor ( n10570 , n10562 , n10569 );
xor ( n10571 , n10570 , n9944 );
buf ( n10572 , n5598 );
xor ( n10573 , n10571 , n10572 );
xor ( n10574 , n10573 , n6875 );
xor ( n10575 , n9731 , n10574 );
not ( n10576 , n6474 );
buf ( n10577 , n5599 );
and ( n10578 , n10576 , n10577 );
buf ( n10579 , n5600 );
xor ( n10580 , n10579 , n10577 );
and ( n10581 , n10580 , n6474 );
or ( n10582 , n10578 , n10581 );
not ( n10583 , n6474 );
buf ( n10584 , n5601 );
and ( n10585 , n10583 , n10584 );
buf ( n10586 , n5602 );
xor ( n10587 , n10586 , n10584 );
and ( n10588 , n10587 , n6474 );
or ( n10589 , n10585 , n10588 );
xor ( n10590 , n10582 , n10589 );
xor ( n10591 , n10590 , n9314 );
buf ( n10592 , n5603 );
xor ( n10593 , n10591 , n10592 );
buf ( n10594 , n5604 );
xor ( n10595 , n10593 , n10594 );
xor ( n10596 , n10575 , n10595 );
not ( n10597 , n10596 );
not ( n10598 , n6474 );
buf ( n10599 , n5605 );
and ( n10600 , n10598 , n10599 );
buf ( n10601 , n5606 );
xor ( n10602 , n10601 , n10599 );
and ( n10603 , n10602 , n6474 );
or ( n10604 , n10600 , n10603 );
not ( n10605 , n6474 );
buf ( n10606 , n5607 );
and ( n10607 , n10605 , n10606 );
buf ( n10608 , n5608 );
xor ( n10609 , n10608 , n10606 );
and ( n10610 , n10609 , n6474 );
or ( n10611 , n10607 , n10610 );
not ( n10612 , n6474 );
buf ( n10613 , n5609 );
and ( n10614 , n10612 , n10613 );
buf ( n10615 , n5610 );
xor ( n10616 , n10615 , n10613 );
and ( n10617 , n10616 , n6474 );
or ( n10618 , n10614 , n10617 );
xor ( n10619 , n10611 , n10618 );
buf ( n10620 , n5611 );
xor ( n10621 , n10619 , n10620 );
buf ( n10622 , n5612 );
xor ( n10623 , n10621 , n10622 );
buf ( n10624 , n5613 );
xor ( n10625 , n10623 , n10624 );
xor ( n10626 , n10604 , n10625 );
xor ( n10627 , n10626 , n7208 );
and ( n10628 , n10597 , n10627 );
xor ( n10629 , n10555 , n10628 );
xor ( n10630 , n10553 , n10629 );
xor ( n10631 , n10179 , n10630 );
not ( n10632 , n6474 );
buf ( n10633 , n5614 );
and ( n10634 , n10632 , n10633 );
buf ( n10635 , n5615 );
xor ( n10636 , n10635 , n10633 );
and ( n10637 , n10636 , n6474 );
or ( n10638 , n10634 , n10637 );
not ( n10639 , n6474 );
buf ( n10640 , n5616 );
and ( n10641 , n10639 , n10640 );
buf ( n10642 , n5617 );
xor ( n10643 , n10642 , n10640 );
and ( n10644 , n10643 , n6474 );
or ( n10645 , n10641 , n10644 );
xor ( n10646 , n10638 , n10645 );
buf ( n10647 , n5618 );
xor ( n10648 , n10646 , n10647 );
buf ( n10649 , n5619 );
xor ( n10650 , n10648 , n10649 );
buf ( n10651 , n5620 );
xor ( n10652 , n10650 , n10651 );
xor ( n10653 , n10485 , n10652 );
not ( n10654 , n6474 );
buf ( n10655 , n5621 );
and ( n10656 , n10654 , n10655 );
buf ( n10657 , n5622 );
xor ( n10658 , n10657 , n10655 );
and ( n10659 , n10658 , n6474 );
or ( n10660 , n10656 , n10659 );
not ( n10661 , n6474 );
buf ( n10662 , n5623 );
and ( n10663 , n10661 , n10662 );
buf ( n10664 , n5624 );
xor ( n10665 , n10664 , n10662 );
and ( n10666 , n10665 , n6474 );
or ( n10667 , n10663 , n10666 );
xor ( n10668 , n10660 , n10667 );
buf ( n10669 , n5625 );
xor ( n10670 , n10668 , n10669 );
buf ( n10671 , n5626 );
xor ( n10672 , n10670 , n10671 );
buf ( n10673 , n5627 );
xor ( n10674 , n10672 , n10673 );
xor ( n10675 , n10653 , n10674 );
buf ( n10676 , n5628 );
not ( n10677 , n6474 );
buf ( n10678 , n5629 );
and ( n10679 , n10677 , n10678 );
buf ( n10680 , n5630 );
xor ( n10681 , n10680 , n10678 );
and ( n10682 , n10681 , n6474 );
or ( n10683 , n10679 , n10682 );
not ( n10684 , n6474 );
buf ( n10685 , n5631 );
and ( n10686 , n10684 , n10685 );
buf ( n10687 , n5632 );
xor ( n10688 , n10687 , n10685 );
and ( n10689 , n10688 , n6474 );
or ( n10690 , n10686 , n10689 );
xor ( n10691 , n10683 , n10690 );
buf ( n10692 , n5633 );
xor ( n10693 , n10691 , n10692 );
buf ( n10694 , n5634 );
xor ( n10695 , n10693 , n10694 );
buf ( n10696 , n5635 );
xor ( n10697 , n10695 , n10696 );
xor ( n10698 , n10676 , n10697 );
not ( n10699 , n6474 );
buf ( n10700 , n5636 );
and ( n10701 , n10699 , n10700 );
buf ( n10702 , n5637 );
xor ( n10703 , n10702 , n10700 );
and ( n10704 , n10703 , n6474 );
or ( n10705 , n10701 , n10704 );
buf ( n10706 , n5638 );
xor ( n10707 , n10705 , n10706 );
buf ( n10708 , n5639 );
xor ( n10709 , n10707 , n10708 );
buf ( n10710 , n5640 );
xor ( n10711 , n10709 , n10710 );
buf ( n10712 , n5641 );
xor ( n10713 , n10711 , n10712 );
xor ( n10714 , n10698 , n10713 );
not ( n10715 , n10714 );
and ( n10716 , n10715 , n8623 );
xor ( n10717 , n10675 , n10716 );
not ( n10718 , n6474 );
buf ( n10719 , n5642 );
and ( n10720 , n10718 , n10719 );
buf ( n10721 , n5643 );
xor ( n10722 , n10721 , n10719 );
and ( n10723 , n10722 , n6474 );
or ( n10724 , n10720 , n10723 );
xor ( n10725 , n10604 , n10724 );
buf ( n10726 , n5644 );
xor ( n10727 , n10725 , n10726 );
buf ( n10728 , n5645 );
xor ( n10729 , n10727 , n10728 );
buf ( n10730 , n5646 );
xor ( n10731 , n10729 , n10730 );
xor ( n10732 , n6535 , n10731 );
not ( n10733 , n6474 );
buf ( n10734 , n5647 );
and ( n10735 , n10733 , n10734 );
buf ( n10736 , n5648 );
xor ( n10737 , n10736 , n10734 );
and ( n10738 , n10737 , n6474 );
or ( n10739 , n10735 , n10738 );
buf ( n10740 , n5649 );
xor ( n10741 , n10739 , n10740 );
xor ( n10742 , n10741 , n9691 );
buf ( n10743 , n5650 );
xor ( n10744 , n10742 , n10743 );
xor ( n10745 , n10744 , n7187 );
xor ( n10746 , n10732 , n10745 );
not ( n10747 , n10746 );
not ( n10748 , n6474 );
buf ( n10749 , n5651 );
and ( n10750 , n10748 , n10749 );
buf ( n10751 , n5652 );
xor ( n10752 , n10751 , n10749 );
and ( n10753 , n10752 , n6474 );
or ( n10754 , n10750 , n10753 );
not ( n10755 , n6474 );
buf ( n10756 , n5653 );
and ( n10757 , n10755 , n10756 );
buf ( n10758 , n5654 );
xor ( n10759 , n10758 , n10756 );
and ( n10760 , n10759 , n6474 );
or ( n10761 , n10757 , n10760 );
xor ( n10762 , n10754 , n10761 );
buf ( n10763 , n5655 );
xor ( n10764 , n10762 , n10763 );
buf ( n10765 , n5656 );
xor ( n10766 , n10764 , n10765 );
buf ( n10767 , n5657 );
xor ( n10768 , n10766 , n10767 );
xor ( n10769 , n10145 , n10768 );
not ( n10770 , n6474 );
buf ( n10771 , n5658 );
and ( n10772 , n10770 , n10771 );
buf ( n10773 , n5659 );
xor ( n10774 , n10773 , n10771 );
and ( n10775 , n10774 , n6474 );
or ( n10776 , n10772 , n10775 );
not ( n10777 , n6474 );
buf ( n10778 , n5660 );
and ( n10779 , n10777 , n10778 );
buf ( n10780 , n5661 );
xor ( n10781 , n10780 , n10778 );
and ( n10782 , n10781 , n6474 );
or ( n10783 , n10779 , n10782 );
xor ( n10784 , n10776 , n10783 );
buf ( n10785 , n5662 );
xor ( n10786 , n10784 , n10785 );
buf ( n10787 , n5663 );
xor ( n10788 , n10786 , n10787 );
buf ( n10789 , n5664 );
xor ( n10790 , n10788 , n10789 );
xor ( n10791 , n10769 , n10790 );
and ( n10792 , n10747 , n10791 );
xor ( n10793 , n8470 , n10792 );
not ( n10794 , n6474 );
buf ( n10795 , n5665 );
and ( n10796 , n10794 , n10795 );
buf ( n10797 , n5666 );
xor ( n10798 , n10797 , n10795 );
and ( n10799 , n10798 , n6474 );
or ( n10800 , n10796 , n10799 );
not ( n10801 , n6474 );
buf ( n10802 , n5667 );
and ( n10803 , n10801 , n10802 );
buf ( n10804 , n5668 );
xor ( n10805 , n10804 , n10802 );
and ( n10806 , n10805 , n6474 );
or ( n10807 , n10803 , n10806 );
xor ( n10808 , n10800 , n10807 );
buf ( n10809 , n5669 );
xor ( n10810 , n10808 , n10809 );
buf ( n10811 , n5670 );
xor ( n10812 , n10810 , n10811 );
buf ( n10813 , n5671 );
xor ( n10814 , n10812 , n10813 );
xor ( n10815 , n7631 , n10814 );
not ( n10816 , n6474 );
buf ( n10817 , n5672 );
and ( n10818 , n10816 , n10817 );
buf ( n10819 , n5673 );
xor ( n10820 , n10819 , n10817 );
and ( n10821 , n10820 , n6474 );
or ( n10822 , n10818 , n10821 );
not ( n10823 , n6474 );
buf ( n10824 , n5674 );
and ( n10825 , n10823 , n10824 );
buf ( n10826 , n5675 );
xor ( n10827 , n10826 , n10824 );
and ( n10828 , n10827 , n6474 );
or ( n10829 , n10825 , n10828 );
xor ( n10830 , n10822 , n10829 );
buf ( n10831 , n5676 );
xor ( n10832 , n10830 , n10831 );
buf ( n10833 , n5677 );
xor ( n10834 , n10832 , n10833 );
buf ( n10835 , n5678 );
xor ( n10836 , n10834 , n10835 );
xor ( n10837 , n10815 , n10836 );
not ( n10838 , n10837 );
buf ( n10839 , n5679 );
xor ( n10840 , n10839 , n8366 );
xor ( n10841 , n10840 , n8388 );
and ( n10842 , n10838 , n10841 );
xor ( n10843 , n8537 , n10842 );
xor ( n10844 , n10793 , n10843 );
not ( n10845 , n6474 );
buf ( n10846 , n5680 );
and ( n10847 , n10845 , n10846 );
buf ( n10848 , n5681 );
xor ( n10849 , n10848 , n10846 );
and ( n10850 , n10849 , n6474 );
or ( n10851 , n10847 , n10850 );
not ( n10852 , n6474 );
buf ( n10853 , n5682 );
and ( n10854 , n10852 , n10853 );
buf ( n10855 , n5683 );
xor ( n10856 , n10855 , n10853 );
and ( n10857 , n10856 , n6474 );
or ( n10858 , n10854 , n10857 );
xor ( n10859 , n10851 , n10858 );
xor ( n10860 , n10859 , n9513 );
buf ( n10861 , n5684 );
xor ( n10862 , n10860 , n10861 );
buf ( n10863 , n5685 );
xor ( n10864 , n10862 , n10863 );
xor ( n10865 , n7250 , n10864 );
xor ( n10866 , n10865 , n7159 );
not ( n10867 , n10866 );
buf ( n10868 , n5686 );
xor ( n10869 , n10868 , n9148 );
xor ( n10870 , n10869 , n9170 );
and ( n10871 , n10867 , n10870 );
xor ( n10872 , n8576 , n10871 );
xor ( n10873 , n10844 , n10872 );
not ( n10874 , n10675 );
and ( n10875 , n10874 , n10714 );
xor ( n10876 , n8665 , n10875 );
xor ( n10877 , n10873 , n10876 );
buf ( n10878 , n5687 );
xor ( n10879 , n10878 , n10394 );
xor ( n10880 , n10879 , n10416 );
not ( n10881 , n10880 );
buf ( n10882 , n5688 );
xor ( n10883 , n10882 , n9850 );
xor ( n10884 , n10883 , n9872 );
and ( n10885 , n10881 , n10884 );
xor ( n10886 , n8765 , n10885 );
xor ( n10887 , n10877 , n10886 );
xor ( n10888 , n10717 , n10887 );
buf ( n10889 , n5689 );
xor ( n10890 , n10889 , n6850 );
xor ( n10891 , n10890 , n6872 );
xor ( n10892 , n8300 , n7537 );
not ( n10893 , n6474 );
buf ( n10894 , n5690 );
and ( n10895 , n10893 , n10894 );
buf ( n10896 , n5691 );
xor ( n10897 , n10896 , n10894 );
and ( n10898 , n10897 , n6474 );
or ( n10899 , n10895 , n10898 );
xor ( n10900 , n10899 , n9829 );
buf ( n10901 , n5692 );
xor ( n10902 , n10900 , n10901 );
buf ( n10903 , n5693 );
xor ( n10904 , n10902 , n10903 );
xor ( n10905 , n10904 , n10882 );
xor ( n10906 , n10892 , n10905 );
not ( n10907 , n10906 );
xor ( n10908 , n7627 , n10814 );
xor ( n10909 , n10908 , n10836 );
and ( n10910 , n10907 , n10909 );
xor ( n10911 , n10891 , n10910 );
buf ( n10912 , n5694 );
xor ( n10913 , n10912 , n8696 );
xor ( n10914 , n10913 , n8710 );
xor ( n10915 , n9981 , n9464 );
not ( n10916 , n6474 );
buf ( n10917 , n5695 );
and ( n10918 , n10916 , n10917 );
buf ( n10919 , n5696 );
xor ( n10920 , n10919 , n10917 );
and ( n10921 , n10920 , n6474 );
or ( n10922 , n10918 , n10921 );
buf ( n10923 , n5697 );
xor ( n10924 , n10922 , n10923 );
buf ( n10925 , n5698 );
xor ( n10926 , n10924 , n10925 );
xor ( n10927 , n10926 , n9773 );
buf ( n10928 , n5699 );
xor ( n10929 , n10927 , n10928 );
xor ( n10930 , n10915 , n10929 );
not ( n10931 , n10930 );
xor ( n10932 , n7919 , n6538 );
xor ( n10933 , n10932 , n6560 );
and ( n10934 , n10931 , n10933 );
xor ( n10935 , n10914 , n10934 );
xor ( n10936 , n10911 , n10935 );
buf ( n10937 , n5700 );
xor ( n10938 , n10937 , n9606 );
xor ( n10939 , n10938 , n9628 );
xor ( n10940 , n10899 , n9850 );
xor ( n10941 , n10940 , n9872 );
not ( n10942 , n10941 );
not ( n10943 , n6474 );
buf ( n10944 , n5701 );
and ( n10945 , n10943 , n10944 );
buf ( n10946 , n5702 );
xor ( n10947 , n10946 , n10944 );
and ( n10948 , n10947 , n6474 );
or ( n10949 , n10945 , n10948 );
not ( n10950 , n6474 );
buf ( n10951 , n5703 );
and ( n10952 , n10950 , n10951 );
buf ( n10953 , n5704 );
xor ( n10954 , n10953 , n10951 );
and ( n10955 , n10954 , n6474 );
or ( n10956 , n10952 , n10955 );
xor ( n10957 , n10949 , n10956 );
buf ( n10958 , n5705 );
xor ( n10959 , n10957 , n10958 );
buf ( n10960 , n5706 );
xor ( n10961 , n10959 , n10960 );
buf ( n10962 , n5707 );
xor ( n10963 , n10961 , n10962 );
xor ( n10964 , n8858 , n10963 );
xor ( n10965 , n10964 , n10864 );
and ( n10966 , n10942 , n10965 );
xor ( n10967 , n10939 , n10966 );
xor ( n10968 , n10936 , n10967 );
buf ( n10969 , n5708 );
not ( n10970 , n6474 );
buf ( n10971 , n5709 );
and ( n10972 , n10970 , n10971 );
buf ( n10973 , n5710 );
xor ( n10974 , n10973 , n10971 );
and ( n10975 , n10974 , n6474 );
or ( n10976 , n10972 , n10975 );
not ( n10977 , n6474 );
buf ( n10978 , n5711 );
and ( n10979 , n10977 , n10978 );
buf ( n10980 , n5712 );
xor ( n10981 , n10980 , n10978 );
and ( n10982 , n10981 , n6474 );
or ( n10983 , n10979 , n10982 );
xor ( n10984 , n10976 , n10983 );
buf ( n10985 , n5713 );
xor ( n10986 , n10984 , n10985 );
buf ( n10987 , n5714 );
xor ( n10988 , n10986 , n10987 );
buf ( n10989 , n5715 );
xor ( n10990 , n10988 , n10989 );
xor ( n10991 , n10969 , n10990 );
xor ( n10992 , n10991 , n10022 );
xor ( n10993 , n7830 , n7399 );
xor ( n10994 , n10993 , n7421 );
not ( n10995 , n10994 );
not ( n10996 , n6474 );
buf ( n10997 , n5716 );
and ( n10998 , n10996 , n10997 );
buf ( n10999 , n5717 );
xor ( n11000 , n10999 , n10997 );
and ( n11001 , n11000 , n6474 );
or ( n11002 , n10998 , n11001 );
xor ( n11003 , n11002 , n7376 );
xor ( n11004 , n11003 , n10465 );
and ( n11005 , n10995 , n11004 );
xor ( n11006 , n10992 , n11005 );
xor ( n11007 , n10968 , n11006 );
buf ( n11008 , n5718 );
xor ( n11009 , n11008 , n9047 );
xor ( n11010 , n11009 , n9338 );
not ( n11011 , n6474 );
buf ( n11012 , n5719 );
and ( n11013 , n11011 , n11012 );
buf ( n11014 , n5720 );
xor ( n11015 , n11014 , n11012 );
and ( n11016 , n11015 , n6474 );
or ( n11017 , n11013 , n11016 );
not ( n11018 , n6474 );
buf ( n11019 , n5721 );
and ( n11020 , n11018 , n11019 );
buf ( n11021 , n5722 );
xor ( n11022 , n11021 , n11019 );
and ( n11023 , n11022 , n6474 );
or ( n11024 , n11020 , n11023 );
xor ( n11025 , n11017 , n11024 );
buf ( n11026 , n5723 );
xor ( n11027 , n11025 , n11026 );
buf ( n11028 , n5724 );
xor ( n11029 , n11027 , n11028 );
buf ( n11030 , n5725 );
xor ( n11031 , n11029 , n11030 );
xor ( n11032 , n7016 , n11031 );
not ( n11033 , n6474 );
buf ( n11034 , n5726 );
and ( n11035 , n11033 , n11034 );
buf ( n11036 , n5727 );
xor ( n11037 , n11036 , n11034 );
and ( n11038 , n11037 , n6474 );
or ( n11039 , n11035 , n11038 );
not ( n11040 , n6474 );
buf ( n11041 , n5728 );
and ( n11042 , n11040 , n11041 );
buf ( n11043 , n5729 );
xor ( n11044 , n11043 , n11041 );
and ( n11045 , n11044 , n6474 );
or ( n11046 , n11042 , n11045 );
xor ( n11047 , n11039 , n11046 );
buf ( n11048 , n5730 );
xor ( n11049 , n11047 , n11048 );
buf ( n11050 , n5731 );
xor ( n11051 , n11049 , n11050 );
xor ( n11052 , n11051 , n7500 );
xor ( n11053 , n11032 , n11052 );
not ( n11054 , n11053 );
not ( n11055 , n6474 );
buf ( n11056 , n5732 );
and ( n11057 , n11055 , n11056 );
buf ( n11058 , n5733 );
xor ( n11059 , n11058 , n11056 );
and ( n11060 , n11059 , n6474 );
or ( n11061 , n11057 , n11060 );
xor ( n11062 , n11061 , n10697 );
xor ( n11063 , n11062 , n10713 );
and ( n11064 , n11054 , n11063 );
xor ( n11065 , n11010 , n11064 );
xor ( n11066 , n11007 , n11065 );
xor ( n11067 , n10888 , n11066 );
not ( n11068 , n11067 );
not ( n11069 , n6474 );
buf ( n11070 , n5734 );
and ( n11071 , n11069 , n11070 );
buf ( n11072 , n5735 );
xor ( n11073 , n11072 , n11070 );
and ( n11074 , n11073 , n6474 );
or ( n11075 , n11071 , n11074 );
not ( n11076 , n6474 );
buf ( n11077 , n5736 );
and ( n11078 , n11076 , n11077 );
buf ( n11079 , n5737 );
xor ( n11080 , n11079 , n11077 );
and ( n11081 , n11080 , n6474 );
or ( n11082 , n11078 , n11081 );
xor ( n11083 , n11075 , n11082 );
buf ( n11084 , n5738 );
xor ( n11085 , n11083 , n11084 );
buf ( n11086 , n5739 );
xor ( n11087 , n11085 , n11086 );
buf ( n11088 , n5740 );
xor ( n11089 , n11087 , n11088 );
xor ( n11090 , n10043 , n11089 );
not ( n11091 , n6474 );
buf ( n11092 , n5741 );
and ( n11093 , n11091 , n11092 );
buf ( n11094 , n5742 );
xor ( n11095 , n11094 , n11092 );
and ( n11096 , n11095 , n6474 );
or ( n11097 , n11093 , n11096 );
not ( n11098 , n6474 );
buf ( n11099 , n5743 );
and ( n11100 , n11098 , n11099 );
buf ( n11101 , n5744 );
xor ( n11102 , n11101 , n11099 );
and ( n11103 , n11102 , n6474 );
or ( n11104 , n11100 , n11103 );
xor ( n11105 , n11097 , n11104 );
buf ( n11106 , n5745 );
xor ( n11107 , n11105 , n11106 );
buf ( n11108 , n5746 );
xor ( n11109 , n11107 , n11108 );
xor ( n11110 , n11109 , n7748 );
xor ( n11111 , n11090 , n11110 );
not ( n11112 , n6474 );
buf ( n11113 , n5747 );
and ( n11114 , n11112 , n11113 );
buf ( n11115 , n5748 );
xor ( n11116 , n11115 , n11113 );
and ( n11117 , n11116 , n6474 );
or ( n11118 , n11114 , n11117 );
not ( n11119 , n6474 );
buf ( n11120 , n5749 );
and ( n11121 , n11119 , n11120 );
buf ( n11122 , n5750 );
xor ( n11123 , n11122 , n11120 );
and ( n11124 , n11123 , n6474 );
or ( n11125 , n11121 , n11124 );
xor ( n11126 , n11118 , n11125 );
buf ( n11127 , n5751 );
xor ( n11128 , n11126 , n11127 );
buf ( n11129 , n5752 );
xor ( n11130 , n11128 , n11129 );
buf ( n11131 , n5753 );
xor ( n11132 , n11130 , n11131 );
xor ( n11133 , n8174 , n11132 );
not ( n11134 , n6474 );
buf ( n11135 , n5754 );
and ( n11136 , n11134 , n11135 );
buf ( n11137 , n5755 );
xor ( n11138 , n11137 , n11135 );
and ( n11139 , n11138 , n6474 );
or ( n11140 , n11136 , n11139 );
xor ( n11141 , n11140 , n11061 );
buf ( n11142 , n5756 );
xor ( n11143 , n11141 , n11142 );
buf ( n11144 , n5757 );
xor ( n11145 , n11143 , n11144 );
xor ( n11146 , n11145 , n10676 );
xor ( n11147 , n11133 , n11146 );
not ( n11148 , n11147 );
not ( n11149 , n6474 );
buf ( n11150 , n5758 );
and ( n11151 , n11149 , n11150 );
buf ( n11152 , n5759 );
xor ( n11153 , n11152 , n11150 );
and ( n11154 , n11153 , n6474 );
or ( n11155 , n11151 , n11154 );
xor ( n11156 , n11155 , n8799 );
not ( n11157 , n6474 );
buf ( n11158 , n5760 );
and ( n11159 , n11157 , n11158 );
buf ( n11160 , n5761 );
xor ( n11161 , n11160 , n11158 );
and ( n11162 , n11161 , n6474 );
or ( n11163 , n11159 , n11162 );
buf ( n11164 , n5762 );
xor ( n11165 , n11163 , n11164 );
buf ( n11166 , n5763 );
xor ( n11167 , n11165 , n11166 );
buf ( n11168 , n5764 );
xor ( n11169 , n11167 , n11168 );
buf ( n11170 , n5765 );
xor ( n11171 , n11169 , n11170 );
xor ( n11172 , n11156 , n11171 );
and ( n11173 , n11148 , n11172 );
xor ( n11174 , n11111 , n11173 );
not ( n11175 , n6474 );
buf ( n11176 , n5766 );
and ( n11177 , n11175 , n11176 );
buf ( n11178 , n5767 );
xor ( n11179 , n11178 , n11176 );
and ( n11180 , n11179 , n6474 );
or ( n11181 , n11177 , n11180 );
xor ( n11182 , n11181 , n7474 );
buf ( n11183 , n5768 );
xor ( n11184 , n11182 , n11183 );
xor ( n11185 , n11184 , n8164 );
buf ( n11186 , n5769 );
xor ( n11187 , n11185 , n11186 );
xor ( n11188 , n10765 , n11187 );
not ( n11189 , n6474 );
buf ( n11190 , n5770 );
and ( n11191 , n11189 , n11190 );
buf ( n11192 , n5771 );
xor ( n11193 , n11192 , n11190 );
and ( n11194 , n11193 , n6474 );
or ( n11195 , n11191 , n11194 );
buf ( n11196 , n5772 );
xor ( n11197 , n11195 , n11196 );
buf ( n11198 , n5773 );
xor ( n11199 , n11197 , n11198 );
xor ( n11200 , n11199 , n6829 );
xor ( n11201 , n11200 , n10889 );
xor ( n11202 , n11188 , n11201 );
xor ( n11203 , n6583 , n7732 );
xor ( n11204 , n11203 , n8076 );
not ( n11205 , n11204 );
xor ( n11206 , n9637 , n10713 );
not ( n11207 , n6474 );
buf ( n11208 , n5774 );
and ( n11209 , n11207 , n11208 );
buf ( n11210 , n5775 );
xor ( n11211 , n11210 , n11208 );
and ( n11212 , n11211 , n6474 );
or ( n11213 , n11209 , n11212 );
not ( n11214 , n6474 );
buf ( n11215 , n5776 );
and ( n11216 , n11214 , n11215 );
buf ( n11217 , n5777 );
xor ( n11218 , n11217 , n11215 );
and ( n11219 , n11218 , n6474 );
or ( n11220 , n11216 , n11219 );
xor ( n11221 , n11213 , n11220 );
buf ( n11222 , n5778 );
xor ( n11223 , n11221 , n11222 );
buf ( n11224 , n5779 );
xor ( n11225 , n11223 , n11224 );
buf ( n11226 , n5780 );
xor ( n11227 , n11225 , n11226 );
xor ( n11228 , n11206 , n11227 );
and ( n11229 , n11205 , n11228 );
xor ( n11230 , n11202 , n11229 );
xor ( n11231 , n10462 , n10246 );
not ( n11232 , n6474 );
buf ( n11233 , n5781 );
and ( n11234 , n11232 , n11233 );
buf ( n11235 , n5782 );
xor ( n11236 , n11235 , n11233 );
and ( n11237 , n11236 , n6474 );
or ( n11238 , n11234 , n11237 );
not ( n11239 , n6474 );
buf ( n11240 , n5783 );
and ( n11241 , n11239 , n11240 );
buf ( n11242 , n5784 );
xor ( n11243 , n11242 , n11240 );
and ( n11244 , n11243 , n6474 );
or ( n11245 , n11241 , n11244 );
xor ( n11246 , n11238 , n11245 );
buf ( n11247 , n5785 );
xor ( n11248 , n11246 , n11247 );
buf ( n11249 , n5786 );
xor ( n11250 , n11248 , n11249 );
buf ( n11251 , n5787 );
xor ( n11252 , n11250 , n11251 );
xor ( n11253 , n11231 , n11252 );
buf ( n11254 , n5788 );
not ( n11255 , n6474 );
buf ( n11256 , n5789 );
and ( n11257 , n11255 , n11256 );
buf ( n11258 , n5790 );
xor ( n11259 , n11258 , n11256 );
and ( n11260 , n11259 , n6474 );
or ( n11261 , n11257 , n11260 );
not ( n11262 , n6474 );
buf ( n11263 , n5791 );
and ( n11264 , n11262 , n11263 );
buf ( n11265 , n5792 );
xor ( n11266 , n11265 , n11263 );
and ( n11267 , n11266 , n6474 );
or ( n11268 , n11264 , n11267 );
xor ( n11269 , n11261 , n11268 );
buf ( n11270 , n5793 );
xor ( n11271 , n11269 , n11270 );
buf ( n11272 , n5794 );
xor ( n11273 , n11271 , n11272 );
buf ( n11274 , n5795 );
xor ( n11275 , n11273 , n11274 );
xor ( n11276 , n11254 , n11275 );
xor ( n11277 , n11276 , n9559 );
not ( n11278 , n11277 );
xor ( n11279 , n6524 , n10731 );
xor ( n11280 , n11279 , n10745 );
and ( n11281 , n11278 , n11280 );
xor ( n11282 , n11253 , n11281 );
xor ( n11283 , n11230 , n11282 );
not ( n11284 , n6474 );
buf ( n11285 , n5796 );
and ( n11286 , n11284 , n11285 );
buf ( n11287 , n5797 );
xor ( n11288 , n11287 , n11285 );
and ( n11289 , n11288 , n6474 );
or ( n11290 , n11286 , n11289 );
not ( n11291 , n6474 );
buf ( n11292 , n5798 );
and ( n11293 , n11291 , n11292 );
buf ( n11294 , n5799 );
xor ( n11295 , n11294 , n11292 );
and ( n11296 , n11295 , n6474 );
or ( n11297 , n11293 , n11296 );
xor ( n11298 , n11290 , n11297 );
buf ( n11299 , n5800 );
xor ( n11300 , n11298 , n11299 );
buf ( n11301 , n5801 );
xor ( n11302 , n11300 , n11301 );
buf ( n11303 , n5802 );
xor ( n11304 , n11302 , n11303 );
xor ( n11305 , n7534 , n11304 );
xor ( n11306 , n11305 , n9850 );
buf ( n11307 , n5803 );
xor ( n11308 , n11307 , n9002 );
not ( n11309 , n6474 );
buf ( n11310 , n5804 );
and ( n11311 , n11309 , n11310 );
buf ( n11312 , n5805 );
xor ( n11313 , n11312 , n11310 );
and ( n11314 , n11313 , n6474 );
or ( n11315 , n11311 , n11314 );
not ( n11316 , n6474 );
buf ( n11317 , n5806 );
and ( n11318 , n11316 , n11317 );
buf ( n11319 , n5807 );
xor ( n11320 , n11319 , n11317 );
and ( n11321 , n11320 , n6474 );
or ( n11322 , n11318 , n11321 );
xor ( n11323 , n11315 , n11322 );
buf ( n11324 , n5808 );
xor ( n11325 , n11323 , n11324 );
buf ( n11326 , n5809 );
xor ( n11327 , n11325 , n11326 );
buf ( n11328 , n5810 );
xor ( n11329 , n11327 , n11328 );
xor ( n11330 , n11308 , n11329 );
not ( n11331 , n11330 );
not ( n11332 , n6474 );
buf ( n11333 , n5811 );
and ( n11334 , n11332 , n11333 );
buf ( n11335 , n5812 );
xor ( n11336 , n11335 , n11333 );
and ( n11337 , n11336 , n6474 );
or ( n11338 , n11334 , n11337 );
xor ( n11339 , n11338 , n10007 );
buf ( n11340 , n5813 );
xor ( n11341 , n11339 , n11340 );
buf ( n11342 , n5814 );
xor ( n11343 , n11341 , n11342 );
buf ( n11344 , n5815 );
xor ( n11345 , n11343 , n11344 );
xor ( n11346 , n11213 , n11345 );
not ( n11347 , n6474 );
buf ( n11348 , n5816 );
and ( n11349 , n11347 , n11348 );
buf ( n11350 , n5817 );
xor ( n11351 , n11350 , n11348 );
and ( n11352 , n11351 , n6474 );
or ( n11353 , n11349 , n11352 );
not ( n11354 , n6474 );
buf ( n11355 , n5818 );
and ( n11356 , n11354 , n11355 );
buf ( n11357 , n5819 );
xor ( n11358 , n11357 , n11355 );
and ( n11359 , n11358 , n6474 );
or ( n11360 , n11356 , n11359 );
xor ( n11361 , n11353 , n11360 );
buf ( n11362 , n5820 );
xor ( n11363 , n11361 , n11362 );
buf ( n11364 , n5821 );
xor ( n11365 , n11363 , n11364 );
buf ( n11366 , n5822 );
xor ( n11367 , n11365 , n11366 );
xor ( n11368 , n11346 , n11367 );
and ( n11369 , n11331 , n11368 );
xor ( n11370 , n11306 , n11369 );
xor ( n11371 , n11283 , n11370 );
xor ( n11372 , n9531 , n6606 );
xor ( n11373 , n11372 , n9123 );
buf ( n11374 , n5823 );
xor ( n11375 , n11374 , n9217 );
xor ( n11376 , n11375 , n9417 );
not ( n11377 , n11376 );
not ( n11378 , n6474 );
buf ( n11379 , n5824 );
and ( n11380 , n11378 , n11379 );
buf ( n11381 , n5825 );
xor ( n11382 , n11381 , n11379 );
and ( n11383 , n11382 , n6474 );
or ( n11384 , n11380 , n11383 );
xor ( n11385 , n11384 , n8495 );
xor ( n11386 , n11385 , n8517 );
and ( n11387 , n11377 , n11386 );
xor ( n11388 , n11373 , n11387 );
xor ( n11389 , n11371 , n11388 );
buf ( n11390 , n5826 );
not ( n11391 , n6474 );
buf ( n11392 , n5827 );
and ( n11393 , n11391 , n11392 );
buf ( n11394 , n5828 );
xor ( n11395 , n11394 , n11392 );
and ( n11396 , n11395 , n6474 );
or ( n11397 , n11393 , n11396 );
buf ( n11398 , n5829 );
xor ( n11399 , n11397 , n11398 );
buf ( n11400 , n5830 );
xor ( n11401 , n11399 , n11400 );
buf ( n11402 , n5831 );
xor ( n11403 , n11401 , n11402 );
buf ( n11404 , n5832 );
xor ( n11405 , n11403 , n11404 );
xor ( n11406 , n11390 , n11405 );
not ( n11407 , n6474 );
buf ( n11408 , n5833 );
and ( n11409 , n11407 , n11408 );
buf ( n11410 , n5834 );
xor ( n11411 , n11410 , n11408 );
and ( n11412 , n11411 , n6474 );
or ( n11413 , n11409 , n11412 );
not ( n11414 , n6474 );
buf ( n11415 , n5835 );
and ( n11416 , n11414 , n11415 );
buf ( n11417 , n5836 );
xor ( n11418 , n11417 , n11415 );
and ( n11419 , n11418 , n6474 );
or ( n11420 , n11416 , n11419 );
xor ( n11421 , n11413 , n11420 );
buf ( n11422 , n5837 );
xor ( n11423 , n11421 , n11422 );
buf ( n11424 , n5838 );
xor ( n11425 , n11423 , n11424 );
buf ( n11426 , n5839 );
xor ( n11427 , n11425 , n11426 );
xor ( n11428 , n11406 , n11427 );
not ( n11429 , n11111 );
and ( n11430 , n11429 , n11147 );
xor ( n11431 , n11428 , n11430 );
xor ( n11432 , n11389 , n11431 );
xor ( n11433 , n11174 , n11432 );
xor ( n11434 , n11338 , n10022 );
xor ( n11435 , n11434 , n10044 );
xor ( n11436 , n10458 , n10246 );
xor ( n11437 , n11436 , n11252 );
not ( n11438 , n11437 );
xor ( n11439 , n9285 , n8660 );
xor ( n11440 , n11439 , n10105 );
and ( n11441 , n11438 , n11440 );
xor ( n11442 , n11435 , n11441 );
not ( n11443 , n6474 );
buf ( n11444 , n5840 );
and ( n11445 , n11443 , n11444 );
buf ( n11446 , n5841 );
xor ( n11447 , n11446 , n11444 );
and ( n11448 , n11447 , n6474 );
or ( n11449 , n11445 , n11448 );
not ( n11450 , n6474 );
buf ( n11451 , n5842 );
and ( n11452 , n11450 , n11451 );
buf ( n11453 , n5843 );
xor ( n11454 , n11453 , n11451 );
and ( n11455 , n11454 , n6474 );
or ( n11456 , n11452 , n11455 );
xor ( n11457 , n11449 , n11456 );
buf ( n11458 , n5844 );
xor ( n11459 , n11457 , n11458 );
xor ( n11460 , n11459 , n6963 );
buf ( n11461 , n5845 );
xor ( n11462 , n11460 , n11461 );
xor ( n11463 , n7194 , n11462 );
xor ( n11464 , n11463 , n10263 );
xor ( n11465 , n10139 , n10768 );
xor ( n11466 , n11465 , n10790 );
not ( n11467 , n11466 );
not ( n11468 , n6474 );
buf ( n11469 , n5846 );
and ( n11470 , n11468 , n11469 );
buf ( n11471 , n5847 );
xor ( n11472 , n11471 , n11469 );
and ( n11473 , n11472 , n6474 );
or ( n11474 , n11470 , n11473 );
buf ( n11475 , n5848 );
xor ( n11476 , n11474 , n11475 );
xor ( n11477 , n11476 , n10148 );
buf ( n11478 , n5849 );
xor ( n11479 , n11477 , n11478 );
buf ( n11480 , n5850 );
xor ( n11481 , n11479 , n11480 );
xor ( n11482 , n8908 , n11481 );
xor ( n11483 , n11482 , n8696 );
and ( n11484 , n11467 , n11483 );
xor ( n11485 , n11464 , n11484 );
xor ( n11486 , n11442 , n11485 );
xor ( n11487 , n10030 , n11089 );
xor ( n11488 , n11487 , n11110 );
xor ( n11489 , n7514 , n8016 );
xor ( n11490 , n11489 , n11304 );
not ( n11491 , n11490 );
not ( n11492 , n6474 );
buf ( n11493 , n5851 );
and ( n11494 , n11492 , n11493 );
buf ( n11495 , n5852 );
xor ( n11496 , n11495 , n11493 );
and ( n11497 , n11496 , n6474 );
or ( n11498 , n11494 , n11497 );
not ( n11499 , n6474 );
buf ( n11500 , n5853 );
and ( n11501 , n11499 , n11500 );
buf ( n11502 , n5854 );
xor ( n11503 , n11502 , n11500 );
and ( n11504 , n11503 , n6474 );
or ( n11505 , n11501 , n11504 );
xor ( n11506 , n11498 , n11505 );
buf ( n11507 , n5855 );
xor ( n11508 , n11506 , n11507 );
buf ( n11509 , n5856 );
xor ( n11510 , n11508 , n11509 );
buf ( n11511 , n5857 );
xor ( n11512 , n11510 , n11511 );
xor ( n11513 , n7856 , n11512 );
xor ( n11514 , n11384 , n8475 );
buf ( n11515 , n5858 );
xor ( n11516 , n11514 , n11515 );
buf ( n11517 , n5859 );
xor ( n11518 , n11516 , n11517 );
buf ( n11519 , n5860 );
xor ( n11520 , n11518 , n11519 );
xor ( n11521 , n11513 , n11520 );
and ( n11522 , n11491 , n11521 );
xor ( n11523 , n11488 , n11522 );
xor ( n11524 , n11486 , n11523 );
xor ( n11525 , n7918 , n6538 );
xor ( n11526 , n11525 , n6560 );
not ( n11527 , n6474 );
buf ( n11528 , n5861 );
and ( n11529 , n11527 , n11528 );
buf ( n11530 , n5862 );
xor ( n11531 , n11530 , n11528 );
and ( n11532 , n11531 , n6474 );
or ( n11533 , n11529 , n11532 );
xor ( n11534 , n11533 , n10929 );
not ( n11535 , n6474 );
buf ( n11536 , n5863 );
and ( n11537 , n11535 , n11536 );
buf ( n11538 , n5864 );
xor ( n11539 , n11538 , n11536 );
and ( n11540 , n11539 , n6474 );
or ( n11541 , n11537 , n11540 );
not ( n11542 , n6474 );
buf ( n11543 , n5865 );
and ( n11544 , n11542 , n11543 );
buf ( n11545 , n5866 );
xor ( n11546 , n11545 , n11543 );
and ( n11547 , n11546 , n6474 );
or ( n11548 , n11544 , n11547 );
xor ( n11549 , n11541 , n11548 );
buf ( n11550 , n5867 );
xor ( n11551 , n11549 , n11550 );
buf ( n11552 , n5868 );
xor ( n11553 , n11551 , n11552 );
buf ( n11554 , n5869 );
xor ( n11555 , n11553 , n11554 );
xor ( n11556 , n11534 , n11555 );
not ( n11557 , n11556 );
xor ( n11558 , n6758 , n9400 );
xor ( n11559 , n11558 , n10309 );
and ( n11560 , n11557 , n11559 );
xor ( n11561 , n11526 , n11560 );
xor ( n11562 , n11524 , n11561 );
not ( n11563 , n6474 );
buf ( n11564 , n5870 );
and ( n11565 , n11563 , n11564 );
buf ( n11566 , n5871 );
xor ( n11567 , n11566 , n11564 );
and ( n11568 , n11567 , n6474 );
or ( n11569 , n11565 , n11568 );
not ( n11570 , n6474 );
buf ( n11571 , n5872 );
and ( n11572 , n11570 , n11571 );
buf ( n11573 , n5873 );
xor ( n11574 , n11573 , n11571 );
and ( n11575 , n11574 , n6474 );
or ( n11576 , n11572 , n11575 );
xor ( n11577 , n11569 , n11576 );
buf ( n11578 , n5874 );
xor ( n11579 , n11577 , n11578 );
buf ( n11580 , n5875 );
xor ( n11581 , n11579 , n11580 );
buf ( n11582 , n5876 );
xor ( n11583 , n11581 , n11582 );
xor ( n11584 , n10683 , n11583 );
not ( n11585 , n6474 );
buf ( n11586 , n5877 );
and ( n11587 , n11585 , n11586 );
buf ( n11588 , n5878 );
xor ( n11589 , n11588 , n11586 );
and ( n11590 , n11589 , n6474 );
or ( n11591 , n11587 , n11590 );
not ( n11592 , n6474 );
buf ( n11593 , n5879 );
and ( n11594 , n11592 , n11593 );
buf ( n11595 , n5880 );
xor ( n11596 , n11595 , n11593 );
and ( n11597 , n11596 , n6474 );
or ( n11598 , n11594 , n11597 );
xor ( n11599 , n11591 , n11598 );
buf ( n11600 , n5881 );
xor ( n11601 , n11599 , n11600 );
buf ( n11602 , n5882 );
xor ( n11603 , n11601 , n11602 );
xor ( n11604 , n11603 , n10969 );
xor ( n11605 , n11584 , n11604 );
not ( n11606 , n6474 );
buf ( n11607 , n5883 );
and ( n11608 , n11606 , n11607 );
buf ( n11609 , n5884 );
xor ( n11610 , n11609 , n11607 );
and ( n11611 , n11610 , n6474 );
or ( n11612 , n11608 , n11611 );
xor ( n11613 , n11612 , n9217 );
xor ( n11614 , n11613 , n9417 );
not ( n11615 , n11614 );
not ( n11616 , n6474 );
buf ( n11617 , n5885 );
and ( n11618 , n11616 , n11617 );
buf ( n11619 , n5886 );
xor ( n11620 , n11619 , n11617 );
and ( n11621 , n11620 , n6474 );
or ( n11622 , n11618 , n11621 );
not ( n11623 , n6474 );
buf ( n11624 , n5887 );
and ( n11625 , n11623 , n11624 );
buf ( n11626 , n5888 );
xor ( n11627 , n11626 , n11624 );
and ( n11628 , n11627 , n6474 );
or ( n11629 , n11625 , n11628 );
xor ( n11630 , n11622 , n11629 );
buf ( n11631 , n5889 );
xor ( n11632 , n11630 , n11631 );
buf ( n11633 , n5890 );
xor ( n11634 , n11632 , n11633 );
buf ( n11635 , n5891 );
xor ( n11636 , n11634 , n11635 );
xor ( n11637 , n6822 , n11636 );
not ( n11638 , n6474 );
buf ( n11639 , n5892 );
and ( n11640 , n11638 , n11639 );
buf ( n11641 , n5893 );
xor ( n11642 , n11641 , n11639 );
and ( n11643 , n11642 , n6474 );
or ( n11644 , n11640 , n11643 );
not ( n11645 , n6474 );
buf ( n11646 , n5894 );
and ( n11647 , n11645 , n11646 );
buf ( n11648 , n5895 );
xor ( n11649 , n11648 , n11646 );
and ( n11650 , n11649 , n6474 );
or ( n11651 , n11647 , n11650 );
xor ( n11652 , n11644 , n11651 );
buf ( n11653 , n5896 );
xor ( n11654 , n11652 , n11653 );
xor ( n11655 , n11654 , n11390 );
buf ( n11656 , n5897 );
xor ( n11657 , n11655 , n11656 );
xor ( n11658 , n11637 , n11657 );
and ( n11659 , n11615 , n11658 );
xor ( n11660 , n11605 , n11659 );
xor ( n11661 , n11562 , n11660 );
xor ( n11662 , n11433 , n11661 );
and ( n11663 , n11068 , n11662 );
xor ( n11664 , n10631 , n11663 );
and ( n11665 , n11664 , n6475 );
or ( n11666 , n9748 , n11665 );
and ( n11667 , n9745 , n11666 );
buf ( n11668 , n11667 );
buf ( n11669 , n11668 );
not ( n11670 , n6469 );
not ( n11671 , n6475 );
and ( n11672 , n11671 , n9661 );
xor ( n11673 , n8682 , n10170 );
xor ( n11674 , n11673 , n7030 );
not ( n11675 , n6474 );
buf ( n11676 , n5898 );
and ( n11677 , n11675 , n11676 );
buf ( n11678 , n5899 );
xor ( n11679 , n11678 , n11676 );
and ( n11680 , n11679 , n6474 );
or ( n11681 , n11677 , n11680 );
not ( n11682 , n6474 );
buf ( n11683 , n5900 );
and ( n11684 , n11682 , n11683 );
buf ( n11685 , n5901 );
xor ( n11686 , n11685 , n11683 );
and ( n11687 , n11686 , n6474 );
or ( n11688 , n11684 , n11687 );
xor ( n11689 , n11681 , n11688 );
buf ( n11690 , n5902 );
xor ( n11691 , n11689 , n11690 );
xor ( n11692 , n11691 , n9948 );
xor ( n11693 , n11692 , n11008 );
xor ( n11694 , n9865 , n11693 );
not ( n11695 , n6474 );
buf ( n11696 , n5903 );
and ( n11697 , n11695 , n11696 );
buf ( n11698 , n5904 );
xor ( n11699 , n11698 , n11696 );
and ( n11700 , n11699 , n6474 );
or ( n11701 , n11697 , n11700 );
not ( n11702 , n6474 );
buf ( n11703 , n5905 );
and ( n11704 , n11702 , n11703 );
buf ( n11705 , n5906 );
xor ( n11706 , n11705 , n11703 );
and ( n11707 , n11706 , n6474 );
or ( n11708 , n11704 , n11707 );
xor ( n11709 , n11701 , n11708 );
buf ( n11710 , n5907 );
xor ( n11711 , n11709 , n11710 );
xor ( n11712 , n11711 , n9318 );
buf ( n11713 , n5908 );
xor ( n11714 , n11712 , n11713 );
xor ( n11715 , n11694 , n11714 );
not ( n11716 , n11715 );
xor ( n11717 , n7203 , n11462 );
xor ( n11718 , n11717 , n10263 );
and ( n11719 , n11716 , n11718 );
xor ( n11720 , n11674 , n11719 );
not ( n11721 , n6474 );
buf ( n11722 , n5909 );
and ( n11723 , n11721 , n11722 );
buf ( n11724 , n5910 );
xor ( n11725 , n11724 , n11722 );
and ( n11726 , n11725 , n6474 );
or ( n11727 , n11723 , n11726 );
not ( n11728 , n6474 );
buf ( n11729 , n5911 );
and ( n11730 , n11728 , n11729 );
buf ( n11731 , n5912 );
xor ( n11732 , n11731 , n11729 );
and ( n11733 , n11732 , n6474 );
or ( n11734 , n11730 , n11733 );
xor ( n11735 , n11727 , n11734 );
buf ( n11736 , n5913 );
xor ( n11737 , n11735 , n11736 );
buf ( n11738 , n5914 );
xor ( n11739 , n11737 , n11738 );
buf ( n11740 , n5915 );
xor ( n11741 , n11739 , n11740 );
xor ( n11742 , n9001 , n11741 );
not ( n11743 , n6474 );
buf ( n11744 , n5916 );
and ( n11745 , n11743 , n11744 );
buf ( n11746 , n5917 );
xor ( n11747 , n11746 , n11744 );
and ( n11748 , n11747 , n6474 );
or ( n11749 , n11745 , n11748 );
not ( n11750 , n6474 );
buf ( n11751 , n5918 );
and ( n11752 , n11750 , n11751 );
buf ( n11753 , n5919 );
xor ( n11754 , n11753 , n11751 );
and ( n11755 , n11754 , n6474 );
or ( n11756 , n11752 , n11755 );
xor ( n11757 , n11749 , n11756 );
buf ( n11758 , n5920 );
xor ( n11759 , n11757 , n11758 );
buf ( n11760 , n5921 );
xor ( n11761 , n11759 , n11760 );
buf ( n11762 , n5922 );
xor ( n11763 , n11761 , n11762 );
xor ( n11764 , n11742 , n11763 );
xor ( n11765 , n8899 , n11481 );
xor ( n11766 , n11765 , n8696 );
not ( n11767 , n11766 );
not ( n11768 , n6474 );
buf ( n11769 , n5923 );
and ( n11770 , n11768 , n11769 );
buf ( n11771 , n5924 );
xor ( n11772 , n11771 , n11769 );
and ( n11773 , n11772 , n6474 );
or ( n11774 , n11770 , n11773 );
not ( n11775 , n6474 );
buf ( n11776 , n5925 );
and ( n11777 , n11775 , n11776 );
buf ( n11778 , n5926 );
xor ( n11779 , n11778 , n11776 );
and ( n11780 , n11779 , n6474 );
or ( n11781 , n11777 , n11780 );
xor ( n11782 , n11774 , n11781 );
buf ( n11783 , n5927 );
xor ( n11784 , n11782 , n11783 );
xor ( n11785 , n11784 , n10878 );
xor ( n11786 , n11785 , n10379 );
xor ( n11787 , n8284 , n11786 );
not ( n11788 , n6474 );
buf ( n11789 , n5928 );
and ( n11790 , n11788 , n11789 );
buf ( n11791 , n5929 );
xor ( n11792 , n11791 , n11789 );
and ( n11793 , n11792 , n6474 );
or ( n11794 , n11790 , n11793 );
not ( n11795 , n6474 );
buf ( n11796 , n5930 );
and ( n11797 , n11795 , n11796 );
buf ( n11798 , n5931 );
xor ( n11799 , n11798 , n11796 );
and ( n11800 , n11799 , n6474 );
or ( n11801 , n11797 , n11800 );
xor ( n11802 , n11794 , n11801 );
buf ( n11803 , n5932 );
xor ( n11804 , n11802 , n11803 );
buf ( n11805 , n5933 );
xor ( n11806 , n11804 , n11805 );
buf ( n11807 , n5934 );
xor ( n11808 , n11806 , n11807 );
xor ( n11809 , n11787 , n11808 );
and ( n11810 , n11767 , n11809 );
xor ( n11811 , n11764 , n11810 );
xor ( n11812 , n9672 , n11227 );
not ( n11813 , n6474 );
buf ( n11814 , n5935 );
and ( n11815 , n11813 , n11814 );
buf ( n11816 , n5936 );
xor ( n11817 , n11816 , n11814 );
and ( n11818 , n11817 , n6474 );
or ( n11819 , n11815 , n11818 );
not ( n11820 , n6474 );
buf ( n11821 , n5937 );
and ( n11822 , n11820 , n11821 );
buf ( n11823 , n5938 );
xor ( n11824 , n11823 , n11821 );
and ( n11825 , n11824 , n6474 );
or ( n11826 , n11822 , n11825 );
xor ( n11827 , n11819 , n11826 );
buf ( n11828 , n5939 );
xor ( n11829 , n11827 , n11828 );
buf ( n11830 , n5940 );
xor ( n11831 , n11829 , n11830 );
buf ( n11832 , n5941 );
xor ( n11833 , n11831 , n11832 );
xor ( n11834 , n11812 , n11833 );
not ( n11835 , n6474 );
buf ( n11836 , n5942 );
and ( n11837 , n11835 , n11836 );
buf ( n11838 , n5943 );
xor ( n11839 , n11838 , n11836 );
and ( n11840 , n11839 , n6474 );
or ( n11841 , n11837 , n11840 );
xor ( n11842 , n11841 , n8574 );
xor ( n11843 , n11842 , n7441 );
not ( n11844 , n11843 );
not ( n11845 , n6474 );
buf ( n11846 , n5944 );
and ( n11847 , n11845 , n11846 );
buf ( n11848 , n5945 );
xor ( n11849 , n11848 , n11846 );
and ( n11850 , n11849 , n6474 );
or ( n11851 , n11847 , n11850 );
not ( n11852 , n6474 );
buf ( n11853 , n5946 );
and ( n11854 , n11852 , n11853 );
buf ( n11855 , n5947 );
xor ( n11856 , n11855 , n11853 );
and ( n11857 , n11856 , n6474 );
or ( n11858 , n11854 , n11857 );
xor ( n11859 , n11851 , n11858 );
buf ( n11860 , n5948 );
xor ( n11861 , n11859 , n11860 );
buf ( n11862 , n5949 );
xor ( n11863 , n11861 , n11862 );
buf ( n11864 , n5950 );
xor ( n11865 , n11863 , n11864 );
xor ( n11866 , n8085 , n11865 );
not ( n11867 , n6474 );
buf ( n11868 , n5951 );
and ( n11869 , n11867 , n11868 );
buf ( n11870 , n5952 );
xor ( n11871 , n11870 , n11868 );
and ( n11872 , n11871 , n6474 );
or ( n11873 , n11869 , n11872 );
xor ( n11874 , n11873 , n9133 );
buf ( n11875 , n5953 );
xor ( n11876 , n11874 , n11875 );
buf ( n11877 , n5954 );
xor ( n11878 , n11876 , n11877 );
xor ( n11879 , n11878 , n10868 );
xor ( n11880 , n11866 , n11879 );
and ( n11881 , n11844 , n11880 );
xor ( n11882 , n11834 , n11881 );
xor ( n11883 , n11811 , n11882 );
xor ( n11884 , n10789 , n11201 );
not ( n11885 , n6474 );
buf ( n11886 , n5955 );
and ( n11887 , n11885 , n11886 );
buf ( n11888 , n5956 );
xor ( n11889 , n11888 , n11886 );
and ( n11890 , n11889 , n6474 );
or ( n11891 , n11887 , n11890 );
not ( n11892 , n6474 );
buf ( n11893 , n5957 );
and ( n11894 , n11892 , n11893 );
buf ( n11895 , n5958 );
xor ( n11896 , n11895 , n11893 );
and ( n11897 , n11896 , n6474 );
or ( n11898 , n11894 , n11897 );
xor ( n11899 , n11891 , n11898 );
buf ( n11900 , n5959 );
xor ( n11901 , n11899 , n11900 );
buf ( n11902 , n5960 );
xor ( n11903 , n11901 , n11902 );
buf ( n11904 , n5961 );
xor ( n11905 , n11903 , n11904 );
xor ( n11906 , n11884 , n11905 );
not ( n11907 , n11674 );
and ( n11908 , n11907 , n11715 );
xor ( n11909 , n11906 , n11908 );
xor ( n11910 , n11883 , n11909 );
xor ( n11911 , n8841 , n6739 );
not ( n11912 , n6474 );
buf ( n11913 , n5962 );
and ( n11914 , n11912 , n11913 );
buf ( n11915 , n5963 );
xor ( n11916 , n11915 , n11913 );
and ( n11917 , n11916 , n6474 );
or ( n11918 , n11914 , n11917 );
buf ( n11919 , n5964 );
buf ( n11920 , n11919 );
xor ( n11921 , n11918 , n11920 );
buf ( n11922 , n5965 );
xor ( n11923 , n11921 , n11922 );
buf ( n11924 , n5966 );
xor ( n11925 , n11923 , n11924 );
buf ( n11926 , n5967 );
xor ( n11927 , n11925 , n11926 );
xor ( n11928 , n11911 , n11927 );
not ( n11929 , n6474 );
buf ( n11930 , n5968 );
and ( n11931 , n11929 , n11930 );
buf ( n11932 , n5969 );
xor ( n11933 , n11932 , n11930 );
and ( n11934 , n11933 , n6474 );
or ( n11935 , n11931 , n11934 );
not ( n11936 , n6474 );
buf ( n11937 , n5970 );
and ( n11938 , n11936 , n11937 );
buf ( n11939 , n5971 );
xor ( n11940 , n11939 , n11937 );
and ( n11941 , n11940 , n6474 );
or ( n11942 , n11938 , n11941 );
xor ( n11943 , n11935 , n11942 );
buf ( n11944 , n5972 );
xor ( n11945 , n11943 , n11944 );
buf ( n11946 , n5973 );
xor ( n11947 , n11945 , n11946 );
buf ( n11948 , n5974 );
xor ( n11949 , n11947 , n11948 );
xor ( n11950 , n9702 , n11949 );
xor ( n11951 , n11950 , n10574 );
not ( n11952 , n11951 );
not ( n11953 , n6474 );
buf ( n11954 , n5975 );
and ( n11955 , n11953 , n11954 );
buf ( n11956 , n5976 );
xor ( n11957 , n11956 , n11954 );
and ( n11958 , n11957 , n6474 );
or ( n11959 , n11955 , n11958 );
xor ( n11960 , n11959 , n6827 );
not ( n11961 , n6474 );
buf ( n11962 , n5977 );
and ( n11963 , n11961 , n11962 );
buf ( n11964 , n5978 );
xor ( n11965 , n11964 , n11962 );
and ( n11966 , n11965 , n6474 );
or ( n11967 , n11963 , n11966 );
not ( n11968 , n6474 );
buf ( n11969 , n5979 );
and ( n11970 , n11968 , n11969 );
buf ( n11971 , n5980 );
xor ( n11972 , n11971 , n11969 );
and ( n11973 , n11972 , n6474 );
or ( n11974 , n11970 , n11973 );
xor ( n11975 , n11967 , n11974 );
buf ( n11976 , n5981 );
xor ( n11977 , n11975 , n11976 );
buf ( n11978 , n5982 );
xor ( n11979 , n11977 , n11978 );
buf ( n11980 , n5983 );
xor ( n11981 , n11979 , n11980 );
xor ( n11982 , n11960 , n11981 );
and ( n11983 , n11952 , n11982 );
xor ( n11984 , n11928 , n11983 );
xor ( n11985 , n11910 , n11984 );
not ( n11986 , n6474 );
buf ( n11987 , n5984 );
and ( n11988 , n11986 , n11987 );
buf ( n11989 , n5985 );
xor ( n11990 , n11989 , n11987 );
and ( n11991 , n11990 , n6474 );
or ( n11992 , n11988 , n11991 );
xor ( n11993 , n7979 , n11992 );
buf ( n11994 , n5986 );
xor ( n11995 , n11993 , n11994 );
xor ( n11996 , n11995 , n10173 );
buf ( n11997 , n5987 );
xor ( n11998 , n11996 , n11997 );
xor ( n11999 , n11030 , n11998 );
xor ( n12000 , n11999 , n7521 );
xor ( n12001 , n11353 , n10044 );
xor ( n12002 , n12001 , n8891 );
not ( n12003 , n12002 );
not ( n12004 , n6474 );
buf ( n12005 , n5988 );
and ( n12006 , n12004 , n12005 );
buf ( n12007 , n5989 );
xor ( n12008 , n12007 , n12005 );
and ( n12009 , n12008 , n6474 );
or ( n12010 , n12006 , n12009 );
not ( n12011 , n6474 );
buf ( n12012 , n5990 );
and ( n12013 , n12011 , n12012 );
buf ( n12014 , n5991 );
xor ( n12015 , n12014 , n12012 );
and ( n12016 , n12015 , n6474 );
or ( n12017 , n12013 , n12016 );
xor ( n12018 , n12017 , n8807 );
buf ( n12019 , n5992 );
xor ( n12020 , n12018 , n12019 );
buf ( n12021 , n5993 );
xor ( n12022 , n12020 , n12021 );
buf ( n12023 , n5994 );
xor ( n12024 , n12022 , n12023 );
xor ( n12025 , n12010 , n12024 );
not ( n12026 , n6474 );
buf ( n12027 , n5995 );
and ( n12028 , n12026 , n12027 );
buf ( n12029 , n5996 );
xor ( n12030 , n12029 , n12027 );
and ( n12031 , n12030 , n6474 );
or ( n12032 , n12028 , n12031 );
buf ( n12033 , n5997 );
xor ( n12034 , n12032 , n12033 );
buf ( n12035 , n5998 );
xor ( n12036 , n12034 , n12035 );
buf ( n12037 , n5999 );
xor ( n12038 , n12036 , n12037 );
buf ( n12039 , n6000 );
xor ( n12040 , n12038 , n12039 );
xor ( n12041 , n12025 , n12040 );
and ( n12042 , n12003 , n12041 );
xor ( n12043 , n12000 , n12042 );
xor ( n12044 , n11985 , n12043 );
xor ( n12045 , n11720 , n12044 );
not ( n12046 , n6474 );
buf ( n12047 , n6001 );
and ( n12048 , n12046 , n12047 );
buf ( n12049 , n6002 );
xor ( n12050 , n12049 , n12047 );
and ( n12051 , n12050 , n6474 );
or ( n12052 , n12048 , n12051 );
not ( n12053 , n6474 );
buf ( n12054 , n6003 );
and ( n12055 , n12053 , n12054 );
buf ( n12056 , n6004 );
xor ( n12057 , n12056 , n12054 );
and ( n12058 , n12057 , n6474 );
or ( n12059 , n12055 , n12058 );
xor ( n12060 , n12052 , n12059 );
buf ( n12061 , n6005 );
xor ( n12062 , n12060 , n12061 );
buf ( n12063 , n6006 );
xor ( n12064 , n12062 , n12063 );
buf ( n12065 , n6007 );
xor ( n12066 , n12064 , n12065 );
xor ( n12067 , n10409 , n12066 );
xor ( n12068 , n12067 , n9895 );
buf ( n12069 , n6008 );
xor ( n12070 , n12069 , n8291 );
xor ( n12071 , n12070 , n9921 );
not ( n12072 , n12071 );
xor ( n12073 , n7858 , n11512 );
xor ( n12074 , n12073 , n11520 );
and ( n12075 , n12072 , n12074 );
xor ( n12076 , n12068 , n12075 );
not ( n12077 , n6474 );
buf ( n12078 , n6009 );
and ( n12079 , n12077 , n12078 );
buf ( n12080 , n6010 );
xor ( n12081 , n12080 , n12078 );
and ( n12082 , n12081 , n6474 );
or ( n12083 , n12079 , n12082 );
not ( n12084 , n6474 );
buf ( n12085 , n6011 );
and ( n12086 , n12084 , n12085 );
buf ( n12087 , n6012 );
xor ( n12088 , n12087 , n12085 );
and ( n12089 , n12088 , n6474 );
or ( n12090 , n12086 , n12089 );
xor ( n12091 , n12083 , n12090 );
buf ( n12092 , n6013 );
xor ( n12093 , n12091 , n12092 );
buf ( n12094 , n6014 );
xor ( n12095 , n12093 , n12094 );
buf ( n12096 , n6015 );
xor ( n12097 , n12095 , n12096 );
xor ( n12098 , n9141 , n12097 );
not ( n12099 , n6474 );
buf ( n12100 , n6016 );
and ( n12101 , n12099 , n12100 );
buf ( n12102 , n6017 );
xor ( n12103 , n12102 , n12100 );
and ( n12104 , n12103 , n6474 );
or ( n12105 , n12101 , n12104 );
xor ( n12106 , n12105 , n9592 );
buf ( n12107 , n6018 );
xor ( n12108 , n12106 , n12107 );
buf ( n12109 , n6019 );
xor ( n12110 , n12108 , n12109 );
xor ( n12111 , n12110 , n10937 );
xor ( n12112 , n12098 , n12111 );
xor ( n12113 , n8309 , n7537 );
xor ( n12114 , n12113 , n10905 );
not ( n12115 , n12114 );
xor ( n12116 , n8444 , n9942 );
xor ( n12117 , n12116 , n10193 );
and ( n12118 , n12115 , n12117 );
xor ( n12119 , n12112 , n12118 );
xor ( n12120 , n12076 , n12119 );
xor ( n12121 , n9332 , n6763 );
xor ( n12122 , n12121 , n6785 );
not ( n12123 , n6474 );
buf ( n12124 , n6020 );
and ( n12125 , n12123 , n12124 );
buf ( n12126 , n6021 );
xor ( n12127 , n12126 , n12124 );
and ( n12128 , n12127 , n6474 );
or ( n12129 , n12125 , n12128 );
not ( n12130 , n6474 );
buf ( n12131 , n6022 );
and ( n12132 , n12130 , n12131 );
buf ( n12133 , n6023 );
xor ( n12134 , n12133 , n12131 );
and ( n12135 , n12134 , n6474 );
or ( n12136 , n12132 , n12135 );
xor ( n12137 , n12129 , n12136 );
buf ( n12138 , n6024 );
xor ( n12139 , n12137 , n12138 );
buf ( n12140 , n6025 );
xor ( n12141 , n12139 , n12140 );
buf ( n12142 , n6026 );
xor ( n12143 , n12141 , n12142 );
xor ( n12144 , n7001 , n12143 );
xor ( n12145 , n12144 , n9710 );
not ( n12146 , n12145 );
buf ( n12147 , n6027 );
xor ( n12148 , n12147 , n7331 );
not ( n12149 , n6474 );
buf ( n12150 , n6028 );
and ( n12151 , n12149 , n12150 );
buf ( n12152 , n6029 );
xor ( n12153 , n12152 , n12150 );
and ( n12154 , n12153 , n6474 );
or ( n12155 , n12151 , n12154 );
xor ( n12156 , n6569 , n12155 );
buf ( n12157 , n6030 );
xor ( n12158 , n12156 , n12157 );
buf ( n12159 , n6031 );
xor ( n12160 , n12158 , n12159 );
buf ( n12161 , n6032 );
xor ( n12162 , n12160 , n12161 );
xor ( n12163 , n12148 , n12162 );
and ( n12164 , n12146 , n12163 );
xor ( n12165 , n12122 , n12164 );
xor ( n12166 , n12120 , n12165 );
xor ( n12167 , n11651 , n11405 );
xor ( n12168 , n12167 , n11427 );
xor ( n12169 , n6601 , n8076 );
not ( n12170 , n6474 );
buf ( n12171 , n6033 );
and ( n12172 , n12170 , n12171 );
buf ( n12173 , n6034 );
xor ( n12174 , n12173 , n12171 );
and ( n12175 , n12174 , n6474 );
or ( n12176 , n12172 , n12175 );
not ( n12177 , n6474 );
buf ( n12178 , n6035 );
and ( n12179 , n12177 , n12178 );
buf ( n12180 , n6036 );
xor ( n12181 , n12180 , n12178 );
and ( n12182 , n12181 , n6474 );
or ( n12183 , n12179 , n12182 );
xor ( n12184 , n12176 , n12183 );
buf ( n12185 , n6037 );
xor ( n12186 , n12184 , n12185 );
buf ( n12187 , n6038 );
xor ( n12188 , n12186 , n12187 );
buf ( n12189 , n6039 );
xor ( n12190 , n12188 , n12189 );
xor ( n12191 , n12169 , n12190 );
not ( n12192 , n12191 );
not ( n12193 , n6474 );
buf ( n12194 , n6040 );
and ( n12195 , n12193 , n12194 );
buf ( n12196 , n6041 );
xor ( n12197 , n12196 , n12194 );
and ( n12198 , n12197 , n6474 );
or ( n12199 , n12195 , n12198 );
not ( n12200 , n6474 );
buf ( n12201 , n6042 );
and ( n12202 , n12200 , n12201 );
buf ( n12203 , n6043 );
xor ( n12204 , n12203 , n12201 );
and ( n12205 , n12204 , n6474 );
or ( n12206 , n12202 , n12205 );
xor ( n12207 , n12199 , n12206 );
buf ( n12208 , n6044 );
xor ( n12209 , n12207 , n12208 );
buf ( n12210 , n6045 );
xor ( n12211 , n12209 , n12210 );
buf ( n12212 , n6046 );
xor ( n12213 , n12211 , n12212 );
xor ( n12214 , n10127 , n12213 );
xor ( n12215 , n12214 , n10768 );
and ( n12216 , n12192 , n12215 );
xor ( n12217 , n12168 , n12216 );
xor ( n12218 , n12166 , n12217 );
xor ( n12219 , n8835 , n6739 );
xor ( n12220 , n12219 , n11927 );
xor ( n12221 , n7371 , n10224 );
xor ( n12222 , n12221 , n10246 );
not ( n12223 , n12222 );
buf ( n12224 , n6047 );
xor ( n12225 , n12224 , n9094 );
not ( n12226 , n6474 );
buf ( n12227 , n6048 );
and ( n12228 , n12226 , n12227 );
buf ( n12229 , n6049 );
xor ( n12230 , n12229 , n12227 );
and ( n12231 , n12230 , n6474 );
or ( n12232 , n12228 , n12231 );
not ( n12233 , n6474 );
buf ( n12234 , n6050 );
and ( n12235 , n12233 , n12234 );
buf ( n12236 , n6051 );
xor ( n12237 , n12236 , n12234 );
and ( n12238 , n12237 , n6474 );
or ( n12239 , n12235 , n12238 );
xor ( n12240 , n12232 , n12239 );
buf ( n12241 , n6052 );
xor ( n12242 , n12240 , n12241 );
buf ( n12243 , n6053 );
xor ( n12244 , n12242 , n12243 );
buf ( n12245 , n6054 );
xor ( n12246 , n12244 , n12245 );
xor ( n12247 , n12225 , n12246 );
and ( n12248 , n12223 , n12247 );
xor ( n12249 , n12220 , n12248 );
xor ( n12250 , n12218 , n12249 );
xor ( n12251 , n12045 , n12250 );
not ( n12252 , n6474 );
buf ( n12253 , n6055 );
and ( n12254 , n12252 , n12253 );
buf ( n12255 , n6056 );
xor ( n12256 , n12255 , n12253 );
and ( n12257 , n12256 , n6474 );
or ( n12258 , n12254 , n12257 );
xor ( n12259 , n12258 , n9002 );
xor ( n12260 , n12259 , n11329 );
not ( n12261 , n6474 );
buf ( n12262 , n6057 );
and ( n12263 , n12261 , n12262 );
buf ( n12264 , n6058 );
xor ( n12265 , n12264 , n12262 );
and ( n12266 , n12265 , n6474 );
or ( n12267 , n12263 , n12266 );
not ( n12268 , n6474 );
buf ( n12269 , n6059 );
and ( n12270 , n12268 , n12269 );
buf ( n12271 , n6060 );
xor ( n12272 , n12271 , n12269 );
and ( n12273 , n12272 , n6474 );
or ( n12274 , n12270 , n12273 );
xor ( n12275 , n12267 , n12274 );
buf ( n12276 , n6061 );
xor ( n12277 , n12275 , n12276 );
buf ( n12278 , n6062 );
xor ( n12279 , n12277 , n12278 );
buf ( n12280 , n6063 );
xor ( n12281 , n12279 , n12280 );
xor ( n12282 , n7129 , n12281 );
not ( n12283 , n6474 );
buf ( n12284 , n6064 );
and ( n12285 , n12283 , n12284 );
buf ( n12286 , n6065 );
xor ( n12287 , n12286 , n12284 );
and ( n12288 , n12287 , n6474 );
or ( n12289 , n12285 , n12288 );
not ( n12290 , n6474 );
buf ( n12291 , n6066 );
and ( n12292 , n12290 , n12291 );
buf ( n12293 , n6067 );
xor ( n12294 , n12293 , n12291 );
and ( n12295 , n12294 , n6474 );
or ( n12296 , n12292 , n12295 );
xor ( n12297 , n12289 , n12296 );
xor ( n12298 , n12297 , n6610 );
buf ( n12299 , n6068 );
xor ( n12300 , n12298 , n12299 );
buf ( n12301 , n6069 );
xor ( n12302 , n12300 , n12301 );
xor ( n12303 , n12282 , n12302 );
not ( n12304 , n12303 );
buf ( n12305 , n6070 );
xor ( n12306 , n12305 , n11275 );
xor ( n12307 , n12306 , n9559 );
and ( n12308 , n12304 , n12307 );
xor ( n12309 , n12260 , n12308 );
not ( n12310 , n6474 );
buf ( n12311 , n6071 );
and ( n12312 , n12310 , n12311 );
buf ( n12313 , n6072 );
xor ( n12314 , n12313 , n12311 );
and ( n12315 , n12314 , n6474 );
or ( n12316 , n12312 , n12315 );
xor ( n12317 , n12316 , n9094 );
xor ( n12318 , n12317 , n12246 );
xor ( n12319 , n9163 , n12111 );
xor ( n12320 , n12319 , n7910 );
not ( n12321 , n12320 );
xor ( n12322 , n6956 , n8114 );
xor ( n12323 , n12322 , n7861 );
and ( n12324 , n12321 , n12323 );
xor ( n12325 , n12318 , n12324 );
xor ( n12326 , n9364 , n9872 );
not ( n12327 , n6474 );
buf ( n12328 , n6073 );
and ( n12329 , n12327 , n12328 );
buf ( n12330 , n6074 );
xor ( n12331 , n12330 , n12328 );
and ( n12332 , n12331 , n6474 );
or ( n12333 , n12329 , n12332 );
buf ( n12334 , n6075 );
xor ( n12335 , n12333 , n12334 );
buf ( n12336 , n6076 );
xor ( n12337 , n12335 , n12336 );
buf ( n12338 , n6077 );
xor ( n12339 , n12337 , n12338 );
buf ( n12340 , n6078 );
xor ( n12341 , n12339 , n12340 );
xor ( n12342 , n12326 , n12341 );
buf ( n12343 , n6079 );
xor ( n12344 , n12343 , n11833 );
not ( n12345 , n6474 );
buf ( n12346 , n6080 );
and ( n12347 , n12345 , n12346 );
buf ( n12348 , n6081 );
xor ( n12349 , n12348 , n12346 );
and ( n12350 , n12349 , n6474 );
or ( n12351 , n12347 , n12350 );
not ( n12352 , n6474 );
buf ( n12353 , n6082 );
and ( n12354 , n12352 , n12353 );
buf ( n12355 , n6083 );
xor ( n12356 , n12355 , n12353 );
and ( n12357 , n12356 , n6474 );
or ( n12358 , n12354 , n12357 );
xor ( n12359 , n12351 , n12358 );
buf ( n12360 , n6084 );
xor ( n12361 , n12359 , n12360 );
buf ( n12362 , n6085 );
xor ( n12363 , n12361 , n12362 );
buf ( n12364 , n6086 );
xor ( n12365 , n12363 , n12364 );
xor ( n12366 , n12344 , n12365 );
not ( n12367 , n12366 );
not ( n12368 , n6474 );
buf ( n12369 , n6087 );
and ( n12370 , n12368 , n12369 );
buf ( n12371 , n6088 );
xor ( n12372 , n12371 , n12369 );
and ( n12373 , n12372 , n6474 );
or ( n12374 , n12370 , n12373 );
xor ( n12375 , n12374 , n9900 );
buf ( n12376 , n6089 );
xor ( n12377 , n12375 , n12376 );
buf ( n12378 , n6090 );
xor ( n12379 , n12377 , n12378 );
buf ( n12380 , n6091 );
xor ( n12381 , n12379 , n12380 );
xor ( n12382 , n12061 , n12381 );
xor ( n12383 , n12382 , n8447 );
and ( n12384 , n12367 , n12383 );
xor ( n12385 , n12342 , n12384 );
xor ( n12386 , n12325 , n12385 );
xor ( n12387 , n12232 , n8764 );
not ( n12388 , n6474 );
buf ( n12389 , n6092 );
and ( n12390 , n12388 , n12389 );
buf ( n12391 , n6093 );
xor ( n12392 , n12391 , n12389 );
and ( n12393 , n12392 , n6474 );
or ( n12394 , n12390 , n12393 );
not ( n12395 , n6474 );
buf ( n12396 , n6094 );
and ( n12397 , n12395 , n12396 );
buf ( n12398 , n6095 );
xor ( n12399 , n12398 , n12396 );
and ( n12400 , n12399 , n6474 );
or ( n12401 , n12397 , n12400 );
xor ( n12402 , n12394 , n12401 );
xor ( n12403 , n12402 , n12069 );
buf ( n12404 , n6096 );
xor ( n12405 , n12403 , n12404 );
buf ( n12406 , n6097 );
xor ( n12407 , n12405 , n12406 );
xor ( n12408 , n12387 , n12407 );
xor ( n12409 , n8049 , n7634 );
xor ( n12410 , n12409 , n7072 );
not ( n12411 , n12410 );
xor ( n12412 , n11048 , n7521 );
xor ( n12413 , n12412 , n7537 );
and ( n12414 , n12411 , n12413 );
xor ( n12415 , n12408 , n12414 );
xor ( n12416 , n12386 , n12415 );
not ( n12417 , n6474 );
buf ( n12418 , n6098 );
and ( n12419 , n12417 , n12418 );
buf ( n12420 , n6099 );
xor ( n12421 , n12420 , n12418 );
and ( n12422 , n12421 , n6474 );
or ( n12423 , n12419 , n12422 );
xor ( n12424 , n12423 , n9026 );
xor ( n12425 , n12424 , n9047 );
not ( n12426 , n12260 );
and ( n12427 , n12426 , n12303 );
xor ( n12428 , n12425 , n12427 );
xor ( n12429 , n12416 , n12428 );
xor ( n12430 , n9276 , n8660 );
xor ( n12431 , n12430 , n10105 );
not ( n12432 , n6474 );
buf ( n12433 , n6100 );
and ( n12434 , n12432 , n12433 );
buf ( n12435 , n6101 );
xor ( n12436 , n12435 , n12433 );
and ( n12437 , n12436 , n6474 );
or ( n12438 , n12434 , n12437 );
not ( n12439 , n6474 );
buf ( n12440 , n6102 );
and ( n12441 , n12439 , n12440 );
buf ( n12442 , n6103 );
xor ( n12443 , n12442 , n12440 );
and ( n12444 , n12443 , n6474 );
or ( n12445 , n12441 , n12444 );
xor ( n12446 , n12438 , n12445 );
buf ( n12447 , n6104 );
xor ( n12448 , n12446 , n12447 );
buf ( n12449 , n6105 );
xor ( n12450 , n12448 , n12449 );
buf ( n12451 , n6106 );
xor ( n12452 , n12450 , n12451 );
xor ( n12453 , n9787 , n12452 );
not ( n12454 , n6474 );
buf ( n12455 , n6107 );
and ( n12456 , n12454 , n12455 );
buf ( n12457 , n6108 );
xor ( n12458 , n12457 , n12455 );
and ( n12459 , n12458 , n6474 );
or ( n12460 , n12456 , n12459 );
buf ( n12461 , n6109 );
xor ( n12462 , n12460 , n12461 );
buf ( n12463 , n6110 );
xor ( n12464 , n12462 , n12463 );
xor ( n12465 , n12464 , n10355 );
buf ( n12466 , n6111 );
xor ( n12467 , n12465 , n12466 );
xor ( n12468 , n12453 , n12467 );
not ( n12469 , n12468 );
xor ( n12470 , n10141 , n10768 );
xor ( n12471 , n12470 , n10790 );
and ( n12472 , n12469 , n12471 );
xor ( n12473 , n12431 , n12472 );
xor ( n12474 , n12429 , n12473 );
xor ( n12475 , n12309 , n12474 );
xor ( n12476 , n11507 , n9170 );
xor ( n12477 , n12476 , n8495 );
not ( n12478 , n6474 );
buf ( n12479 , n6112 );
and ( n12480 , n12478 , n12479 );
buf ( n12481 , n6113 );
xor ( n12482 , n12481 , n12479 );
and ( n12483 , n12482 , n6474 );
or ( n12484 , n12480 , n12483 );
xor ( n12485 , n8345 , n12484 );
buf ( n12486 , n6114 );
xor ( n12487 , n12485 , n12486 );
buf ( n12488 , n6115 );
xor ( n12489 , n12487 , n12488 );
xor ( n12490 , n12489 , n10839 );
xor ( n12491 , n7790 , n12490 );
not ( n12492 , n6474 );
buf ( n12493 , n6116 );
and ( n12494 , n12492 , n12493 );
buf ( n12495 , n6117 );
xor ( n12496 , n12495 , n12493 );
and ( n12497 , n12496 , n6474 );
or ( n12498 , n12494 , n12497 );
buf ( n12499 , n6118 );
xor ( n12500 , n12498 , n12499 );
buf ( n12501 , n6119 );
xor ( n12502 , n12500 , n12501 );
buf ( n12503 , n6120 );
xor ( n12504 , n12502 , n12503 );
buf ( n12505 , n6121 );
xor ( n12506 , n12504 , n12505 );
xor ( n12507 , n12491 , n12506 );
not ( n12508 , n12507 );
xor ( n12509 , n11926 , n9511 );
not ( n12510 , n6474 );
buf ( n12511 , n6122 );
and ( n12512 , n12510 , n12511 );
buf ( n12513 , n6123 );
xor ( n12514 , n12513 , n12511 );
and ( n12515 , n12514 , n6474 );
or ( n12516 , n12512 , n12515 );
not ( n12517 , n6474 );
buf ( n12518 , n6124 );
and ( n12519 , n12517 , n12518 );
buf ( n12520 , n6125 );
xor ( n12521 , n12520 , n12518 );
and ( n12522 , n12521 , n6474 );
or ( n12523 , n12519 , n12522 );
xor ( n12524 , n12516 , n12523 );
buf ( n12525 , n6126 );
xor ( n12526 , n12524 , n12525 );
buf ( n12527 , n6127 );
xor ( n12528 , n12526 , n12527 );
buf ( n12529 , n6128 );
xor ( n12530 , n12528 , n12529 );
xor ( n12531 , n12509 , n12530 );
and ( n12532 , n12508 , n12531 );
xor ( n12533 , n12477 , n12532 );
not ( n12534 , n6474 );
buf ( n12535 , n6129 );
and ( n12536 , n12534 , n12535 );
buf ( n12537 , n6130 );
xor ( n12538 , n12537 , n12535 );
and ( n12539 , n12538 , n6474 );
or ( n12540 , n12536 , n12539 );
buf ( n12541 , n6131 );
xor ( n12542 , n12540 , n12541 );
buf ( n12543 , n6132 );
xor ( n12544 , n12542 , n12543 );
buf ( n12545 , n6133 );
xor ( n12546 , n12544 , n12545 );
buf ( n12547 , n6134 );
xor ( n12548 , n12546 , n12547 );
xor ( n12549 , n9937 , n12548 );
xor ( n12550 , n12549 , n9238 );
xor ( n12551 , n10622 , n8517 );
xor ( n12552 , n12551 , n11462 );
not ( n12553 , n12552 );
xor ( n12554 , n9289 , n8660 );
xor ( n12555 , n12554 , n10105 );
and ( n12556 , n12553 , n12555 );
xor ( n12557 , n12550 , n12556 );
xor ( n12558 , n12533 , n12557 );
xor ( n12559 , n11299 , n8159 );
xor ( n12560 , n12423 , n9005 );
buf ( n12561 , n6135 );
xor ( n12562 , n12560 , n12561 );
buf ( n12563 , n6136 );
xor ( n12564 , n12562 , n12563 );
buf ( n12565 , n6137 );
xor ( n12566 , n12564 , n12565 );
xor ( n12567 , n12559 , n12566 );
not ( n12568 , n6474 );
buf ( n12569 , n6138 );
and ( n12570 , n12568 , n12569 );
buf ( n12571 , n6139 );
xor ( n12572 , n12571 , n12569 );
and ( n12573 , n12572 , n6474 );
or ( n12574 , n12570 , n12573 );
xor ( n12575 , n12574 , n11155 );
buf ( n12576 , n6140 );
xor ( n12577 , n12575 , n12576 );
buf ( n12578 , n6141 );
xor ( n12579 , n12577 , n12578 );
buf ( n12580 , n6142 );
xor ( n12581 , n12579 , n12580 );
xor ( n12582 , n7109 , n12581 );
xor ( n12583 , n12582 , n12281 );
not ( n12584 , n12583 );
xor ( n12585 , n11344 , n10022 );
xor ( n12586 , n12585 , n10044 );
and ( n12587 , n12584 , n12586 );
xor ( n12588 , n12567 , n12587 );
xor ( n12589 , n12558 , n12588 );
not ( n12590 , n6474 );
buf ( n12591 , n6143 );
and ( n12592 , n12590 , n12591 );
buf ( n12593 , n6144 );
xor ( n12594 , n12593 , n12591 );
and ( n12595 , n12594 , n6474 );
or ( n12596 , n12592 , n12595 );
not ( n12597 , n6474 );
buf ( n12598 , n6145 );
and ( n12599 , n12597 , n12598 );
buf ( n12600 , n6146 );
xor ( n12601 , n12600 , n12598 );
and ( n12602 , n12601 , n6474 );
or ( n12603 , n12599 , n12602 );
xor ( n12604 , n12596 , n12603 );
xor ( n12605 , n12604 , n9402 );
buf ( n12606 , n6147 );
xor ( n12607 , n12605 , n12606 );
buf ( n12608 , n6148 );
xor ( n12609 , n12607 , n12608 );
xor ( n12610 , n6626 , n12609 );
xor ( n12611 , n12610 , n10334 );
xor ( n12612 , n8185 , n11132 );
xor ( n12613 , n12612 , n11146 );
not ( n12614 , n12613 );
buf ( n12615 , n6149 );
xor ( n12616 , n12615 , n6811 );
xor ( n12617 , n12616 , n6827 );
and ( n12618 , n12614 , n12617 );
xor ( n12619 , n12611 , n12618 );
xor ( n12620 , n12589 , n12619 );
xor ( n12621 , n11198 , n6850 );
xor ( n12622 , n12621 , n6872 );
xor ( n12623 , n6936 , n8092 );
xor ( n12624 , n12623 , n8114 );
not ( n12625 , n12624 );
xor ( n12626 , n10415 , n12066 );
xor ( n12627 , n12626 , n9895 );
and ( n12628 , n12625 , n12627 );
xor ( n12629 , n12622 , n12628 );
xor ( n12630 , n12620 , n12629 );
xor ( n12631 , n12475 , n12630 );
not ( n12632 , n12631 );
xor ( n12633 , n10925 , n9794 );
xor ( n12634 , n12633 , n9816 );
not ( n12635 , n6474 );
buf ( n12636 , n6150 );
and ( n12637 , n12635 , n12636 );
buf ( n12638 , n6151 );
xor ( n12639 , n12638 , n12636 );
and ( n12640 , n12639 , n6474 );
or ( n12641 , n12637 , n12640 );
buf ( n12642 , n6152 );
xor ( n12643 , n12641 , n12642 );
buf ( n12644 , n6153 );
xor ( n12645 , n12643 , n12644 );
buf ( n12646 , n6154 );
xor ( n12647 , n12645 , n12646 );
buf ( n12648 , n6155 );
xor ( n12649 , n12647 , n12648 );
xor ( n12650 , n10064 , n12649 );
not ( n12651 , n6474 );
buf ( n12652 , n6156 );
and ( n12653 , n12651 , n12652 );
buf ( n12654 , n6157 );
xor ( n12655 , n12654 , n12652 );
and ( n12656 , n12655 , n6474 );
or ( n12657 , n12653 , n12656 );
not ( n12658 , n6474 );
buf ( n12659 , n6158 );
and ( n12660 , n12658 , n12659 );
buf ( n12661 , n6159 );
xor ( n12662 , n12661 , n12659 );
and ( n12663 , n12662 , n6474 );
or ( n12664 , n12660 , n12663 );
xor ( n12665 , n12657 , n12664 );
buf ( n12666 , n6160 );
xor ( n12667 , n12665 , n12666 );
buf ( n12668 , n6161 );
xor ( n12669 , n12667 , n12668 );
buf ( n12670 , n6162 );
xor ( n12671 , n12669 , n12670 );
xor ( n12672 , n12650 , n12671 );
not ( n12673 , n12672 );
buf ( n12674 , n6163 );
xor ( n12675 , n12674 , n9651 );
xor ( n12676 , n12675 , n9673 );
and ( n12677 , n12673 , n12676 );
xor ( n12678 , n12634 , n12677 );
not ( n12679 , n6474 );
buf ( n12680 , n6164 );
and ( n12681 , n12679 , n12680 );
buf ( n12682 , n6165 );
xor ( n12683 , n12682 , n12680 );
and ( n12684 , n12683 , n6474 );
or ( n12685 , n12681 , n12684 );
not ( n12686 , n6474 );
buf ( n12687 , n6166 );
and ( n12688 , n12686 , n12687 );
buf ( n12689 , n6167 );
xor ( n12690 , n12689 , n12687 );
and ( n12691 , n12690 , n6474 );
or ( n12692 , n12688 , n12691 );
xor ( n12693 , n12685 , n12692 );
buf ( n12694 , n6168 );
xor ( n12695 , n12693 , n12694 );
buf ( n12696 , n6169 );
xor ( n12697 , n12695 , n12696 );
buf ( n12698 , n6170 );
xor ( n12699 , n12697 , n12698 );
xor ( n12700 , n11420 , n12699 );
xor ( n12701 , n12700 , n7360 );
buf ( n12702 , n6171 );
xor ( n12703 , n12702 , n11981 );
xor ( n12704 , n12703 , n7566 );
not ( n12705 , n12704 );
buf ( n12706 , n6172 );
not ( n12707 , n6474 );
buf ( n12708 , n6173 );
and ( n12709 , n12707 , n12708 );
buf ( n12710 , n6174 );
xor ( n12711 , n12710 , n12708 );
and ( n12712 , n12711 , n6474 );
or ( n12713 , n12709 , n12712 );
not ( n12714 , n6474 );
buf ( n12715 , n6175 );
and ( n12716 , n12714 , n12715 );
buf ( n12717 , n6176 );
xor ( n12718 , n12717 , n12715 );
and ( n12719 , n12718 , n6474 );
or ( n12720 , n12716 , n12719 );
xor ( n12721 , n12713 , n12720 );
buf ( n12722 , n6177 );
xor ( n12723 , n12721 , n12722 );
buf ( n12724 , n6178 );
xor ( n12725 , n12723 , n12724 );
buf ( n12726 , n6179 );
xor ( n12727 , n12725 , n12726 );
xor ( n12728 , n12706 , n12727 );
not ( n12729 , n6474 );
buf ( n12730 , n6180 );
and ( n12731 , n12729 , n12730 );
buf ( n12732 , n6181 );
xor ( n12733 , n12732 , n12730 );
and ( n12734 , n12733 , n6474 );
or ( n12735 , n12731 , n12734 );
buf ( n12736 , n6182 );
xor ( n12737 , n12735 , n12736 );
buf ( n12738 , n6183 );
xor ( n12739 , n12737 , n12738 );
buf ( n12740 , n6184 );
xor ( n12741 , n12739 , n12740 );
xor ( n12742 , n12741 , n7927 );
xor ( n12743 , n12728 , n12742 );
and ( n12744 , n12705 , n12743 );
xor ( n12745 , n12701 , n12744 );
xor ( n12746 , n8995 , n11741 );
xor ( n12747 , n12746 , n11763 );
xor ( n12748 , n11340 , n10022 );
xor ( n12749 , n12748 , n10044 );
not ( n12750 , n12749 );
buf ( n12751 , n6185 );
xor ( n12752 , n12751 , n7588 );
xor ( n12753 , n12752 , n9290 );
and ( n12754 , n12750 , n12753 );
xor ( n12755 , n12747 , n12754 );
xor ( n12756 , n12745 , n12755 );
xor ( n12757 , n12484 , n8366 );
xor ( n12758 , n12757 , n8388 );
not ( n12759 , n6474 );
buf ( n12760 , n6186 );
and ( n12761 , n12759 , n12760 );
buf ( n12762 , n6187 );
xor ( n12763 , n12762 , n12760 );
and ( n12764 , n12763 , n6474 );
or ( n12765 , n12761 , n12764 );
not ( n12766 , n6474 );
buf ( n12767 , n6188 );
and ( n12768 , n12766 , n12767 );
buf ( n12769 , n6189 );
xor ( n12770 , n12769 , n12767 );
and ( n12771 , n12770 , n6474 );
or ( n12772 , n12768 , n12771 );
xor ( n12773 , n12765 , n12772 );
buf ( n12774 , n6190 );
xor ( n12775 , n12773 , n12774 );
buf ( n12776 , n6191 );
xor ( n12777 , n12775 , n12776 );
buf ( n12778 , n6192 );
xor ( n12779 , n12777 , n12778 );
xor ( n12780 , n10669 , n12779 );
xor ( n12781 , n12780 , n8092 );
not ( n12782 , n12781 );
xor ( n12783 , n7991 , n8710 );
xor ( n12784 , n12783 , n8137 );
and ( n12785 , n12782 , n12784 );
xor ( n12786 , n12758 , n12785 );
xor ( n12787 , n12756 , n12786 );
buf ( n12788 , n6193 );
xor ( n12789 , n8586 , n12788 );
buf ( n12790 , n6194 );
xor ( n12791 , n12789 , n12790 );
buf ( n12792 , n6195 );
xor ( n12793 , n12791 , n12792 );
buf ( n12794 , n6196 );
xor ( n12795 , n12793 , n12794 );
xor ( n12796 , n8242 , n12795 );
xor ( n12797 , n12796 , n9973 );
xor ( n12798 , n8410 , n8314 );
xor ( n12799 , n12798 , n8336 );
not ( n12800 , n12799 );
buf ( n12801 , n6197 );
xor ( n12802 , n12801 , n7710 );
xor ( n12803 , n12802 , n7732 );
and ( n12804 , n12800 , n12803 );
xor ( n12805 , n12797 , n12804 );
xor ( n12806 , n12787 , n12805 );
xor ( n12807 , n7065 , n10836 );
not ( n12808 , n6474 );
buf ( n12809 , n6198 );
and ( n12810 , n12808 , n12809 );
buf ( n12811 , n6199 );
xor ( n12812 , n12811 , n12809 );
and ( n12813 , n12812 , n6474 );
or ( n12814 , n12810 , n12813 );
buf ( n12815 , n6200 );
xor ( n12816 , n12814 , n12815 );
buf ( n12817 , n6201 );
xor ( n12818 , n12816 , n12817 );
buf ( n12819 , n6202 );
xor ( n12820 , n12818 , n12819 );
buf ( n12821 , n6203 );
xor ( n12822 , n12820 , n12821 );
xor ( n12823 , n12807 , n12822 );
not ( n12824 , n12634 );
and ( n12825 , n12824 , n12672 );
xor ( n12826 , n12823 , n12825 );
xor ( n12827 , n12806 , n12826 );
xor ( n12828 , n12678 , n12827 );
xor ( n12829 , n7945 , n10130 );
xor ( n12830 , n12829 , n10146 );
buf ( n12831 , n6204 );
xor ( n12832 , n12831 , n7331 );
xor ( n12833 , n12832 , n12162 );
not ( n12834 , n12833 );
xor ( n12835 , n9567 , n8204 );
not ( n12836 , n6474 );
buf ( n12837 , n6205 );
and ( n12838 , n12836 , n12837 );
buf ( n12839 , n6206 );
xor ( n12840 , n12839 , n12837 );
and ( n12841 , n12840 , n6474 );
or ( n12842 , n12838 , n12841 );
not ( n12843 , n6474 );
buf ( n12844 , n6207 );
and ( n12845 , n12843 , n12844 );
buf ( n12846 , n6208 );
xor ( n12847 , n12846 , n12844 );
and ( n12848 , n12847 , n6474 );
or ( n12849 , n12845 , n12848 );
xor ( n12850 , n12842 , n12849 );
xor ( n12851 , n12850 , n9630 );
buf ( n12852 , n6209 );
xor ( n12853 , n12851 , n12852 );
xor ( n12854 , n12853 , n12674 );
xor ( n12855 , n12835 , n12854 );
and ( n12856 , n12834 , n12855 );
xor ( n12857 , n12830 , n12856 );
not ( n12858 , n6474 );
buf ( n12859 , n6210 );
and ( n12860 , n12858 , n12859 );
buf ( n12861 , n6211 );
xor ( n12862 , n12861 , n12859 );
and ( n12863 , n12862 , n6474 );
or ( n12864 , n12860 , n12863 );
xor ( n12865 , n12864 , n11002 );
buf ( n12866 , n6212 );
xor ( n12867 , n12865 , n12866 );
buf ( n12868 , n6213 );
xor ( n12869 , n12867 , n12868 );
buf ( n12870 , n6214 );
xor ( n12871 , n12869 , n12870 );
xor ( n12872 , n8657 , n12871 );
xor ( n12873 , n12872 , n9079 );
xor ( n12874 , n6738 , n9489 );
xor ( n12875 , n12874 , n9511 );
not ( n12876 , n12875 );
xor ( n12877 , n8482 , n7910 );
xor ( n12878 , n12877 , n7925 );
and ( n12879 , n12876 , n12878 );
xor ( n12880 , n12873 , n12879 );
xor ( n12881 , n12857 , n12880 );
xor ( n12882 , n7043 , n11052 );
xor ( n12883 , n12882 , n8314 );
xor ( n12884 , n7658 , n6673 );
xor ( n12885 , n12884 , n6695 );
not ( n12886 , n12885 );
xor ( n12887 , n12842 , n9651 );
xor ( n12888 , n12887 , n9673 );
and ( n12889 , n12886 , n12888 );
xor ( n12890 , n12883 , n12889 );
xor ( n12891 , n12881 , n12890 );
xor ( n12892 , n8862 , n10963 );
xor ( n12893 , n12892 , n10864 );
xor ( n12894 , n12580 , n8799 );
xor ( n12895 , n12894 , n11171 );
not ( n12896 , n12895 );
xor ( n12897 , n9599 , n7861 );
xor ( n12898 , n12897 , n7883 );
and ( n12899 , n12896 , n12898 );
xor ( n12900 , n12893 , n12899 );
xor ( n12901 , n12891 , n12900 );
buf ( n12902 , n6215 );
xor ( n12903 , n12902 , n6827 );
xor ( n12904 , n12903 , n11981 );
xor ( n12905 , n11226 , n11345 );
xor ( n12906 , n12905 , n11367 );
not ( n12907 , n12906 );
not ( n12908 , n6474 );
buf ( n12909 , n6216 );
and ( n12910 , n12908 , n12909 );
buf ( n12911 , n6217 );
xor ( n12912 , n12911 , n12909 );
and ( n12913 , n12912 , n6474 );
or ( n12914 , n12910 , n12913 );
xor ( n12915 , n12914 , n11275 );
xor ( n12916 , n12915 , n9559 );
and ( n12917 , n12907 , n12916 );
xor ( n12918 , n12904 , n12917 );
xor ( n12919 , n12901 , n12918 );
xor ( n12920 , n12828 , n12919 );
and ( n12921 , n12632 , n12920 );
xor ( n12922 , n12251 , n12921 );
and ( n12923 , n12922 , n6475 );
or ( n12924 , n11672 , n12923 );
and ( n12925 , n11670 , n12924 );
buf ( n12926 , n12925 );
buf ( n12927 , n12926 );
not ( n12928 , n6469 );
not ( n12929 , n6475 );
and ( n12930 , n12929 , n10437 );
not ( n12931 , n9897 );
not ( n12932 , n6474 );
buf ( n12933 , n6218 );
and ( n12934 , n12932 , n12933 );
buf ( n12935 , n6219 );
xor ( n12936 , n12935 , n12933 );
and ( n12937 , n12936 , n6474 );
or ( n12938 , n12934 , n12937 );
xor ( n12939 , n7339 , n12938 );
buf ( n12940 , n6220 );
xor ( n12941 , n12939 , n12940 );
buf ( n12942 , n6221 );
xor ( n12943 , n12941 , n12942 );
buf ( n12944 , n6222 );
xor ( n12945 , n12943 , n12944 );
xor ( n12946 , n8637 , n12945 );
xor ( n12947 , n12946 , n12871 );
and ( n12948 , n12931 , n12947 );
xor ( n12949 , n9875 , n12948 );
xor ( n12950 , n12949 , n10178 );
xor ( n12951 , n12950 , n10630 );
xor ( n12952 , n7768 , n12365 );
xor ( n12953 , n12952 , n12490 );
xor ( n12954 , n12726 , n11329 );
xor ( n12955 , n12954 , n7948 );
not ( n12956 , n12955 );
not ( n12957 , n6474 );
buf ( n12958 , n6223 );
and ( n12959 , n12957 , n12958 );
buf ( n12960 , n6224 );
xor ( n12961 , n12960 , n12958 );
and ( n12962 , n12961 , n6474 );
or ( n12963 , n12959 , n12962 );
xor ( n12964 , n12963 , n9895 );
xor ( n12965 , n12964 , n7612 );
and ( n12966 , n12956 , n12965 );
xor ( n12967 , n12953 , n12966 );
xor ( n12968 , n9668 , n11227 );
xor ( n12969 , n12968 , n11833 );
xor ( n12970 , n12942 , n7360 );
xor ( n12971 , n12970 , n7376 );
not ( n12972 , n12971 );
xor ( n12973 , n6515 , n9995 );
not ( n12974 , n6474 );
buf ( n12975 , n6225 );
and ( n12976 , n12974 , n12975 );
buf ( n12977 , n6226 );
xor ( n12978 , n12977 , n12975 );
and ( n12979 , n12978 , n6474 );
or ( n12980 , n12976 , n12979 );
xor ( n12981 , n12980 , n11533 );
buf ( n12982 , n6227 );
xor ( n12983 , n12981 , n12982 );
buf ( n12984 , n6228 );
xor ( n12985 , n12983 , n12984 );
buf ( n12986 , n6229 );
xor ( n12987 , n12985 , n12986 );
xor ( n12988 , n12973 , n12987 );
and ( n12989 , n12972 , n12988 );
xor ( n12990 , n12969 , n12989 );
xor ( n12991 , n11875 , n9148 );
xor ( n12992 , n12991 , n9170 );
not ( n12993 , n12953 );
and ( n12994 , n12993 , n12955 );
xor ( n12995 , n12992 , n12994 );
xor ( n12996 , n12990 , n12995 );
buf ( n12997 , n6230 );
not ( n12998 , n6474 );
buf ( n12999 , n6231 );
and ( n13000 , n12998 , n12999 );
buf ( n13001 , n6232 );
xor ( n13002 , n13001 , n12999 );
and ( n13003 , n13002 , n6474 );
or ( n13004 , n13000 , n13003 );
not ( n13005 , n6474 );
buf ( n13006 , n6233 );
and ( n13007 , n13005 , n13006 );
buf ( n13008 , n6234 );
xor ( n13009 , n13008 , n13006 );
and ( n13010 , n13009 , n6474 );
or ( n13011 , n13007 , n13010 );
xor ( n13012 , n13004 , n13011 );
buf ( n13013 , n6235 );
xor ( n13014 , n13012 , n13013 );
buf ( n13015 , n6236 );
xor ( n13016 , n13014 , n13015 );
buf ( n13017 , n6237 );
xor ( n13018 , n13016 , n13017 );
xor ( n13019 , n12997 , n13018 );
xor ( n13020 , n13019 , n10394 );
xor ( n13021 , n10260 , n7006 );
xor ( n13022 , n13021 , n10439 );
not ( n13023 , n13022 );
buf ( n13024 , n6238 );
xor ( n13025 , n13024 , n6827 );
xor ( n13026 , n13025 , n11981 );
and ( n13027 , n13023 , n13026 );
xor ( n13028 , n13020 , n13027 );
xor ( n13029 , n12996 , n13028 );
xor ( n13030 , n9727 , n10574 );
xor ( n13031 , n13030 , n10595 );
not ( n13032 , n6474 );
buf ( n13033 , n6239 );
and ( n13034 , n13032 , n13033 );
buf ( n13035 , n6240 );
xor ( n13036 , n13035 , n13033 );
and ( n13037 , n13036 , n6474 );
or ( n13038 , n13034 , n13037 );
not ( n13039 , n6474 );
buf ( n13040 , n6241 );
and ( n13041 , n13039 , n13040 );
buf ( n13042 , n6242 );
xor ( n13043 , n13042 , n13040 );
and ( n13044 , n13043 , n6474 );
or ( n13045 , n13041 , n13044 );
xor ( n13046 , n13038 , n13045 );
buf ( n13047 , n6243 );
xor ( n13048 , n13046 , n13047 );
buf ( n13049 , n6244 );
xor ( n13050 , n13048 , n13049 );
buf ( n13051 , n6245 );
xor ( n13052 , n13050 , n13051 );
xor ( n13053 , n12449 , n13052 );
xor ( n13054 , n13053 , n10376 );
not ( n13055 , n13054 );
xor ( n13056 , n7731 , n8865 );
xor ( n13057 , n13056 , n7253 );
and ( n13058 , n13055 , n13057 );
xor ( n13059 , n13031 , n13058 );
xor ( n13060 , n13029 , n13059 );
xor ( n13061 , n11922 , n9511 );
xor ( n13062 , n13061 , n12530 );
xor ( n13063 , n9578 , n8204 );
xor ( n13064 , n13063 , n12854 );
not ( n13065 , n13064 );
buf ( n13066 , n6246 );
xor ( n13067 , n13066 , n6939 );
xor ( n13068 , n13067 , n6961 );
and ( n13069 , n13065 , n13068 );
xor ( n13070 , n13062 , n13069 );
xor ( n13071 , n13060 , n13070 );
xor ( n13072 , n12967 , n13071 );
xor ( n13073 , n10928 , n9794 );
xor ( n13074 , n13073 , n9816 );
xor ( n13075 , n6858 , n10504 );
not ( n13076 , n6474 );
buf ( n13077 , n6247 );
and ( n13078 , n13076 , n13077 );
buf ( n13079 , n6248 );
xor ( n13080 , n13079 , n13077 );
and ( n13081 , n13080 , n6474 );
or ( n13082 , n13078 , n13081 );
not ( n13083 , n6474 );
buf ( n13084 , n6249 );
and ( n13085 , n13083 , n13084 );
buf ( n13086 , n6250 );
xor ( n13087 , n13086 , n13084 );
and ( n13088 , n13087 , n6474 );
or ( n13089 , n13085 , n13088 );
xor ( n13090 , n13082 , n13089 );
xor ( n13091 , n13090 , n6918 );
buf ( n13092 , n6251 );
xor ( n13093 , n13091 , n13092 );
xor ( n13094 , n13093 , n13066 );
xor ( n13095 , n13075 , n13094 );
not ( n13096 , n13095 );
xor ( n13097 , n7762 , n12365 );
xor ( n13098 , n13097 , n12490 );
and ( n13099 , n13096 , n13098 );
xor ( n13100 , n13074 , n13099 );
xor ( n13101 , n10129 , n12213 );
xor ( n13102 , n13101 , n10768 );
xor ( n13103 , n8455 , n10193 );
xor ( n13104 , n13103 , n10209 );
not ( n13105 , n13104 );
xor ( n13106 , n8631 , n12945 );
xor ( n13107 , n13106 , n12871 );
and ( n13108 , n13105 , n13107 );
xor ( n13109 , n13102 , n13108 );
xor ( n13110 , n13100 , n13109 );
xor ( n13111 , n11656 , n11405 );
xor ( n13112 , n13111 , n11427 );
xor ( n13113 , n13082 , n6939 );
xor ( n13114 , n13113 , n6961 );
not ( n13115 , n13114 );
xor ( n13116 , n11456 , n6984 );
xor ( n13117 , n13116 , n7006 );
and ( n13118 , n13115 , n13117 );
xor ( n13119 , n13112 , n13118 );
xor ( n13120 , n13110 , n13119 );
xor ( n13121 , n10863 , n9534 );
xor ( n13122 , n13121 , n9543 );
not ( n13123 , n6474 );
buf ( n13124 , n6252 );
and ( n13125 , n13123 , n13124 );
buf ( n13126 , n6253 );
xor ( n13127 , n13126 , n13124 );
and ( n13128 , n13127 , n6474 );
or ( n13129 , n13125 , n13128 );
xor ( n13130 , n12963 , n13129 );
buf ( n13131 , n6254 );
xor ( n13132 , n13130 , n13131 );
xor ( n13133 , n13132 , n9877 );
buf ( n13134 , n6255 );
xor ( n13135 , n13133 , n13134 );
xor ( n13136 , n12540 , n13135 );
xor ( n13137 , n13136 , n8034 );
not ( n13138 , n13137 );
xor ( n13139 , n6710 , n10350 );
xor ( n13140 , n13139 , n9489 );
and ( n13141 , n13138 , n13140 );
xor ( n13142 , n13122 , n13141 );
xor ( n13143 , n13120 , n13142 );
xor ( n13144 , n8113 , n11879 );
xor ( n13145 , n13144 , n11512 );
xor ( n13146 , n11181 , n7494 );
xor ( n13147 , n13146 , n6850 );
not ( n13148 , n13147 );
xor ( n13149 , n7725 , n8865 );
xor ( n13150 , n13149 , n7253 );
and ( n13151 , n13148 , n13150 );
xor ( n13152 , n13145 , n13151 );
xor ( n13153 , n13143 , n13152 );
xor ( n13154 , n13072 , n13153 );
not ( n13155 , n13154 );
not ( n13156 , n8160 );
xor ( n13157 , n10303 , n7309 );
xor ( n13158 , n13157 , n7331 );
and ( n13159 , n13156 , n13158 );
xor ( n13160 , n8115 , n13159 );
xor ( n13161 , n13160 , n8392 );
xor ( n13162 , n13161 , n8768 );
and ( n13163 , n13155 , n13162 );
xor ( n13164 , n12951 , n13163 );
and ( n13165 , n13164 , n6475 );
or ( n13166 , n12930 , n13165 );
and ( n13167 , n12928 , n13166 );
buf ( n13168 , n13167 );
buf ( n13169 , n13168 );
not ( n13170 , n6469 );
not ( n13171 , n6475 );
and ( n13172 , n13171 , n9198 );
xor ( n13173 , n8837 , n6739 );
xor ( n13174 , n13173 , n11927 );
xor ( n13175 , n8635 , n12945 );
xor ( n13176 , n13175 , n12871 );
not ( n13177 , n13176 );
buf ( n13178 , n6256 );
xor ( n13179 , n13178 , n8935 );
xor ( n13180 , n13179 , n8950 );
and ( n13181 , n13177 , n13180 );
xor ( n13182 , n13174 , n13181 );
xor ( n13183 , n6599 , n8076 );
xor ( n13184 , n13183 , n12190 );
xor ( n13185 , n8860 , n10963 );
xor ( n13186 , n13185 , n10864 );
not ( n13187 , n13186 );
buf ( n13188 , n6257 );
xor ( n13189 , n13188 , n9217 );
xor ( n13190 , n13189 , n9417 );
and ( n13191 , n13187 , n13190 );
xor ( n13192 , n13184 , n13191 );
xor ( n13193 , n7105 , n12581 );
xor ( n13194 , n13193 , n12281 );
xor ( n13195 , n9811 , n12467 );
not ( n13196 , n6474 );
buf ( n13197 , n6258 );
and ( n13198 , n13196 , n13197 );
buf ( n13199 , n6259 );
xor ( n13200 , n13199 , n13197 );
and ( n13201 , n13200 , n6474 );
or ( n13202 , n13198 , n13201 );
not ( n13203 , n6474 );
buf ( n13204 , n6260 );
and ( n13205 , n13203 , n13204 );
buf ( n13206 , n6261 );
xor ( n13207 , n13206 , n13204 );
and ( n13208 , n13207 , n6474 );
or ( n13209 , n13205 , n13208 );
xor ( n13210 , n13202 , n13209 );
xor ( n13211 , n13210 , n10046 );
buf ( n13212 , n6262 );
xor ( n13213 , n13211 , n13212 );
buf ( n13214 , n6263 );
xor ( n13215 , n13213 , n13214 );
xor ( n13216 , n13195 , n13215 );
not ( n13217 , n13216 );
xor ( n13218 , n7272 , n7159 );
xor ( n13219 , n13218 , n7181 );
and ( n13220 , n13217 , n13219 );
xor ( n13221 , n13194 , n13220 );
xor ( n13222 , n13192 , n13221 );
not ( n13223 , n6474 );
buf ( n13224 , n6264 );
and ( n13225 , n13223 , n13224 );
buf ( n13226 , n6265 );
xor ( n13227 , n13226 , n13224 );
and ( n13228 , n13227 , n6474 );
or ( n13229 , n13225 , n13228 );
xor ( n13230 , n13229 , n11981 );
xor ( n13231 , n13230 , n7566 );
not ( n13232 , n13174 );
and ( n13233 , n13232 , n13176 );
xor ( n13234 , n13231 , n13233 );
xor ( n13235 , n13222 , n13234 );
xor ( n13236 , n8130 , n7046 );
xor ( n13237 , n13236 , n8414 );
xor ( n13238 , n10460 , n10246 );
xor ( n13239 , n13238 , n11252 );
not ( n13240 , n13239 );
xor ( n13241 , n9893 , n8447 );
xor ( n13242 , n13241 , n8469 );
and ( n13243 , n13240 , n13242 );
xor ( n13244 , n13237 , n13243 );
xor ( n13245 , n13235 , n13244 );
xor ( n13246 , n7854 , n11512 );
xor ( n13247 , n13246 , n11520 );
xor ( n13248 , n8530 , n9378 );
xor ( n13249 , n13248 , n9400 );
not ( n13250 , n13249 );
buf ( n13251 , n6266 );
xor ( n13252 , n13251 , n9354 );
xor ( n13253 , n13252 , n7710 );
and ( n13254 , n13250 , n13253 );
xor ( n13255 , n13247 , n13254 );
xor ( n13256 , n13245 , n13255 );
xor ( n13257 , n13182 , n13256 );
xor ( n13258 , n10524 , n12302 );
not ( n13259 , n6474 );
buf ( n13260 , n6267 );
and ( n13261 , n13259 , n13260 );
buf ( n13262 , n6268 );
xor ( n13263 , n13262 , n13260 );
and ( n13264 , n13263 , n6474 );
or ( n13265 , n13261 , n13264 );
buf ( n13266 , n6269 );
xor ( n13267 , n13265 , n13266 );
buf ( n13268 , n6270 );
xor ( n13269 , n13267 , n13268 );
buf ( n13270 , n6271 );
xor ( n13271 , n13269 , n13270 );
buf ( n13272 , n6272 );
xor ( n13273 , n13271 , n13272 );
xor ( n13274 , n13258 , n13273 );
xor ( n13275 , n12547 , n13135 );
xor ( n13276 , n13275 , n8034 );
not ( n13277 , n13276 );
xor ( n13278 , n7407 , n6516 );
xor ( n13279 , n13278 , n13052 );
and ( n13280 , n13277 , n13279 );
xor ( n13281 , n13274 , n13280 );
buf ( n13282 , n6273 );
xor ( n13283 , n13282 , n7659 );
xor ( n13284 , n13283 , n7681 );
xor ( n13285 , n10594 , n6913 );
xor ( n13286 , n13285 , n8600 );
not ( n13287 , n13286 );
xor ( n13288 , n11591 , n10990 );
xor ( n13289 , n13288 , n10022 );
and ( n13290 , n13287 , n13289 );
xor ( n13291 , n13284 , n13290 );
xor ( n13292 , n13281 , n13291 );
xor ( n13293 , n7373 , n10224 );
xor ( n13294 , n13293 , n10246 );
xor ( n13295 , n7094 , n12822 );
not ( n13296 , n6474 );
buf ( n13297 , n6274 );
and ( n13298 , n13296 , n13297 );
buf ( n13299 , n6275 );
xor ( n13300 , n13299 , n13297 );
and ( n13301 , n13300 , n6474 );
or ( n13302 , n13298 , n13301 );
not ( n13303 , n6474 );
buf ( n13304 , n6276 );
and ( n13305 , n13303 , n13304 );
buf ( n13306 , n6277 );
xor ( n13307 , n13306 , n13304 );
and ( n13308 , n13307 , n6474 );
or ( n13309 , n13305 , n13308 );
xor ( n13310 , n13302 , n13309 );
buf ( n13311 , n6278 );
xor ( n13312 , n13310 , n13311 );
buf ( n13313 , n6279 );
xor ( n13314 , n13312 , n13313 );
xor ( n13315 , n13314 , n9175 );
xor ( n13316 , n13295 , n13315 );
not ( n13317 , n13316 );
xor ( n13318 , n13038 , n12987 );
not ( n13319 , n6474 );
buf ( n13320 , n6280 );
and ( n13321 , n13319 , n13320 );
buf ( n13322 , n6281 );
xor ( n13323 , n13322 , n13320 );
and ( n13324 , n13323 , n6474 );
or ( n13325 , n13321 , n13324 );
not ( n13326 , n6474 );
buf ( n13327 , n6282 );
and ( n13328 , n13326 , n13327 );
buf ( n13329 , n6283 );
xor ( n13330 , n13329 , n13327 );
and ( n13331 , n13330 , n6474 );
or ( n13332 , n13328 , n13331 );
xor ( n13333 , n13325 , n13332 );
buf ( n13334 , n6284 );
xor ( n13335 , n13333 , n13334 );
buf ( n13336 , n6285 );
xor ( n13337 , n13335 , n13336 );
buf ( n13338 , n6286 );
xor ( n13339 , n13337 , n13338 );
xor ( n13340 , n13318 , n13339 );
and ( n13341 , n13317 , n13340 );
xor ( n13342 , n13294 , n13341 );
xor ( n13343 , n13292 , n13342 );
xor ( n13344 , n10190 , n9238 );
xor ( n13345 , n13344 , n9260 );
xor ( n13346 , n6537 , n10731 );
xor ( n13347 , n13346 , n10745 );
not ( n13348 , n13347 );
xor ( n13349 , n8196 , n11146 );
xor ( n13350 , n13349 , n9651 );
and ( n13351 , n13348 , n13350 );
xor ( n13352 , n13345 , n13351 );
xor ( n13353 , n13343 , n13352 );
buf ( n13354 , n6287 );
not ( n13355 , n6474 );
buf ( n13356 , n6288 );
and ( n13357 , n13355 , n13356 );
buf ( n13358 , n6289 );
xor ( n13359 , n13358 , n13356 );
and ( n13360 , n13359 , n6474 );
or ( n13361 , n13357 , n13360 );
buf ( n13362 , n6290 );
xor ( n13363 , n13361 , n13362 );
buf ( n13364 , n6291 );
xor ( n13365 , n13363 , n13364 );
xor ( n13366 , n13365 , n12147 );
xor ( n13367 , n13366 , n12831 );
xor ( n13368 , n13354 , n13367 );
xor ( n13369 , n13368 , n10963 );
xor ( n13370 , n11554 , n9816 );
xor ( n13371 , n13370 , n6811 );
not ( n13372 , n13371 );
xor ( n13373 , n7808 , n7463 );
xor ( n13374 , n13373 , n7399 );
and ( n13375 , n13372 , n13374 );
xor ( n13376 , n13369 , n13375 );
xor ( n13377 , n13353 , n13376 );
xor ( n13378 , n13257 , n13377 );
xor ( n13379 , n10728 , n10625 );
xor ( n13380 , n13379 , n7208 );
not ( n13381 , n6474 );
buf ( n13382 , n6292 );
and ( n13383 , n13381 , n13382 );
buf ( n13384 , n6293 );
xor ( n13385 , n13384 , n13382 );
and ( n13386 , n13385 , n6474 );
or ( n13387 , n13383 , n13386 );
xor ( n13388 , n8675 , n13387 );
buf ( n13389 , n6294 );
xor ( n13390 , n13388 , n13389 );
xor ( n13391 , n13390 , n9676 );
xor ( n13392 , n13391 , n10912 );
xor ( n13393 , n8387 , n13392 );
xor ( n13394 , n13393 , n7994 );
not ( n13395 , n13394 );
xor ( n13396 , n6819 , n11636 );
xor ( n13397 , n13396 , n11657 );
and ( n13398 , n13395 , n13397 );
xor ( n13399 , n13380 , n13398 );
xor ( n13400 , n9212 , n7134 );
xor ( n13401 , n13400 , n10527 );
xor ( n13402 , n8597 , n7822 );
xor ( n13403 , n13402 , n7837 );
not ( n13404 , n13403 );
xor ( n13405 , n11519 , n8495 );
xor ( n13406 , n13405 , n8517 );
and ( n13407 , n13404 , n13406 );
xor ( n13408 , n13401 , n13407 );
xor ( n13409 , n7153 , n9543 );
not ( n13410 , n6474 );
buf ( n13411 , n6295 );
and ( n13412 , n13410 , n13411 );
buf ( n13413 , n6296 );
xor ( n13414 , n13413 , n13411 );
and ( n13415 , n13414 , n6474 );
or ( n13416 , n13412 , n13415 );
not ( n13417 , n6474 );
buf ( n13418 , n6297 );
and ( n13419 , n13417 , n13418 );
buf ( n13420 , n6298 );
xor ( n13421 , n13420 , n13418 );
and ( n13422 , n13421 , n6474 );
or ( n13423 , n13419 , n13422 );
xor ( n13424 , n13416 , n13423 );
xor ( n13425 , n13424 , n8663 );
xor ( n13426 , n13425 , n13282 );
xor ( n13427 , n13426 , n7639 );
xor ( n13428 , n13409 , n13427 );
xor ( n13429 , n9436 , n10549 );
xor ( n13430 , n13429 , n12024 );
not ( n13431 , n13430 );
xor ( n13432 , n9871 , n11693 );
xor ( n13433 , n13432 , n11714 );
and ( n13434 , n13431 , n13433 );
xor ( n13435 , n13428 , n13434 );
xor ( n13436 , n13408 , n13435 );
xor ( n13437 , n10371 , n13339 );
xor ( n13438 , n13437 , n12649 );
xor ( n13439 , n10143 , n10768 );
xor ( n13440 , n13439 , n10790 );
not ( n13441 , n13440 );
xor ( n13442 , n10438 , n9710 );
xor ( n13443 , n13442 , n9732 );
and ( n13444 , n13441 , n13443 );
xor ( n13445 , n13438 , n13444 );
xor ( n13446 , n13436 , n13445 );
xor ( n13447 , n11900 , n6872 );
not ( n13448 , n6474 );
buf ( n13449 , n6299 );
and ( n13450 , n13448 , n13449 );
buf ( n13451 , n6300 );
xor ( n13452 , n13451 , n13449 );
and ( n13453 , n13452 , n6474 );
or ( n13454 , n13450 , n13453 );
not ( n13455 , n6474 );
buf ( n13456 , n6301 );
and ( n13457 , n13455 , n13456 );
buf ( n13458 , n6302 );
xor ( n13459 , n13458 , n13456 );
and ( n13460 , n13459 , n6474 );
or ( n13461 , n13457 , n13460 );
xor ( n13462 , n13454 , n13461 );
buf ( n13463 , n6303 );
xor ( n13464 , n13462 , n13463 );
buf ( n13465 , n6304 );
xor ( n13466 , n13464 , n13465 );
buf ( n13467 , n6305 );
xor ( n13468 , n13466 , n13467 );
xor ( n13469 , n13447 , n13468 );
not ( n13470 , n13380 );
and ( n13471 , n13470 , n13394 );
xor ( n13472 , n13469 , n13471 );
xor ( n13473 , n13446 , n13472 );
xor ( n13474 , n10204 , n9260 );
not ( n13475 , n6474 );
buf ( n13476 , n6306 );
and ( n13477 , n13475 , n13476 );
buf ( n13478 , n6307 );
xor ( n13479 , n13478 , n13476 );
and ( n13480 , n13479 , n6474 );
or ( n13481 , n13477 , n13480 );
xor ( n13482 , n8921 , n13481 );
buf ( n13483 , n6308 );
xor ( n13484 , n13482 , n13483 );
buf ( n13485 , n6309 );
xor ( n13486 , n13484 , n13485 );
xor ( n13487 , n13486 , n13178 );
xor ( n13488 , n13474 , n13487 );
xor ( n13489 , n7092 , n12822 );
xor ( n13490 , n13489 , n13315 );
not ( n13491 , n13490 );
xor ( n13492 , n6605 , n8076 );
xor ( n13493 , n13492 , n12190 );
and ( n13494 , n13491 , n13493 );
xor ( n13495 , n13488 , n13494 );
xor ( n13496 , n13473 , n13495 );
xor ( n13497 , n13399 , n13496 );
not ( n13498 , n6607 );
xor ( n13499 , n9432 , n10549 );
xor ( n13500 , n13499 , n12024 );
and ( n13501 , n13498 , n13500 );
xor ( n13502 , n6561 , n13501 );
not ( n13503 , n6474 );
buf ( n13504 , n6310 );
and ( n13505 , n13503 , n13504 );
buf ( n13506 , n6311 );
xor ( n13507 , n13506 , n13504 );
and ( n13508 , n13507 , n6474 );
or ( n13509 , n13505 , n13508 );
not ( n13510 , n6474 );
buf ( n13511 , n6312 );
and ( n13512 , n13510 , n13511 );
buf ( n13513 , n6313 );
xor ( n13514 , n13513 , n13511 );
and ( n13515 , n13514 , n6474 );
or ( n13516 , n13512 , n13515 );
xor ( n13517 , n13509 , n13516 );
buf ( n13518 , n6314 );
xor ( n13519 , n13517 , n13518 );
buf ( n13520 , n6315 );
xor ( n13521 , n13519 , n13520 );
buf ( n13522 , n6316 );
xor ( n13523 , n13521 , n13522 );
xor ( n13524 , n7552 , n13523 );
xor ( n13525 , n13524 , n8638 );
not ( n13526 , n13525 );
xor ( n13527 , n12788 , n8600 );
xor ( n13528 , n13527 , n8622 );
and ( n13529 , n13526 , n13528 );
xor ( n13530 , n6786 , n13529 );
xor ( n13531 , n13502 , n13530 );
xor ( n13532 , n6592 , n8076 );
xor ( n13533 , n13532 , n12190 );
not ( n13534 , n13533 );
xor ( n13535 , n10123 , n12213 );
xor ( n13536 , n13535 , n10768 );
and ( n13537 , n13534 , n13536 );
xor ( n13538 , n6914 , n13537 );
xor ( n13539 , n13531 , n13538 );
not ( n13540 , n6474 );
buf ( n13541 , n6317 );
and ( n13542 , n13540 , n13541 );
buf ( n13543 , n6318 );
xor ( n13544 , n13543 , n13541 );
and ( n13545 , n13544 , n6474 );
or ( n13546 , n13542 , n13545 );
not ( n13547 , n6474 );
buf ( n13548 , n6319 );
and ( n13549 , n13547 , n13548 );
buf ( n13550 , n6320 );
xor ( n13551 , n13550 , n13548 );
and ( n13552 , n13551 , n6474 );
or ( n13553 , n13549 , n13552 );
xor ( n13554 , n13546 , n13553 );
buf ( n13555 , n6321 );
xor ( n13556 , n13554 , n13555 );
buf ( n13557 , n6322 );
xor ( n13558 , n13556 , n13557 );
buf ( n13559 , n6323 );
xor ( n13560 , n13558 , n13559 );
xor ( n13561 , n11397 , n13560 );
xor ( n13562 , n13561 , n12699 );
not ( n13563 , n13562 );
xor ( n13564 , n9935 , n12548 );
xor ( n13565 , n13564 , n9238 );
and ( n13566 , n13563 , n13565 );
xor ( n13567 , n7047 , n13566 );
xor ( n13568 , n13539 , n13567 );
xor ( n13569 , n10296 , n7309 );
xor ( n13570 , n13569 , n7331 );
not ( n13571 , n13570 );
xor ( n13572 , n8381 , n13392 );
xor ( n13573 , n13572 , n7994 );
and ( n13574 , n13571 , n13573 );
xor ( n13575 , n7182 , n13574 );
xor ( n13576 , n13568 , n13575 );
xor ( n13577 , n13497 , n13576 );
not ( n13578 , n13577 );
not ( n13579 , n8389 );
not ( n13580 , n6474 );
buf ( n13581 , n6324 );
and ( n13582 , n13580 , n13581 );
buf ( n13583 , n6325 );
xor ( n13584 , n13583 , n13581 );
and ( n13585 , n13584 , n6474 );
or ( n13586 , n13582 , n13585 );
xor ( n13587 , n12914 , n13586 );
buf ( n13588 , n6326 );
xor ( n13589 , n13587 , n13588 );
xor ( n13590 , n13589 , n12305 );
xor ( n13591 , n13590 , n11254 );
xor ( n13592 , n9504 , n13591 );
not ( n13593 , n6474 );
buf ( n13594 , n6327 );
and ( n13595 , n13593 , n13594 );
buf ( n13596 , n6328 );
xor ( n13597 , n13596 , n13594 );
and ( n13598 , n13597 , n6474 );
or ( n13599 , n13595 , n13598 );
buf ( n13600 , n6329 );
xor ( n13601 , n13599 , n13600 );
buf ( n13602 , n6330 );
xor ( n13603 , n13601 , n13602 );
xor ( n13604 , n13603 , n9546 );
buf ( n13605 , n6331 );
xor ( n13606 , n13604 , n13605 );
xor ( n13607 , n13592 , n13606 );
and ( n13608 , n13579 , n13607 );
xor ( n13609 , n8337 , n13608 );
xor ( n13610 , n13609 , n8392 );
xor ( n13611 , n13610 , n8768 );
and ( n13612 , n13578 , n13611 );
xor ( n13613 , n13378 , n13612 );
and ( n13614 , n13613 , n6475 );
or ( n13615 , n13172 , n13614 );
and ( n13616 , n13170 , n13615 );
buf ( n13617 , n13616 );
buf ( n13618 , n13617 );
not ( n13619 , n6469 );
not ( n13620 , n6475 );
and ( n13621 , n13620 , n7091 );
xor ( n13622 , n9709 , n11949 );
xor ( n13623 , n13622 , n10574 );
xor ( n13624 , n7646 , n6673 );
xor ( n13625 , n13624 , n6695 );
not ( n13626 , n13625 );
not ( n13627 , n6474 );
buf ( n13628 , n6332 );
and ( n13629 , n13627 , n13628 );
buf ( n13630 , n6333 );
xor ( n13631 , n13630 , n13628 );
and ( n13632 , n13631 , n6474 );
or ( n13633 , n13629 , n13632 );
not ( n13634 , n6474 );
buf ( n13635 , n6334 );
and ( n13636 , n13634 , n13635 );
buf ( n13637 , n6335 );
xor ( n13638 , n13637 , n13635 );
and ( n13639 , n13638 , n6474 );
or ( n13640 , n13636 , n13639 );
xor ( n13641 , n13633 , n13640 );
buf ( n13642 , n6336 );
xor ( n13643 , n13641 , n13642 );
buf ( n13644 , n6337 );
xor ( n13645 , n13643 , n13644 );
buf ( n13646 , n6338 );
xor ( n13647 , n13645 , n13646 );
xor ( n13648 , n11268 , n13647 );
xor ( n13649 , n13648 , n8188 );
and ( n13650 , n13626 , n13649 );
xor ( n13651 , n13623 , n13650 );
xor ( n13652 , n10373 , n13339 );
xor ( n13653 , n13652 , n12649 );
not ( n13654 , n13623 );
and ( n13655 , n13654 , n13625 );
xor ( n13656 , n13653 , n13655 );
xor ( n13657 , n11129 , n12530 );
xor ( n13658 , n13657 , n10697 );
xor ( n13659 , n8864 , n10963 );
xor ( n13660 , n13659 , n10864 );
not ( n13661 , n13660 );
xor ( n13662 , n10099 , n9079 );
xor ( n13663 , n13662 , n9094 );
and ( n13664 , n13661 , n13663 );
xor ( n13665 , n13658 , n13664 );
xor ( n13666 , n13656 , n13665 );
xor ( n13667 , n9145 , n12097 );
xor ( n13668 , n13667 , n12111 );
xor ( n13669 , n8621 , n7837 );
not ( n13670 , n6474 );
buf ( n13671 , n6339 );
and ( n13672 , n13670 , n13671 );
buf ( n13673 , n6340 );
xor ( n13674 , n13673 , n13671 );
and ( n13675 , n13674 , n6474 );
or ( n13676 , n13672 , n13675 );
not ( n13677 , n6474 );
buf ( n13678 , n6341 );
and ( n13679 , n13677 , n13678 );
buf ( n13680 , n6342 );
xor ( n13681 , n13680 , n13678 );
and ( n13682 , n13681 , n6474 );
or ( n13683 , n13679 , n13682 );
xor ( n13684 , n13676 , n13683 );
buf ( n13685 , n6343 );
xor ( n13686 , n13684 , n13685 );
buf ( n13687 , n6344 );
xor ( n13688 , n13686 , n13687 );
buf ( n13689 , n6345 );
xor ( n13690 , n13688 , n13689 );
xor ( n13691 , n13669 , n13690 );
not ( n13692 , n13691 );
not ( n13693 , n6474 );
buf ( n13694 , n6346 );
and ( n13695 , n13693 , n13694 );
buf ( n13696 , n6347 );
xor ( n13697 , n13696 , n13694 );
and ( n13698 , n13697 , n6474 );
or ( n13699 , n13695 , n13698 );
xor ( n13700 , n13699 , n12258 );
buf ( n13701 , n6348 );
xor ( n13702 , n13700 , n13701 );
buf ( n13703 , n6349 );
xor ( n13704 , n13702 , n13703 );
xor ( n13705 , n13704 , n11307 );
xor ( n13706 , n6681 , n13705 );
xor ( n13707 , n13706 , n12727 );
and ( n13708 , n13692 , n13707 );
xor ( n13709 , n13668 , n13708 );
xor ( n13710 , n13666 , n13709 );
xor ( n13711 , n8571 , n9732 );
xor ( n13712 , n13711 , n8227 );
xor ( n13713 , n9025 , n8336 );
xor ( n13714 , n13713 , n8535 );
not ( n13715 , n13714 );
xor ( n13716 , n7368 , n10224 );
xor ( n13717 , n13716 , n10246 );
and ( n13718 , n13715 , n13717 );
xor ( n13719 , n13712 , n13718 );
xor ( n13720 , n13710 , n13719 );
xor ( n13721 , n10546 , n13273 );
xor ( n13722 , n13721 , n8820 );
xor ( n13723 , n11328 , n11763 );
xor ( n13724 , n13723 , n10130 );
not ( n13725 , n13724 );
xor ( n13726 , n9520 , n6606 );
xor ( n13727 , n13726 , n9123 );
and ( n13728 , n13725 , n13727 );
xor ( n13729 , n13722 , n13728 );
xor ( n13730 , n13720 , n13729 );
xor ( n13731 , n13651 , n13730 );
xor ( n13732 , n13699 , n9002 );
xor ( n13733 , n13732 , n11329 );
xor ( n13734 , n11125 , n12530 );
xor ( n13735 , n13734 , n10697 );
not ( n13736 , n13735 );
xor ( n13737 , n13588 , n11275 );
xor ( n13738 , n13737 , n9559 );
and ( n13739 , n13736 , n13738 );
xor ( n13740 , n13733 , n13739 );
xor ( n13741 , n8729 , n11252 );
xor ( n13742 , n13741 , n8269 );
xor ( n13743 , n12461 , n10376 );
xor ( n13744 , n13743 , n10067 );
not ( n13745 , n13744 );
xor ( n13746 , n7965 , n10146 );
xor ( n13747 , n13746 , n10652 );
and ( n13748 , n13745 , n13747 );
xor ( n13749 , n13742 , n13748 );
xor ( n13750 , n13740 , n13749 );
xor ( n13751 , n11315 , n11763 );
xor ( n13752 , n13751 , n10130 );
xor ( n13753 , n13461 , n13094 );
xor ( n13754 , n13753 , n12097 );
not ( n13755 , n13754 );
xor ( n13756 , n12940 , n7360 );
xor ( n13757 , n13756 , n7376 );
and ( n13758 , n13755 , n13757 );
xor ( n13759 , n13752 , n13758 );
xor ( n13760 , n13750 , n13759 );
xor ( n13761 , n9298 , n10105 );
not ( n13762 , n6474 );
buf ( n13763 , n6350 );
and ( n13764 , n13762 , n13763 );
buf ( n13765 , n6351 );
xor ( n13766 , n13765 , n13763 );
and ( n13767 , n13766 , n6474 );
or ( n13768 , n13764 , n13767 );
xor ( n13769 , n12316 , n13768 );
buf ( n13770 , n6352 );
xor ( n13771 , n13769 , n13770 );
xor ( n13772 , n13771 , n12224 );
buf ( n13773 , n6353 );
xor ( n13774 , n13772 , n13773 );
xor ( n13775 , n13761 , n13774 );
xor ( n13776 , n7087 , n12822 );
xor ( n13777 , n13776 , n13315 );
not ( n13778 , n13777 );
xor ( n13779 , n10620 , n8517 );
xor ( n13780 , n13779 , n11462 );
and ( n13781 , n13778 , n13780 );
xor ( n13782 , n13775 , n13781 );
xor ( n13783 , n13760 , n13782 );
xor ( n13784 , n12176 , n7274 );
not ( n13785 , n6474 );
buf ( n13786 , n6354 );
and ( n13787 , n13785 , n13786 );
buf ( n13788 , n6355 );
xor ( n13789 , n13788 , n13786 );
and ( n13790 , n13789 , n6474 );
or ( n13791 , n13787 , n13790 );
xor ( n13792 , n8986 , n13791 );
buf ( n13793 , n6356 );
xor ( n13794 , n13792 , n13793 );
buf ( n13795 , n6357 );
xor ( n13796 , n13794 , n13795 );
buf ( n13797 , n6358 );
xor ( n13798 , n13796 , n13797 );
xor ( n13799 , n13784 , n13798 );
xor ( n13800 , n9019 , n8336 );
xor ( n13801 , n13800 , n8535 );
not ( n13802 , n13801 );
xor ( n13803 , n9412 , n10527 );
xor ( n13804 , n13803 , n10549 );
and ( n13805 , n13802 , n13804 );
xor ( n13806 , n13799 , n13805 );
xor ( n13807 , n13783 , n13806 );
xor ( n13808 , n13731 , n13807 );
not ( n13809 , n6474 );
buf ( n13810 , n6359 );
and ( n13811 , n13809 , n13810 );
buf ( n13812 , n6360 );
xor ( n13813 , n13812 , n13810 );
and ( n13814 , n13813 , n6474 );
or ( n13815 , n13811 , n13814 );
xor ( n13816 , n13815 , n9770 );
xor ( n13817 , n13816 , n7112 );
xor ( n13818 , n9088 , n8743 );
xor ( n13819 , n13818 , n8764 );
not ( n13820 , n13819 );
xor ( n13821 , n6555 , n10745 );
not ( n13822 , n6474 );
buf ( n13823 , n6361 );
and ( n13824 , n13822 , n13823 );
buf ( n13825 , n6362 );
xor ( n13826 , n13825 , n13823 );
and ( n13827 , n13826 , n6474 );
or ( n13828 , n13824 , n13827 );
not ( n13829 , n6474 );
buf ( n13830 , n6363 );
and ( n13831 , n13829 , n13830 );
buf ( n13832 , n6364 );
xor ( n13833 , n13832 , n13830 );
and ( n13834 , n13833 , n6474 );
or ( n13835 , n13831 , n13834 );
xor ( n13836 , n13828 , n13835 );
buf ( n13837 , n6365 );
xor ( n13838 , n13836 , n13837 );
buf ( n13839 , n6366 );
xor ( n13840 , n13838 , n13839 );
buf ( n13841 , n6367 );
xor ( n13842 , n13840 , n13841 );
xor ( n13843 , n13821 , n13842 );
and ( n13844 , n13820 , n13843 );
xor ( n13845 , n13817 , n13844 );
xor ( n13846 , n6826 , n11636 );
xor ( n13847 , n13846 , n11657 );
xor ( n13848 , n12105 , n9606 );
xor ( n13849 , n13848 , n9628 );
not ( n13850 , n13849 );
xor ( n13851 , n11024 , n11998 );
xor ( n13852 , n13851 , n7521 );
and ( n13853 , n13850 , n13852 );
xor ( n13854 , n13847 , n13853 );
xor ( n13855 , n12778 , n11905 );
xor ( n13856 , n13855 , n11865 );
not ( n13857 , n13817 );
and ( n13858 , n13857 , n13819 );
xor ( n13859 , n13856 , n13858 );
xor ( n13860 , n13854 , n13859 );
xor ( n13861 , n12870 , n7376 );
xor ( n13862 , n13861 , n10465 );
xor ( n13863 , n9614 , n7883 );
xor ( n13864 , n13863 , n10731 );
not ( n13865 , n13864 );
xor ( n13866 , n8567 , n9732 );
xor ( n13867 , n13866 , n8227 );
and ( n13868 , n13865 , n13867 );
xor ( n13869 , n13862 , n13868 );
xor ( n13870 , n13860 , n13869 );
xor ( n13871 , n11740 , n7681 );
not ( n13872 , n6474 );
buf ( n13873 , n6368 );
and ( n13874 , n13872 , n13873 );
buf ( n13875 , n6369 );
xor ( n13876 , n13875 , n13873 );
and ( n13877 , n13876 , n6474 );
or ( n13878 , n13874 , n13877 );
buf ( n13879 , n6370 );
xor ( n13880 , n13878 , n13879 );
buf ( n13881 , n6371 );
xor ( n13882 , n13880 , n13881 );
buf ( n13883 , n6372 );
xor ( n13884 , n13882 , n13883 );
buf ( n13885 , n6373 );
xor ( n13886 , n13884 , n13885 );
xor ( n13887 , n13871 , n13886 );
xor ( n13888 , n8928 , n7072 );
xor ( n13889 , n13888 , n7095 );
not ( n13890 , n13889 );
xor ( n13891 , n12523 , n13606 );
xor ( n13892 , n13891 , n11583 );
and ( n13893 , n13890 , n13892 );
xor ( n13894 , n13887 , n13893 );
xor ( n13895 , n13870 , n13894 );
xor ( n13896 , n10624 , n8517 );
xor ( n13897 , n13896 , n11462 );
xor ( n13898 , n13454 , n13094 );
xor ( n13899 , n13898 , n12097 );
not ( n13900 , n13899 );
xor ( n13901 , n13791 , n7181 );
xor ( n13902 , n13901 , n9002 );
and ( n13903 , n13900 , n13902 );
xor ( n13904 , n13897 , n13903 );
xor ( n13905 , n13895 , n13904 );
xor ( n13906 , n13845 , n13905 );
xor ( n13907 , n8009 , n8137 );
xor ( n13908 , n13907 , n8159 );
xor ( n13909 , n7025 , n11031 );
xor ( n13910 , n13909 , n11052 );
not ( n13911 , n13910 );
buf ( n13912 , n6374 );
xor ( n13913 , n13912 , n12407 );
xor ( n13914 , n13913 , n12381 );
and ( n13915 , n13911 , n13914 );
xor ( n13916 , n13908 , n13915 );
not ( n13917 , n6474 );
buf ( n13918 , n6375 );
and ( n13919 , n13917 , n13918 );
buf ( n13920 , n6376 );
xor ( n13921 , n13920 , n13918 );
and ( n13922 , n13921 , n6474 );
or ( n13923 , n13919 , n13922 );
not ( n13924 , n6474 );
buf ( n13925 , n6377 );
and ( n13926 , n13924 , n13925 );
buf ( n13927 , n6378 );
xor ( n13928 , n13927 , n13925 );
and ( n13929 , n13928 , n6474 );
or ( n13930 , n13926 , n13929 );
xor ( n13931 , n13923 , n13930 );
xor ( n13932 , n13931 , n12997 );
buf ( n13933 , n6379 );
xor ( n13934 , n13932 , n13933 );
buf ( n13935 , n6380 );
xor ( n13936 , n13934 , n13935 );
xor ( n13937 , n8262 , n13936 );
xor ( n13938 , n13937 , n11786 );
xor ( n13939 , n7225 , n10263 );
xor ( n13940 , n13939 , n10285 );
not ( n13941 , n13940 );
xor ( n13942 , n8412 , n8314 );
xor ( n13943 , n13942 , n8336 );
and ( n13944 , n13941 , n13943 );
xor ( n13945 , n13938 , n13944 );
xor ( n13946 , n13916 , n13945 );
xor ( n13947 , n10589 , n6913 );
xor ( n13948 , n13947 , n8600 );
xor ( n13949 , n9255 , n8056 );
xor ( n13950 , n13949 , n8935 );
not ( n13951 , n13950 );
xor ( n13952 , n7834 , n7399 );
xor ( n13953 , n13952 , n7421 );
and ( n13954 , n13951 , n13953 );
xor ( n13955 , n13948 , n13954 );
xor ( n13956 , n13946 , n13955 );
xor ( n13957 , n9574 , n8204 );
xor ( n13958 , n13957 , n12854 );
xor ( n13959 , n13047 , n12987 );
xor ( n13960 , n13959 , n13339 );
not ( n13961 , n13960 );
xor ( n13962 , n13520 , n11427 );
xor ( n13963 , n13962 , n12945 );
and ( n13964 , n13961 , n13963 );
xor ( n13965 , n13958 , n13964 );
xor ( n13966 , n13956 , n13965 );
xor ( n13967 , n11734 , n7681 );
xor ( n13968 , n13967 , n13886 );
buf ( n13969 , n6381 );
xor ( n13970 , n13969 , n11833 );
xor ( n13971 , n13970 , n12365 );
not ( n13972 , n13971 );
xor ( n13973 , n8910 , n11481 );
xor ( n13974 , n13973 , n8696 );
and ( n13975 , n13972 , n13974 );
xor ( n13976 , n13968 , n13975 );
xor ( n13977 , n13966 , n13976 );
xor ( n13978 , n13906 , n13977 );
not ( n13979 , n13978 );
xor ( n13980 , n7023 , n11031 );
xor ( n13981 , n13980 , n11052 );
xor ( n13982 , n12092 , n6961 );
xor ( n13983 , n13982 , n9606 );
not ( n13984 , n13983 );
and ( n13985 , n13984 , n11306 );
xor ( n13986 , n13981 , n13985 );
xor ( n13987 , n8653 , n12871 );
xor ( n13988 , n13987 , n9079 );
not ( n13989 , n13988 );
not ( n13990 , n6474 );
buf ( n13991 , n6382 );
and ( n13992 , n13990 , n13991 );
buf ( n13993 , n6383 );
xor ( n13994 , n13993 , n13991 );
and ( n13995 , n13994 , n6474 );
or ( n13996 , n13992 , n13995 );
not ( n13997 , n6474 );
buf ( n13998 , n6384 );
and ( n13999 , n13997 , n13998 );
buf ( n14000 , n6385 );
xor ( n14001 , n14000 , n13998 );
and ( n14002 , n14001 , n6474 );
or ( n14003 , n13999 , n14002 );
xor ( n14004 , n13996 , n14003 );
buf ( n14005 , n6386 );
xor ( n14006 , n14004 , n14005 );
xor ( n14007 , n14006 , n12751 );
buf ( n14008 , n6387 );
xor ( n14009 , n14007 , n14008 );
xor ( n14010 , n7355 , n14009 );
xor ( n14011 , n14010 , n10224 );
and ( n14012 , n13989 , n14011 );
xor ( n14013 , n11228 , n14012 );
xor ( n14014 , n12736 , n7948 );
xor ( n14015 , n14014 , n7970 );
not ( n14016 , n14015 );
not ( n14017 , n6474 );
buf ( n14018 , n6388 );
and ( n14019 , n14017 , n14018 );
buf ( n14020 , n6389 );
xor ( n14021 , n14020 , n14018 );
and ( n14022 , n14021 , n6474 );
or ( n14023 , n14019 , n14022 );
buf ( n14024 , n6390 );
xor ( n14025 , n14023 , n14024 );
buf ( n14026 , n6391 );
xor ( n14027 , n14025 , n14026 );
buf ( n14028 , n6392 );
xor ( n14029 , n14027 , n14028 );
xor ( n14030 , n14029 , n8870 );
xor ( n14031 , n12360 , n14030 );
xor ( n14032 , n14031 , n8366 );
and ( n14033 , n14016 , n14032 );
xor ( n14034 , n11280 , n14033 );
xor ( n14035 , n14013 , n14034 );
not ( n14036 , n13981 );
and ( n14037 , n14036 , n13983 );
xor ( n14038 , n11368 , n14037 );
xor ( n14039 , n14035 , n14038 );
xor ( n14040 , n7414 , n6516 );
xor ( n14041 , n14040 , n13052 );
not ( n14042 , n14041 );
xor ( n14043 , n11690 , n9047 );
xor ( n14044 , n14043 , n9338 );
and ( n14045 , n14042 , n14044 );
xor ( n14046 , n11386 , n14045 );
xor ( n14047 , n14039 , n14046 );
not ( n14048 , n11172 );
not ( n14049 , n6474 );
buf ( n14050 , n6393 );
and ( n14051 , n14049 , n14050 );
buf ( n14052 , n6394 );
xor ( n14053 , n14052 , n14050 );
and ( n14054 , n14053 , n6474 );
or ( n14055 , n14051 , n14054 );
not ( n14056 , n6474 );
buf ( n14057 , n6395 );
and ( n14058 , n14056 , n14057 );
buf ( n14059 , n6396 );
xor ( n14060 , n14059 , n14057 );
and ( n14061 , n14060 , n6474 );
or ( n14062 , n14058 , n14061 );
xor ( n14063 , n14055 , n14062 );
xor ( n14064 , n14063 , n6790 );
buf ( n14065 , n6397 );
xor ( n14066 , n14064 , n14065 );
xor ( n14067 , n14066 , n12615 );
xor ( n14068 , n12644 , n14067 );
not ( n14069 , n6474 );
buf ( n14070 , n6398 );
and ( n14071 , n14069 , n14070 );
buf ( n14072 , n6399 );
xor ( n14073 , n14072 , n14070 );
and ( n14074 , n14073 , n6474 );
or ( n14075 , n14071 , n14074 );
xor ( n14076 , n14075 , n11959 );
buf ( n14077 , n6400 );
xor ( n14078 , n14076 , n14077 );
xor ( n14079 , n14078 , n12902 );
xor ( n14080 , n14079 , n13024 );
xor ( n14081 , n14068 , n14080 );
and ( n14082 , n14048 , n14081 );
xor ( n14083 , n11147 , n14082 );
xor ( n14084 , n14047 , n14083 );
xor ( n14085 , n13986 , n14084 );
xor ( n14086 , n6847 , n10488 );
xor ( n14087 , n14086 , n10504 );
not ( n14088 , n14087 );
xor ( n14089 , n7252 , n10864 );
xor ( n14090 , n14089 , n7159 );
and ( n14091 , n14088 , n14090 );
xor ( n14092 , n11440 , n14091 );
buf ( n14093 , n6401 );
xor ( n14094 , n14093 , n13774 );
xor ( n14095 , n14094 , n13018 );
not ( n14096 , n14095 );
xor ( n14097 , n8187 , n11132 );
xor ( n14098 , n14097 , n11146 );
and ( n14099 , n14096 , n14098 );
xor ( n14100 , n11483 , n14099 );
xor ( n14101 , n14092 , n14100 );
xor ( n14102 , n12563 , n9026 );
xor ( n14103 , n14102 , n9047 );
not ( n14104 , n14103 );
xor ( n14105 , n11762 , n13886 );
xor ( n14106 , n14105 , n12213 );
and ( n14107 , n14104 , n14106 );
xor ( n14108 , n11521 , n14107 );
xor ( n14109 , n14101 , n14108 );
xor ( n14110 , n12187 , n7274 );
xor ( n14111 , n14110 , n13798 );
not ( n14112 , n14111 );
xor ( n14113 , n10526 , n12302 );
xor ( n14114 , n14113 , n13273 );
and ( n14115 , n14112 , n14114 );
xor ( n14116 , n11559 , n14115 );
xor ( n14117 , n14109 , n14116 );
buf ( n14118 , n6402 );
xor ( n14119 , n7545 , n14118 );
buf ( n14120 , n6403 );
xor ( n14121 , n14119 , n14120 );
buf ( n14122 , n6404 );
xor ( n14123 , n14121 , n14122 );
buf ( n14124 , n6405 );
xor ( n14125 , n14123 , n14124 );
xor ( n14126 , n12696 , n14125 );
xor ( n14127 , n14126 , n14009 );
not ( n14128 , n14127 );
xor ( n14129 , n7770 , n12365 );
xor ( n14130 , n14129 , n12490 );
and ( n14131 , n14128 , n14130 );
xor ( n14132 , n11658 , n14131 );
xor ( n14133 , n14117 , n14132 );
xor ( n14134 , n14085 , n14133 );
and ( n14135 , n13979 , n14134 );
xor ( n14136 , n13808 , n14135 );
and ( n14137 , n14136 , n6475 );
or ( n14138 , n13621 , n14137 );
and ( n14139 , n13619 , n14138 );
buf ( n14140 , n14139 );
buf ( n14141 , n14140 );
not ( n14142 , n6469 );
not ( n14143 , n6475 );
and ( n14144 , n14143 , n7157 );
not ( n14145 , n6654 );
and ( n14146 , n14145 , n6517 );
xor ( n14147 , n13500 , n14146 );
not ( n14148 , n6696 );
and ( n14149 , n14148 , n6740 );
xor ( n14150 , n13528 , n14149 );
xor ( n14151 , n14147 , n14150 );
not ( n14152 , n6828 );
and ( n14153 , n14152 , n6873 );
xor ( n14154 , n13536 , n14153 );
xor ( n14155 , n14151 , n14154 );
not ( n14156 , n6962 );
and ( n14157 , n14156 , n7007 );
xor ( n14158 , n13565 , n14157 );
xor ( n14159 , n14155 , n14158 );
not ( n14160 , n7096 );
and ( n14161 , n14160 , n7135 );
xor ( n14162 , n13573 , n14161 );
xor ( n14163 , n14159 , n14162 );
xor ( n14164 , n6657 , n14163 );
xor ( n14165 , n9992 , n9464 );
xor ( n14166 , n14165 , n10929 );
not ( n14167 , n7231 );
and ( n14168 , n14167 , n7275 );
xor ( n14169 , n14166 , n14168 );
not ( n14170 , n6474 );
buf ( n14171 , n6406 );
and ( n14172 , n14170 , n14171 );
buf ( n14173 , n6407 );
xor ( n14174 , n14173 , n14171 );
and ( n14175 , n14174 , n6474 );
or ( n14176 , n14172 , n14175 );
not ( n14177 , n6474 );
buf ( n14178 , n6408 );
and ( n14179 , n14177 , n14178 );
buf ( n14180 , n6409 );
xor ( n14181 , n14180 , n14178 );
and ( n14182 , n14181 , n6474 );
or ( n14183 , n14179 , n14182 );
xor ( n14184 , n14176 , n14183 );
buf ( n14185 , n6410 );
xor ( n14186 , n14184 , n14185 );
buf ( n14187 , n6411 );
xor ( n14188 , n14186 , n14187 );
buf ( n14189 , n6412 );
xor ( n14190 , n14188 , n14189 );
xor ( n14191 , n9486 , n14190 );
xor ( n14192 , n14191 , n13591 );
not ( n14193 , n7332 );
and ( n14194 , n14193 , n7377 );
xor ( n14195 , n14192 , n14194 );
xor ( n14196 , n14169 , n14195 );
xor ( n14197 , n10501 , n10674 );
xor ( n14198 , n14197 , n6939 );
not ( n14199 , n7464 );
and ( n14200 , n14199 , n7466 );
xor ( n14201 , n14198 , n14200 );
xor ( n14202 , n14196 , n14201 );
xor ( n14203 , n12140 , n13842 );
xor ( n14204 , n14203 , n11949 );
not ( n14205 , n7538 );
and ( n14206 , n14205 , n7589 );
xor ( n14207 , n14204 , n14206 );
xor ( n14208 , n14202 , n14207 );
xor ( n14209 , n12278 , n11171 );
xor ( n14210 , n14209 , n6631 );
not ( n14211 , n7682 );
and ( n14212 , n14211 , n7733 );
xor ( n14213 , n14210 , n14212 );
xor ( n14214 , n14208 , n14213 );
xor ( n14215 , n14164 , n14214 );
not ( n14216 , n10841 );
and ( n14217 , n14216 , n8474 );
xor ( n14218 , n10837 , n14217 );
xor ( n14219 , n14218 , n10887 );
xor ( n14220 , n14219 , n11066 );
not ( n14221 , n14220 );
xor ( n14222 , n9849 , n12566 );
xor ( n14223 , n14222 , n11693 );
xor ( n14224 , n7120 , n12281 );
xor ( n14225 , n14224 , n12302 );
not ( n14226 , n14225 );
xor ( n14227 , n13586 , n11275 );
xor ( n14228 , n14227 , n9559 );
and ( n14229 , n14226 , n14228 );
xor ( n14230 , n14223 , n14229 );
xor ( n14231 , n6782 , n10309 );
xor ( n14232 , n14231 , n13367 );
xor ( n14233 , n12505 , n8388 );
xor ( n14234 , n14233 , n11998 );
not ( n14235 , n14234 );
xor ( n14236 , n9182 , n7112 );
xor ( n14237 , n14236 , n7134 );
and ( n14238 , n14235 , n14237 );
xor ( n14239 , n14232 , n14238 );
xor ( n14240 , n13687 , n7421 );
xor ( n14241 , n14240 , n12452 );
xor ( n14242 , n8055 , n7634 );
xor ( n14243 , n14242 , n7072 );
not ( n14244 , n14243 );
not ( n14245 , n6474 );
buf ( n14246 , n6413 );
and ( n14247 , n14245 , n14246 );
buf ( n14248 , n6414 );
xor ( n14249 , n14248 , n14246 );
and ( n14250 , n14249 , n6474 );
or ( n14251 , n14247 , n14250 );
xor ( n14252 , n14251 , n12727 );
xor ( n14253 , n14252 , n12742 );
and ( n14254 , n14244 , n14253 );
xor ( n14255 , n14241 , n14254 );
xor ( n14256 , n14239 , n14255 );
xor ( n14257 , n8201 , n11146 );
xor ( n14258 , n14257 , n9651 );
not ( n14259 , n14223 );
and ( n14260 , n14259 , n14225 );
xor ( n14261 , n14258 , n14260 );
xor ( n14262 , n14256 , n14261 );
xor ( n14263 , n7027 , n11031 );
xor ( n14264 , n14263 , n11052 );
xor ( n14265 , n13935 , n13018 );
xor ( n14266 , n14265 , n10394 );
not ( n14267 , n14266 );
xor ( n14268 , n8994 , n11741 );
xor ( n14269 , n14268 , n11763 );
and ( n14270 , n14267 , n14269 );
xor ( n14271 , n14264 , n14270 );
xor ( n14272 , n14262 , n14271 );
xor ( n14273 , n10572 , n6891 );
xor ( n14274 , n14273 , n6913 );
xor ( n14275 , n6630 , n12609 );
xor ( n14276 , n14275 , n10334 );
not ( n14277 , n14276 );
not ( n14278 , n6474 );
buf ( n14279 , n6415 );
and ( n14280 , n14278 , n14279 );
buf ( n14281 , n6416 );
xor ( n14282 , n14281 , n14279 );
and ( n14283 , n14282 , n6474 );
or ( n14284 , n14280 , n14283 );
not ( n14285 , n6474 );
buf ( n14286 , n6417 );
and ( n14287 , n14285 , n14286 );
buf ( n14288 , n6418 );
xor ( n14289 , n14288 , n14286 );
and ( n14290 , n14289 , n6474 );
or ( n14291 , n14287 , n14290 );
xor ( n14292 , n14284 , n14291 );
buf ( n14293 , n6419 );
xor ( n14294 , n14292 , n14293 );
buf ( n14295 , n6420 );
xor ( n14296 , n14294 , n14295 );
buf ( n14297 , n6421 );
xor ( n14298 , n14296 , n14297 );
xor ( n14299 , n10822 , n14298 );
not ( n14300 , n6474 );
buf ( n14301 , n6422 );
and ( n14302 , n14300 , n14301 );
buf ( n14303 , n6423 );
xor ( n14304 , n14303 , n14301 );
and ( n14305 , n14304 , n6474 );
or ( n14306 , n14302 , n14305 );
xor ( n14307 , n13815 , n14306 );
xor ( n14308 , n14307 , n9749 );
buf ( n14309 , n6424 );
xor ( n14310 , n14308 , n14309 );
buf ( n14311 , n6425 );
xor ( n14312 , n14310 , n14311 );
xor ( n14313 , n14299 , n14312 );
and ( n14314 , n14277 , n14313 );
xor ( n14315 , n14274 , n14314 );
xor ( n14316 , n14272 , n14315 );
xor ( n14317 , n14230 , n14316 );
xor ( n14318 , n12267 , n11171 );
xor ( n14319 , n14318 , n6631 );
xor ( n14320 , n13683 , n7421 );
xor ( n14321 , n14320 , n12452 );
not ( n14322 , n14321 );
xor ( n14323 , n6495 , n9973 );
xor ( n14324 , n14323 , n9995 );
and ( n14325 , n14322 , n14324 );
xor ( n14326 , n14319 , n14325 );
xor ( n14327 , n7934 , n10130 );
xor ( n14328 , n14327 , n10146 );
xor ( n14329 , n9347 , n6785 );
not ( n14330 , n6474 );
buf ( n14331 , n6426 );
and ( n14332 , n14330 , n14331 );
buf ( n14333 , n6427 );
xor ( n14334 , n14333 , n14331 );
and ( n14335 , n14334 , n6474 );
or ( n14336 , n14332 , n14335 );
not ( n14337 , n6474 );
buf ( n14338 , n6428 );
and ( n14339 , n14337 , n14338 );
buf ( n14340 , n6429 );
xor ( n14341 , n14340 , n14338 );
and ( n14342 , n14341 , n6474 );
or ( n14343 , n14339 , n14342 );
xor ( n14344 , n14336 , n14343 );
buf ( n14345 , n6430 );
xor ( n14346 , n14344 , n14345 );
xor ( n14347 , n14346 , n13354 );
buf ( n14348 , n6431 );
xor ( n14349 , n14347 , n14348 );
xor ( n14350 , n14329 , n14349 );
not ( n14351 , n14350 );
xor ( n14352 , n6712 , n10350 );
xor ( n14353 , n14352 , n9489 );
and ( n14354 , n14351 , n14353 );
xor ( n14355 , n14328 , n14354 );
xor ( n14356 , n14326 , n14355 );
xor ( n14357 , n6617 , n12609 );
xor ( n14358 , n14357 , n10334 );
xor ( n14359 , n8181 , n11132 );
xor ( n14360 , n14359 , n11146 );
not ( n14361 , n14360 );
xor ( n14362 , n13793 , n7181 );
xor ( n14363 , n14362 , n9002 );
and ( n14364 , n14361 , n14363 );
xor ( n14365 , n14358 , n14364 );
xor ( n14366 , n14356 , n14365 );
not ( n14367 , n6474 );
buf ( n14368 , n6432 );
and ( n14369 , n14367 , n14368 );
buf ( n14370 , n6433 );
xor ( n14371 , n14370 , n14368 );
and ( n14372 , n14371 , n6474 );
or ( n14373 , n14369 , n14372 );
xor ( n14374 , n14251 , n14373 );
buf ( n14375 , n6434 );
xor ( n14376 , n14374 , n14375 );
xor ( n14377 , n14376 , n12706 );
buf ( n14378 , n6435 );
xor ( n14379 , n14377 , n14378 );
xor ( n14380 , n13878 , n14379 );
not ( n14381 , n6474 );
buf ( n14382 , n6436 );
and ( n14383 , n14381 , n14382 );
buf ( n14384 , n6437 );
xor ( n14385 , n14384 , n14382 );
and ( n14386 , n14385 , n6474 );
or ( n14387 , n14383 , n14386 );
not ( n14388 , n6474 );
buf ( n14389 , n6438 );
and ( n14390 , n14388 , n14389 );
buf ( n14391 , n6439 );
xor ( n14392 , n14391 , n14389 );
and ( n14393 , n14392 , n6474 );
or ( n14394 , n14390 , n14393 );
xor ( n14395 , n14387 , n14394 );
buf ( n14396 , n6440 );
xor ( n14397 , n14395 , n14396 );
buf ( n14398 , n6441 );
xor ( n14399 , n14397 , n14398 );
buf ( n14400 , n6442 );
xor ( n14401 , n14399 , n14400 );
xor ( n14402 , n14380 , n14401 );
xor ( n14403 , n8510 , n7925 );
xor ( n14404 , n14403 , n6984 );
not ( n14405 , n14404 );
xor ( n14406 , n10039 , n11089 );
xor ( n14407 , n14406 , n11110 );
and ( n14408 , n14405 , n14407 );
xor ( n14409 , n14402 , n14408 );
xor ( n14410 , n14366 , n14409 );
xor ( n14411 , n9756 , n8950 );
xor ( n14412 , n14411 , n12581 );
xor ( n14413 , n13930 , n13018 );
xor ( n14414 , n14413 , n10394 );
not ( n14415 , n14414 );
xor ( n14416 , n9705 , n11949 );
xor ( n14417 , n14416 , n10574 );
and ( n14418 , n14415 , n14417 );
xor ( n14419 , n14412 , n14418 );
xor ( n14420 , n14410 , n14419 );
xor ( n14421 , n14317 , n14420 );
and ( n14422 , n14221 , n14421 );
xor ( n14423 , n14215 , n14422 );
and ( n14424 , n14423 , n6475 );
or ( n14425 , n14144 , n14424 );
and ( n14426 , n14142 , n14425 );
buf ( n14427 , n14426 );
buf ( n14428 , n14427 );
not ( n14429 , n6469 );
not ( n14430 , n6475 );
and ( n14431 , n14430 , n6887 );
xor ( n14432 , n11342 , n10022 );
xor ( n14433 , n14432 , n10044 );
xor ( n14434 , n9169 , n12111 );
xor ( n14435 , n14434 , n7910 );
not ( n14436 , n14435 );
xor ( n14437 , n10474 , n10652 );
xor ( n14438 , n14437 , n10674 );
and ( n14439 , n14436 , n14438 );
xor ( n14440 , n14433 , n14439 );
xor ( n14441 , n11106 , n7771 );
xor ( n14442 , n14441 , n7793 );
xor ( n14443 , n10103 , n9079 );
xor ( n14444 , n14443 , n9094 );
not ( n14445 , n14444 );
xor ( n14446 , n12466 , n10376 );
xor ( n14447 , n14446 , n10067 );
and ( n14448 , n14445 , n14447 );
xor ( n14449 , n14442 , n14448 );
xor ( n14450 , n7878 , n11520 );
xor ( n14451 , n14450 , n10625 );
xor ( n14452 , n8693 , n10170 );
xor ( n14453 , n14452 , n7030 );
not ( n14454 , n14453 );
xor ( n14455 , n11186 , n7494 );
xor ( n14456 , n14455 , n6850 );
and ( n14457 , n14454 , n14456 );
xor ( n14458 , n14451 , n14457 );
xor ( n14459 , n14449 , n14458 );
xor ( n14460 , n9916 , n11808 );
xor ( n14461 , n14460 , n12548 );
not ( n14462 , n6474 );
buf ( n14463 , n6443 );
and ( n14464 , n14462 , n14463 );
buf ( n14465 , n6444 );
xor ( n14466 , n14465 , n14463 );
and ( n14467 , n14466 , n6474 );
or ( n14468 , n14464 , n14467 );
xor ( n14469 , n11841 , n14468 );
xor ( n14470 , n14469 , n8553 );
buf ( n14471 , n6445 );
xor ( n14472 , n14470 , n14471 );
buf ( n14473 , n6446 );
xor ( n14474 , n14472 , n14473 );
xor ( n14475 , n6888 , n14474 );
xor ( n14476 , n14475 , n8972 );
not ( n14477 , n14476 );
xor ( n14478 , n12698 , n14125 );
xor ( n14479 , n14478 , n14009 );
and ( n14480 , n14477 , n14479 );
xor ( n14481 , n14461 , n14480 );
xor ( n14482 , n14459 , n14481 );
xor ( n14483 , n7458 , n8249 );
xor ( n14484 , n14483 , n6500 );
xor ( n14485 , n6808 , n13215 );
xor ( n14486 , n14485 , n11636 );
not ( n14487 , n14486 );
xor ( n14488 , n9122 , n12190 );
xor ( n14489 , n14488 , n6673 );
and ( n14490 , n14487 , n14489 );
xor ( n14491 , n14484 , n14490 );
xor ( n14492 , n14482 , n14491 );
xor ( n14493 , n8199 , n11146 );
xor ( n14494 , n14493 , n9651 );
not ( n14495 , n14433 );
and ( n14496 , n14495 , n14435 );
xor ( n14497 , n14494 , n14496 );
xor ( n14498 , n14492 , n14497 );
xor ( n14499 , n14440 , n14498 );
xor ( n14500 , n12648 , n14067 );
xor ( n14501 , n14500 , n14080 );
xor ( n14502 , n11873 , n9148 );
xor ( n14503 , n14502 , n9170 );
not ( n14504 , n14503 );
xor ( n14505 , n8689 , n10170 );
xor ( n14506 , n14505 , n7030 );
and ( n14507 , n14504 , n14506 );
xor ( n14508 , n14501 , n14507 );
xor ( n14509 , n10487 , n10652 );
xor ( n14510 , n14509 , n10674 );
xor ( n14511 , n7058 , n10836 );
xor ( n14512 , n14511 , n12822 );
not ( n14513 , n14512 );
xor ( n14514 , n9299 , n10105 );
xor ( n14515 , n14514 , n13774 );
and ( n14516 , n14513 , n14515 );
xor ( n14517 , n14510 , n14516 );
xor ( n14518 , n14508 , n14517 );
xor ( n14519 , n7587 , n8638 );
xor ( n14520 , n14519 , n8660 );
xor ( n14521 , n9156 , n12111 );
xor ( n14522 , n14521 , n7910 );
not ( n14523 , n14522 );
not ( n14524 , n6474 );
buf ( n14525 , n6447 );
and ( n14526 , n14524 , n14525 );
buf ( n14527 , n6448 );
xor ( n14528 , n14527 , n14525 );
and ( n14529 , n14528 , n6474 );
or ( n14530 , n14526 , n14529 );
xor ( n14531 , n14530 , n10285 );
xor ( n14532 , n14531 , n14474 );
and ( n14533 , n14523 , n14532 );
xor ( n14534 , n14520 , n14533 );
xor ( n14535 , n14518 , n14534 );
xor ( n14536 , n13797 , n7181 );
xor ( n14537 , n14536 , n9002 );
xor ( n14538 , n10201 , n9260 );
xor ( n14539 , n14538 , n13487 );
not ( n14540 , n14539 );
xor ( n14541 , n13640 , n11927 );
xor ( n14542 , n14541 , n11132 );
and ( n14543 , n14540 , n14542 );
xor ( n14544 , n14537 , n14543 );
xor ( n14545 , n14535 , n14544 );
xor ( n14546 , n9627 , n7883 );
xor ( n14547 , n14546 , n10731 );
xor ( n14548 , n12765 , n11905 );
xor ( n14549 , n14548 , n11865 );
not ( n14550 , n14549 );
xor ( n14551 , n9116 , n12190 );
xor ( n14552 , n14551 , n6673 );
and ( n14553 , n14550 , n14552 );
xor ( n14554 , n14547 , n14553 );
xor ( n14555 , n14545 , n14554 );
xor ( n14556 , n14499 , n14555 );
xor ( n14557 , n12565 , n9026 );
xor ( n14558 , n14557 , n9047 );
xor ( n14559 , n6703 , n10350 );
xor ( n14560 , n14559 , n9489 );
not ( n14561 , n14560 );
xor ( n14562 , n13209 , n10067 );
xor ( n14563 , n14562 , n10089 );
and ( n14564 , n14561 , n14563 );
xor ( n14565 , n14558 , n14564 );
xor ( n14566 , n9120 , n12190 );
xor ( n14567 , n14566 , n6673 );
not ( n14568 , n14558 );
and ( n14569 , n14568 , n14560 );
xor ( n14570 , n14567 , n14569 );
xor ( n14571 , n12668 , n14080 );
not ( n14572 , n6474 );
buf ( n14573 , n6449 );
and ( n14574 , n14572 , n14573 );
buf ( n14575 , n6450 );
xor ( n14576 , n14575 , n14573 );
and ( n14577 , n14576 , n6474 );
or ( n14578 , n14574 , n14577 );
xor ( n14579 , n14578 , n13229 );
xor ( n14580 , n14579 , n12702 );
buf ( n14581 , n6451 );
xor ( n14582 , n14580 , n14581 );
buf ( n14583 , n6452 );
xor ( n14584 , n14582 , n14583 );
xor ( n14585 , n14571 , n14584 );
xor ( n14586 , n9216 , n7134 );
xor ( n14587 , n14586 , n10527 );
not ( n14588 , n14587 );
xor ( n14589 , n10660 , n12779 );
xor ( n14590 , n14589 , n8092 );
and ( n14591 , n14588 , n14590 );
xor ( n14592 , n14585 , n14591 );
xor ( n14593 , n14570 , n14592 );
xor ( n14594 , n14028 , n8891 );
xor ( n14595 , n14594 , n8913 );
xor ( n14596 , n14348 , n13367 );
xor ( n14597 , n14596 , n10963 );
not ( n14598 , n14597 );
xor ( n14599 , n9475 , n14190 );
xor ( n14600 , n14599 , n13591 );
and ( n14601 , n14598 , n14600 );
xor ( n14602 , n14595 , n14601 );
xor ( n14603 , n14593 , n14602 );
xor ( n14604 , n9869 , n11693 );
xor ( n14605 , n14604 , n11714 );
xor ( n14606 , n8468 , n10193 );
xor ( n14607 , n14606 , n10209 );
not ( n14608 , n14607 );
xor ( n14609 , n11195 , n6850 );
xor ( n14610 , n14609 , n6872 );
and ( n14611 , n14608 , n14610 );
xor ( n14612 , n14605 , n14611 );
xor ( n14613 , n14603 , n14612 );
xor ( n14614 , n7418 , n6516 );
xor ( n14615 , n14614 , n13052 );
xor ( n14616 , n11274 , n13647 );
xor ( n14617 , n14616 , n8188 );
not ( n14618 , n14617 );
xor ( n14619 , n12289 , n6631 );
xor ( n14620 , n14619 , n6653 );
and ( n14621 , n14618 , n14620 );
xor ( n14622 , n14615 , n14621 );
xor ( n14623 , n14613 , n14622 );
xor ( n14624 , n14565 , n14623 );
xor ( n14625 , n14176 , n12040 );
xor ( n14626 , n14625 , n11275 );
xor ( n14627 , n12664 , n14080 );
xor ( n14628 , n14627 , n14584 );
not ( n14629 , n14628 );
xor ( n14630 , n6806 , n13215 );
xor ( n14631 , n14630 , n11636 );
and ( n14632 , n14629 , n14631 );
xor ( n14633 , n14626 , n14632 );
xor ( n14634 , n11851 , n13468 );
xor ( n14635 , n14634 , n9148 );
xor ( n14636 , n9536 , n9123 );
xor ( n14637 , n14636 , n7659 );
not ( n14638 , n14637 );
xor ( n14639 , n9576 , n8204 );
xor ( n14640 , n14639 , n12854 );
and ( n14641 , n14638 , n14640 );
xor ( n14642 , n14635 , n14641 );
xor ( n14643 , n14633 , n14642 );
xor ( n14644 , n11261 , n13647 );
xor ( n14645 , n14644 , n8188 );
xor ( n14646 , n11360 , n10044 );
xor ( n14647 , n14646 , n8891 );
not ( n14648 , n14647 );
xor ( n14649 , n10763 , n11187 );
xor ( n14650 , n14649 , n11201 );
and ( n14651 , n14648 , n14650 );
xor ( n14652 , n14645 , n14651 );
xor ( n14653 , n14643 , n14652 );
xor ( n14654 , n10496 , n10674 );
xor ( n14655 , n14654 , n6939 );
xor ( n14656 , n10569 , n6891 );
xor ( n14657 , n14656 , n6913 );
not ( n14658 , n14657 );
xor ( n14659 , n11026 , n11998 );
xor ( n14660 , n14659 , n7521 );
and ( n14661 , n14658 , n14660 );
xor ( n14662 , n14655 , n14661 );
xor ( n14663 , n14653 , n14662 );
xor ( n14664 , n10320 , n9439 );
not ( n14665 , n6474 );
buf ( n14666 , n6453 );
and ( n14667 , n14665 , n14666 );
buf ( n14668 , n6454 );
xor ( n14669 , n14668 , n14666 );
and ( n14670 , n14669 , n6474 );
or ( n14671 , n14667 , n14670 );
xor ( n14672 , n14671 , n12010 );
buf ( n14673 , n6455 );
xor ( n14674 , n14672 , n14673 );
buf ( n14675 , n6456 );
xor ( n14676 , n14674 , n14675 );
buf ( n14677 , n6457 );
xor ( n14678 , n14676 , n14677 );
xor ( n14679 , n14664 , n14678 );
xor ( n14680 , n8462 , n10193 );
xor ( n14681 , n14680 , n10209 );
not ( n14682 , n14681 );
xor ( n14683 , n7832 , n7399 );
xor ( n14684 , n14683 , n7421 );
and ( n14685 , n14682 , n14684 );
xor ( n14686 , n14679 , n14685 );
xor ( n14687 , n14663 , n14686 );
xor ( n14688 , n14624 , n14687 );
not ( n14689 , n14688 );
not ( n14690 , n11880 );
xor ( n14691 , n8132 , n7046 );
xor ( n14692 , n14691 , n8414 );
and ( n14693 , n14690 , n14692 );
xor ( n14694 , n11843 , n14693 );
xor ( n14695 , n14694 , n12044 );
xor ( n14696 , n14695 , n12250 );
and ( n14697 , n14689 , n14696 );
xor ( n14698 , n14556 , n14697 );
and ( n14699 , n14698 , n6475 );
or ( n14700 , n14431 , n14699 );
and ( n14701 , n14429 , n14700 );
buf ( n14702 , n14701 );
buf ( n14703 , n14702 );
not ( n14704 , n6469 );
not ( n14705 , n6475 );
and ( n14706 , n14705 , n11919 );
xor ( n14707 , n7436 , n8227 );
xor ( n14708 , n14707 , n8249 );
xor ( n14709 , n8619 , n7837 );
xor ( n14710 , n14709 , n13690 );
not ( n14711 , n14710 );
xor ( n14712 , n9488 , n14190 );
xor ( n14713 , n14712 , n13591 );
and ( n14714 , n14711 , n14713 );
xor ( n14715 , n14708 , n14714 );
xor ( n14716 , n11548 , n9816 );
xor ( n14717 , n14716 , n6811 );
xor ( n14718 , n12447 , n13052 );
xor ( n14719 , n14718 , n10376 );
not ( n14720 , n14719 );
xor ( n14721 , n10861 , n9534 );
xor ( n14722 , n14721 , n9543 );
and ( n14723 , n14720 , n14722 );
xor ( n14724 , n14717 , n14723 );
xor ( n14725 , n6577 , n7732 );
xor ( n14726 , n14725 , n8076 );
xor ( n14727 , n13642 , n11927 );
xor ( n14728 , n14727 , n11132 );
not ( n14729 , n14728 );
xor ( n14730 , n13212 , n10067 );
xor ( n14731 , n14730 , n10089 );
and ( n14732 , n14729 , n14731 );
xor ( n14733 , n14726 , n14732 );
xor ( n14734 , n14724 , n14733 );
xor ( n14735 , n10983 , n12854 );
not ( n14736 , n6474 );
buf ( n14737 , n6458 );
and ( n14738 , n14736 , n14737 );
buf ( n14739 , n6459 );
xor ( n14740 , n14739 , n14737 );
and ( n14741 , n14740 , n6474 );
or ( n14742 , n14738 , n14741 );
not ( n14743 , n6474 );
buf ( n14744 , n6460 );
and ( n14745 , n14743 , n14744 );
buf ( n14746 , n6461 );
xor ( n14747 , n14746 , n14744 );
and ( n14748 , n14747 , n6474 );
or ( n14749 , n14745 , n14748 );
xor ( n14750 , n14742 , n14749 );
buf ( n14751 , n6462 );
xor ( n14752 , n14750 , n14751 );
buf ( n14753 , n6463 );
xor ( n14754 , n14752 , n14753 );
buf ( n14755 , n6464 );
xor ( n14756 , n14754 , n14755 );
xor ( n14757 , n14735 , n14756 );
xor ( n14758 , n14375 , n12727 );
xor ( n14759 , n14758 , n12742 );
not ( n14760 , n14759 );
buf ( n14761 , n6465 );
xor ( n14762 , n14761 , n11833 );
xor ( n14763 , n14762 , n12365 );
and ( n14764 , n14760 , n14763 );
xor ( n14765 , n14757 , n14764 );
xor ( n14766 , n14734 , n14765 );
xor ( n14767 , n7223 , n10263 );
xor ( n14768 , n14767 , n10285 );
xor ( n14769 , n8361 , n8913 );
xor ( n14770 , n14769 , n13392 );
not ( n14771 , n14770 );
xor ( n14772 , n8333 , n10905 );
xor ( n14773 , n14772 , n9378 );
and ( n14774 , n14771 , n14773 );
xor ( n14775 , n14768 , n14774 );
xor ( n14776 , n14766 , n14775 );
xor ( n14777 , n9914 , n11808 );
xor ( n14778 , n14777 , n12548 );
not ( n14779 , n14708 );
and ( n14780 , n14779 , n14710 );
xor ( n14781 , n14778 , n14780 );
xor ( n14782 , n14776 , n14781 );
xor ( n14783 , n14715 , n14782 );
xor ( n14784 , n14783 , n14623 );
xor ( n14785 , n8740 , n11252 );
xor ( n14786 , n14785 , n8269 );
not ( n14787 , n14501 );
and ( n14788 , n14787 , n14503 );
xor ( n14789 , n14786 , n14788 );
xor ( n14790 , n12486 , n8366 );
xor ( n14791 , n14790 , n8388 );
not ( n14792 , n14786 );
and ( n14793 , n14792 , n14501 );
xor ( n14794 , n14791 , n14793 );
xor ( n14795 , n8512 , n7925 );
xor ( n14796 , n14795 , n6984 );
xor ( n14797 , n11028 , n11998 );
xor ( n14798 , n14797 , n7521 );
not ( n14799 , n14798 );
and ( n14800 , n14799 , n14510 );
xor ( n14801 , n14796 , n14800 );
xor ( n14802 , n14794 , n14801 );
xor ( n14803 , n13131 , n9895 );
xor ( n14804 , n14803 , n7612 );
xor ( n14805 , n7438 , n8227 );
xor ( n14806 , n14805 , n8249 );
not ( n14807 , n14806 );
and ( n14808 , n14807 , n14520 );
xor ( n14809 , n14804 , n14808 );
xor ( n14810 , n14802 , n14809 );
xor ( n14811 , n9969 , n8622 );
xor ( n14812 , n14811 , n9464 );
xor ( n14813 , n10086 , n12671 );
xor ( n14814 , n14813 , n13560 );
not ( n14815 , n14814 );
and ( n14816 , n14815 , n14537 );
xor ( n14817 , n14812 , n14816 );
xor ( n14818 , n14810 , n14817 );
xor ( n14819 , n10708 , n11604 );
xor ( n14820 , n14819 , n11345 );
not ( n14821 , n6474 );
buf ( n14822 , n6466 );
and ( n14823 , n14821 , n14822 );
buf ( n14824 , n6467 );
xor ( n14825 , n14824 , n14822 );
and ( n14826 , n14825 , n6474 );
or ( n14827 , n14823 , n14826 );
xor ( n14828 , n14827 , n12343 );
xor ( n14829 , n14828 , n13969 );
xor ( n14830 , n14829 , n14761 );
buf ( n14831 , n6468 );
xor ( n14832 , n14830 , n14831 );
xor ( n14833 , n11086 , n14832 );
xor ( n14834 , n14833 , n7771 );
not ( n14835 , n14834 );
and ( n14836 , n14835 , n14547 );
xor ( n14837 , n14820 , n14836 );
xor ( n14838 , n14818 , n14837 );
xor ( n14839 , n14789 , n14838 );
xor ( n14840 , n14839 , n13905 );
not ( n14841 , n14840 );
not ( n14842 , n13663 );
xor ( n14843 , n10923 , n9794 );
xor ( n14844 , n14843 , n9816 );
and ( n14845 , n14842 , n14844 );
xor ( n14846 , n13660 , n14845 );
xor ( n14847 , n14846 , n13730 );
xor ( n14848 , n14847 , n13807 );
and ( n14849 , n14841 , n14848 );
xor ( n14850 , n14784 , n14849 );
and ( n14851 , n14850 , n6475 );
or ( n14852 , n14706 , n14851 );
and ( n14853 , n14704 , n14852 );
buf ( n14854 , n14853 );
buf ( n14855 , n14854 );
not ( n14856 , n6469 );
not ( n14857 , n6475 );
and ( n14858 , n14857 , n6860 );
xor ( n14859 , n11301 , n8159 );
xor ( n14860 , n14859 , n12566 );
xor ( n14861 , n10021 , n14756 );
xor ( n14862 , n14861 , n11089 );
not ( n14863 , n14862 );
xor ( n14864 , n8027 , n7612 );
xor ( n14865 , n14864 , n7634 );
and ( n14866 , n14863 , n14865 );
xor ( n14867 , n14860 , n14866 );
xor ( n14868 , n12138 , n13842 );
xor ( n14869 , n14868 , n11949 );
not ( n14870 , n14860 );
and ( n14871 , n14870 , n14862 );
xor ( n14872 , n14869 , n14871 );
xor ( n14873 , n7089 , n12822 );
xor ( n14874 , n14873 , n13315 );
xor ( n14875 , n9729 , n10574 );
xor ( n14876 , n14875 , n10595 );
not ( n14877 , n14876 );
xor ( n14878 , n12406 , n8291 );
xor ( n14879 , n14878 , n9921 );
and ( n14880 , n14877 , n14879 );
xor ( n14881 , n14874 , n14880 );
xor ( n14882 , n14872 , n14881 );
xor ( n14883 , n6780 , n10309 );
xor ( n14884 , n14883 , n13367 );
xor ( n14885 , n10347 , n14678 );
xor ( n14886 , n14885 , n14190 );
not ( n14887 , n14886 );
xor ( n14888 , n10169 , n12506 );
xor ( n14889 , n14888 , n11031 );
and ( n14890 , n14887 , n14889 );
xor ( n14891 , n14884 , n14890 );
xor ( n14892 , n14882 , n14891 );
xor ( n14893 , n11270 , n13647 );
xor ( n14894 , n14893 , n8188 );
xor ( n14895 , n11364 , n10044 );
xor ( n14896 , n14895 , n8891 );
not ( n14897 , n14896 );
xor ( n14898 , n12944 , n7360 );
xor ( n14899 , n14898 , n7376 );
and ( n14900 , n14897 , n14899 );
xor ( n14901 , n14894 , n14900 );
xor ( n14902 , n14892 , n14901 );
xor ( n14903 , n9601 , n7861 );
xor ( n14904 , n14903 , n7883 );
xor ( n14905 , n8514 , n7925 );
xor ( n14906 , n14905 , n6984 );
not ( n14907 , n14906 );
xor ( n14908 , n14297 , n13487 );
xor ( n14909 , n14908 , n9770 );
and ( n14910 , n14907 , n14909 );
xor ( n14911 , n14904 , n14910 );
xor ( n14912 , n14902 , n14911 );
xor ( n14913 , n14867 , n14912 );
xor ( n14914 , n14831 , n11833 );
xor ( n14915 , n14914 , n12365 );
xor ( n14916 , n10800 , n10209 );
xor ( n14917 , n14916 , n14298 );
not ( n14918 , n14917 );
xor ( n14919 , n9725 , n10574 );
xor ( n14920 , n14919 , n10595 );
and ( n14921 , n14918 , n14920 );
xor ( n14922 , n14915 , n14921 );
xor ( n14923 , n11807 , n10416 );
xor ( n14924 , n14923 , n13135 );
xor ( n14925 , n9109 , n12190 );
xor ( n14926 , n14925 , n6673 );
not ( n14927 , n14926 );
xor ( n14928 , n7530 , n11304 );
xor ( n14929 , n14928 , n9850 );
and ( n14930 , n14927 , n14929 );
xor ( n14931 , n14924 , n14930 );
xor ( n14932 , n14922 , n14931 );
xor ( n14933 , n11997 , n7994 );
xor ( n14934 , n14933 , n8016 );
xor ( n14935 , n14284 , n13487 );
xor ( n14936 , n14935 , n9770 );
not ( n14937 , n14936 );
xor ( n14938 , n10327 , n9439 );
xor ( n14939 , n14938 , n14678 );
and ( n14940 , n14937 , n14939 );
xor ( n14941 , n14934 , n14940 );
xor ( n14942 , n14932 , n14941 );
xor ( n14943 , n10223 , n9290 );
xor ( n14944 , n14943 , n9306 );
xor ( n14945 , n7245 , n10864 );
xor ( n14946 , n14945 , n7159 );
not ( n14947 , n14946 );
xor ( n14948 , n6932 , n8092 );
xor ( n14949 , n14948 , n8114 );
and ( n14950 , n14947 , n14949 );
xor ( n14951 , n14944 , n14950 );
xor ( n14952 , n14942 , n14951 );
xor ( n14953 , n8949 , n7095 );
xor ( n14954 , n14953 , n8799 );
xor ( n14955 , n9883 , n8447 );
xor ( n14956 , n14955 , n8469 );
not ( n14957 , n14956 );
xor ( n14958 , n12938 , n7360 );
xor ( n14959 , n14958 , n7376 );
and ( n14960 , n14957 , n14959 );
xor ( n14961 , n14954 , n14960 );
xor ( n14962 , n14952 , n14961 );
xor ( n14963 , n14913 , n14962 );
xor ( n14964 , n10088 , n12671 );
xor ( n14965 , n14964 , n13560 );
xor ( n14966 , n11039 , n7521 );
xor ( n14967 , n14966 , n7537 );
not ( n14968 , n14967 );
xor ( n14969 , n8197 , n11146 );
xor ( n14970 , n14969 , n9651 );
and ( n14971 , n14968 , n14970 );
xor ( n14972 , n14965 , n14971 );
xor ( n14973 , n11602 , n10990 );
xor ( n14974 , n14973 , n10022 );
xor ( n14975 , n9416 , n10527 );
xor ( n14976 , n14975 , n10549 );
not ( n14977 , n14976 );
xor ( n14978 , n7574 , n8638 );
xor ( n14979 , n14978 , n8660 );
and ( n14980 , n14977 , n14979 );
xor ( n14981 , n14974 , n14980 );
xor ( n14982 , n13092 , n6939 );
xor ( n14983 , n14982 , n6961 );
not ( n14984 , n14965 );
and ( n14985 , n14984 , n14967 );
xor ( n14986 , n14983 , n14985 );
xor ( n14987 , n14981 , n14986 );
xor ( n14988 , n7609 , n8469 );
xor ( n14989 , n14988 , n10814 );
xor ( n14990 , n13646 , n11927 );
xor ( n14991 , n14990 , n11132 );
not ( n14992 , n14991 );
xor ( n14993 , n8646 , n12871 );
xor ( n14994 , n14993 , n9079 );
and ( n14995 , n14992 , n14994 );
xor ( n14996 , n14989 , n14995 );
xor ( n14997 , n14987 , n14996 );
xor ( n14998 , n10331 , n9439 );
xor ( n14999 , n14998 , n14678 );
xor ( n15000 , n7398 , n6500 );
xor ( n15001 , n15000 , n6516 );
not ( n15002 , n15001 );
xor ( n15003 , n7986 , n8710 );
xor ( n15004 , n15003 , n8137 );
and ( n15005 , n15002 , n15004 );
xor ( n15006 , n14999 , n15005 );
xor ( n15007 , n14997 , n15006 );
xor ( n15008 , n14398 , n12742 );
xor ( n15009 , n15008 , n7494 );
xor ( n15010 , n10464 , n10246 );
xor ( n15011 , n15010 , n11252 );
not ( n15012 , n15011 );
xor ( n15013 , n14578 , n11981 );
xor ( n15014 , n15013 , n7566 );
and ( n15015 , n15012 , n15014 );
xor ( n15016 , n15009 , n15015 );
xor ( n15017 , n15007 , n15016 );
xor ( n15018 , n14972 , n15017 );
xor ( n15019 , n12864 , n7376 );
xor ( n15020 , n15019 , n10465 );
xor ( n15021 , n13089 , n6939 );
xor ( n15022 , n15021 , n6961 );
not ( n15023 , n15022 );
xor ( n15024 , n12774 , n11905 );
xor ( n15025 , n15024 , n11865 );
and ( n15026 , n15023 , n15025 );
xor ( n15027 , n15020 , n15026 );
xor ( n15028 , n11290 , n8159 );
xor ( n15029 , n15028 , n12566 );
xor ( n15030 , n10706 , n11604 );
xor ( n15031 , n15030 , n11345 );
not ( n15032 , n15031 );
xor ( n15033 , n8760 , n8269 );
xor ( n15034 , n15033 , n8291 );
and ( n15035 , n15032 , n15034 );
xor ( n15036 , n15029 , n15035 );
xor ( n15037 , n15027 , n15036 );
xor ( n15038 , n10451 , n10246 );
xor ( n15039 , n15038 , n11252 );
xor ( n15040 , n9890 , n8447 );
xor ( n15041 , n15040 , n8469 );
not ( n15042 , n15041 );
xor ( n15043 , n8383 , n13392 );
xor ( n15044 , n15043 , n7994 );
and ( n15045 , n15042 , n15044 );
xor ( n15046 , n15039 , n15045 );
xor ( n15047 , n15037 , n15046 );
xor ( n15048 , n7038 , n11052 );
xor ( n15049 , n15048 , n8314 );
xor ( n15050 , n7151 , n9543 );
xor ( n15051 , n15050 , n13427 );
not ( n15052 , n15051 );
xor ( n15053 , n8945 , n7095 );
xor ( n15054 , n15053 , n8799 );
and ( n15055 , n15052 , n15054 );
xor ( n15056 , n15049 , n15055 );
xor ( n15057 , n15047 , n15056 );
xor ( n15058 , n13509 , n11427 );
xor ( n15059 , n15058 , n12945 );
xor ( n15060 , n7393 , n6500 );
xor ( n15061 , n15060 , n6516 );
not ( n15062 , n15061 );
xor ( n15063 , n13881 , n14379 );
xor ( n15064 , n15063 , n14401 );
and ( n15065 , n15062 , n15064 );
xor ( n15066 , n15059 , n15065 );
xor ( n15067 , n15057 , n15066 );
xor ( n15068 , n15018 , n15067 );
not ( n15069 , n15068 );
not ( n15070 , n13867 );
xor ( n15071 , n8464 , n10193 );
xor ( n15072 , n15071 , n10209 );
and ( n15073 , n15070 , n15072 );
xor ( n15074 , n13864 , n15073 );
xor ( n15075 , n15074 , n13905 );
xor ( n15076 , n15075 , n13977 );
and ( n15077 , n15069 , n15076 );
xor ( n15078 , n14963 , n15077 );
and ( n15079 , n15078 , n6475 );
or ( n15080 , n14858 , n15079 );
and ( n15081 , n14856 , n15080 );
buf ( n15082 , n15081 );
buf ( n15083 , n15082 );
endmodule

